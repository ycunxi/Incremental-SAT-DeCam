module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1191(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1192(.a(gate16inter0), .b(s_92), .O(gate16inter1));
  and2  gate1193(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1194(.a(s_92), .O(gate16inter3));
  inv1  gate1195(.a(s_93), .O(gate16inter4));
  nand2 gate1196(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1197(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1198(.a(G15), .O(gate16inter7));
  inv1  gate1199(.a(G16), .O(gate16inter8));
  nand2 gate1200(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1201(.a(s_93), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1202(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1203(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1204(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate757(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate758(.a(gate21inter0), .b(s_30), .O(gate21inter1));
  and2  gate759(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate760(.a(s_30), .O(gate21inter3));
  inv1  gate761(.a(s_31), .O(gate21inter4));
  nand2 gate762(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate763(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate764(.a(G25), .O(gate21inter7));
  inv1  gate765(.a(G26), .O(gate21inter8));
  nand2 gate766(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate767(.a(s_31), .b(gate21inter3), .O(gate21inter10));
  nor2  gate768(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate769(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate770(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1681(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1682(.a(gate27inter0), .b(s_162), .O(gate27inter1));
  and2  gate1683(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1684(.a(s_162), .O(gate27inter3));
  inv1  gate1685(.a(s_163), .O(gate27inter4));
  nand2 gate1686(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1687(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1688(.a(G2), .O(gate27inter7));
  inv1  gate1689(.a(G6), .O(gate27inter8));
  nand2 gate1690(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1691(.a(s_163), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1692(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1693(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1694(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1849(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1850(.a(gate34inter0), .b(s_186), .O(gate34inter1));
  and2  gate1851(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1852(.a(s_186), .O(gate34inter3));
  inv1  gate1853(.a(s_187), .O(gate34inter4));
  nand2 gate1854(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1855(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1856(.a(G25), .O(gate34inter7));
  inv1  gate1857(.a(G29), .O(gate34inter8));
  nand2 gate1858(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1859(.a(s_187), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1860(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1861(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1862(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1121(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1122(.a(gate38inter0), .b(s_82), .O(gate38inter1));
  and2  gate1123(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1124(.a(s_82), .O(gate38inter3));
  inv1  gate1125(.a(s_83), .O(gate38inter4));
  nand2 gate1126(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1127(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1128(.a(G27), .O(gate38inter7));
  inv1  gate1129(.a(G31), .O(gate38inter8));
  nand2 gate1130(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1131(.a(s_83), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1132(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1133(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1134(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1037(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1038(.a(gate39inter0), .b(s_70), .O(gate39inter1));
  and2  gate1039(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1040(.a(s_70), .O(gate39inter3));
  inv1  gate1041(.a(s_71), .O(gate39inter4));
  nand2 gate1042(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1043(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1044(.a(G20), .O(gate39inter7));
  inv1  gate1045(.a(G24), .O(gate39inter8));
  nand2 gate1046(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1047(.a(s_71), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1048(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1049(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1050(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1093(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1094(.a(gate44inter0), .b(s_78), .O(gate44inter1));
  and2  gate1095(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1096(.a(s_78), .O(gate44inter3));
  inv1  gate1097(.a(s_79), .O(gate44inter4));
  nand2 gate1098(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1099(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1100(.a(G4), .O(gate44inter7));
  inv1  gate1101(.a(G269), .O(gate44inter8));
  nand2 gate1102(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1103(.a(s_79), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1104(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1105(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1106(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1247(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1248(.a(gate46inter0), .b(s_100), .O(gate46inter1));
  and2  gate1249(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1250(.a(s_100), .O(gate46inter3));
  inv1  gate1251(.a(s_101), .O(gate46inter4));
  nand2 gate1252(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1253(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1254(.a(G6), .O(gate46inter7));
  inv1  gate1255(.a(G272), .O(gate46inter8));
  nand2 gate1256(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1257(.a(s_101), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1258(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1259(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1260(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate701(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate702(.a(gate50inter0), .b(s_22), .O(gate50inter1));
  and2  gate703(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate704(.a(s_22), .O(gate50inter3));
  inv1  gate705(.a(s_23), .O(gate50inter4));
  nand2 gate706(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate707(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate708(.a(G10), .O(gate50inter7));
  inv1  gate709(.a(G278), .O(gate50inter8));
  nand2 gate710(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate711(.a(s_23), .b(gate50inter3), .O(gate50inter10));
  nor2  gate712(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate713(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate714(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate645(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate646(.a(gate52inter0), .b(s_14), .O(gate52inter1));
  and2  gate647(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate648(.a(s_14), .O(gate52inter3));
  inv1  gate649(.a(s_15), .O(gate52inter4));
  nand2 gate650(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate651(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate652(.a(G12), .O(gate52inter7));
  inv1  gate653(.a(G281), .O(gate52inter8));
  nand2 gate654(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate655(.a(s_15), .b(gate52inter3), .O(gate52inter10));
  nor2  gate656(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate657(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate658(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate715(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate716(.a(gate54inter0), .b(s_24), .O(gate54inter1));
  and2  gate717(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate718(.a(s_24), .O(gate54inter3));
  inv1  gate719(.a(s_25), .O(gate54inter4));
  nand2 gate720(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate721(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate722(.a(G14), .O(gate54inter7));
  inv1  gate723(.a(G284), .O(gate54inter8));
  nand2 gate724(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate725(.a(s_25), .b(gate54inter3), .O(gate54inter10));
  nor2  gate726(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate727(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate728(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1527(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1528(.a(gate55inter0), .b(s_140), .O(gate55inter1));
  and2  gate1529(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1530(.a(s_140), .O(gate55inter3));
  inv1  gate1531(.a(s_141), .O(gate55inter4));
  nand2 gate1532(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1533(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1534(.a(G15), .O(gate55inter7));
  inv1  gate1535(.a(G287), .O(gate55inter8));
  nand2 gate1536(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1537(.a(s_141), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1538(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1539(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1540(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1723(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1724(.a(gate56inter0), .b(s_168), .O(gate56inter1));
  and2  gate1725(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1726(.a(s_168), .O(gate56inter3));
  inv1  gate1727(.a(s_169), .O(gate56inter4));
  nand2 gate1728(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1729(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1730(.a(G16), .O(gate56inter7));
  inv1  gate1731(.a(G287), .O(gate56inter8));
  nand2 gate1732(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1733(.a(s_169), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1734(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1735(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1736(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1779(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1780(.a(gate60inter0), .b(s_176), .O(gate60inter1));
  and2  gate1781(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1782(.a(s_176), .O(gate60inter3));
  inv1  gate1783(.a(s_177), .O(gate60inter4));
  nand2 gate1784(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1785(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1786(.a(G20), .O(gate60inter7));
  inv1  gate1787(.a(G293), .O(gate60inter8));
  nand2 gate1788(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1789(.a(s_177), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1790(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1791(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1792(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1107(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1108(.a(gate72inter0), .b(s_80), .O(gate72inter1));
  and2  gate1109(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1110(.a(s_80), .O(gate72inter3));
  inv1  gate1111(.a(s_81), .O(gate72inter4));
  nand2 gate1112(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1113(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1114(.a(G32), .O(gate72inter7));
  inv1  gate1115(.a(G311), .O(gate72inter8));
  nand2 gate1116(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1117(.a(s_81), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1118(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1119(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1120(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1653(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1654(.a(gate81inter0), .b(s_158), .O(gate81inter1));
  and2  gate1655(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1656(.a(s_158), .O(gate81inter3));
  inv1  gate1657(.a(s_159), .O(gate81inter4));
  nand2 gate1658(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1659(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1660(.a(G3), .O(gate81inter7));
  inv1  gate1661(.a(G326), .O(gate81inter8));
  nand2 gate1662(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1663(.a(s_159), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1664(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1665(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1666(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate869(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate870(.a(gate86inter0), .b(s_46), .O(gate86inter1));
  and2  gate871(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate872(.a(s_46), .O(gate86inter3));
  inv1  gate873(.a(s_47), .O(gate86inter4));
  nand2 gate874(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate875(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate876(.a(G8), .O(gate86inter7));
  inv1  gate877(.a(G332), .O(gate86inter8));
  nand2 gate878(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate879(.a(s_47), .b(gate86inter3), .O(gate86inter10));
  nor2  gate880(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate881(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate882(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1499(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1500(.a(gate93inter0), .b(s_136), .O(gate93inter1));
  and2  gate1501(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1502(.a(s_136), .O(gate93inter3));
  inv1  gate1503(.a(s_137), .O(gate93inter4));
  nand2 gate1504(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1505(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1506(.a(G18), .O(gate93inter7));
  inv1  gate1507(.a(G344), .O(gate93inter8));
  nand2 gate1508(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1509(.a(s_137), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1510(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1511(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1512(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1709(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1710(.a(gate96inter0), .b(s_166), .O(gate96inter1));
  and2  gate1711(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1712(.a(s_166), .O(gate96inter3));
  inv1  gate1713(.a(s_167), .O(gate96inter4));
  nand2 gate1714(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1715(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1716(.a(G30), .O(gate96inter7));
  inv1  gate1717(.a(G347), .O(gate96inter8));
  nand2 gate1718(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1719(.a(s_167), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1720(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1721(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1722(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1177(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1178(.a(gate105inter0), .b(s_90), .O(gate105inter1));
  and2  gate1179(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1180(.a(s_90), .O(gate105inter3));
  inv1  gate1181(.a(s_91), .O(gate105inter4));
  nand2 gate1182(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1183(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1184(.a(G362), .O(gate105inter7));
  inv1  gate1185(.a(G363), .O(gate105inter8));
  nand2 gate1186(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1187(.a(s_91), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1188(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1189(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1190(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate953(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate954(.a(gate108inter0), .b(s_58), .O(gate108inter1));
  and2  gate955(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate956(.a(s_58), .O(gate108inter3));
  inv1  gate957(.a(s_59), .O(gate108inter4));
  nand2 gate958(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate959(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate960(.a(G368), .O(gate108inter7));
  inv1  gate961(.a(G369), .O(gate108inter8));
  nand2 gate962(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate963(.a(s_59), .b(gate108inter3), .O(gate108inter10));
  nor2  gate964(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate965(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate966(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1135(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1136(.a(gate115inter0), .b(s_84), .O(gate115inter1));
  and2  gate1137(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1138(.a(s_84), .O(gate115inter3));
  inv1  gate1139(.a(s_85), .O(gate115inter4));
  nand2 gate1140(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1141(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1142(.a(G382), .O(gate115inter7));
  inv1  gate1143(.a(G383), .O(gate115inter8));
  nand2 gate1144(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1145(.a(s_85), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1146(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1147(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1148(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1373(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1374(.a(gate124inter0), .b(s_118), .O(gate124inter1));
  and2  gate1375(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1376(.a(s_118), .O(gate124inter3));
  inv1  gate1377(.a(s_119), .O(gate124inter4));
  nand2 gate1378(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1379(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1380(.a(G400), .O(gate124inter7));
  inv1  gate1381(.a(G401), .O(gate124inter8));
  nand2 gate1382(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1383(.a(s_119), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1384(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1385(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1386(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1051(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1052(.a(gate127inter0), .b(s_72), .O(gate127inter1));
  and2  gate1053(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1054(.a(s_72), .O(gate127inter3));
  inv1  gate1055(.a(s_73), .O(gate127inter4));
  nand2 gate1056(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1057(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1058(.a(G406), .O(gate127inter7));
  inv1  gate1059(.a(G407), .O(gate127inter8));
  nand2 gate1060(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1061(.a(s_73), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1062(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1063(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1064(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate813(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate814(.a(gate132inter0), .b(s_38), .O(gate132inter1));
  and2  gate815(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate816(.a(s_38), .O(gate132inter3));
  inv1  gate817(.a(s_39), .O(gate132inter4));
  nand2 gate818(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate819(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate820(.a(G416), .O(gate132inter7));
  inv1  gate821(.a(G417), .O(gate132inter8));
  nand2 gate822(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate823(.a(s_39), .b(gate132inter3), .O(gate132inter10));
  nor2  gate824(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate825(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate826(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1541(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1542(.a(gate134inter0), .b(s_142), .O(gate134inter1));
  and2  gate1543(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1544(.a(s_142), .O(gate134inter3));
  inv1  gate1545(.a(s_143), .O(gate134inter4));
  nand2 gate1546(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1547(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1548(.a(G420), .O(gate134inter7));
  inv1  gate1549(.a(G421), .O(gate134inter8));
  nand2 gate1550(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1551(.a(s_143), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1552(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1553(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1554(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate771(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate772(.a(gate136inter0), .b(s_32), .O(gate136inter1));
  and2  gate773(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate774(.a(s_32), .O(gate136inter3));
  inv1  gate775(.a(s_33), .O(gate136inter4));
  nand2 gate776(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate777(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate778(.a(G424), .O(gate136inter7));
  inv1  gate779(.a(G425), .O(gate136inter8));
  nand2 gate780(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate781(.a(s_33), .b(gate136inter3), .O(gate136inter10));
  nor2  gate782(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate783(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate784(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate981(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate982(.a(gate140inter0), .b(s_62), .O(gate140inter1));
  and2  gate983(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate984(.a(s_62), .O(gate140inter3));
  inv1  gate985(.a(s_63), .O(gate140inter4));
  nand2 gate986(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate987(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate988(.a(G444), .O(gate140inter7));
  inv1  gate989(.a(G447), .O(gate140inter8));
  nand2 gate990(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate991(.a(s_63), .b(gate140inter3), .O(gate140inter10));
  nor2  gate992(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate993(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate994(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1457(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1458(.a(gate145inter0), .b(s_130), .O(gate145inter1));
  and2  gate1459(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1460(.a(s_130), .O(gate145inter3));
  inv1  gate1461(.a(s_131), .O(gate145inter4));
  nand2 gate1462(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1463(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1464(.a(G474), .O(gate145inter7));
  inv1  gate1465(.a(G477), .O(gate145inter8));
  nand2 gate1466(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1467(.a(s_131), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1468(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1469(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1470(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1835(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1836(.a(gate148inter0), .b(s_184), .O(gate148inter1));
  and2  gate1837(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1838(.a(s_184), .O(gate148inter3));
  inv1  gate1839(.a(s_185), .O(gate148inter4));
  nand2 gate1840(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1841(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1842(.a(G492), .O(gate148inter7));
  inv1  gate1843(.a(G495), .O(gate148inter8));
  nand2 gate1844(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1845(.a(s_185), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1846(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1847(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1848(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate1583(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1584(.a(gate149inter0), .b(s_148), .O(gate149inter1));
  and2  gate1585(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1586(.a(s_148), .O(gate149inter3));
  inv1  gate1587(.a(s_149), .O(gate149inter4));
  nand2 gate1588(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1589(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1590(.a(G498), .O(gate149inter7));
  inv1  gate1591(.a(G501), .O(gate149inter8));
  nand2 gate1592(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1593(.a(s_149), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1594(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1595(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1596(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1471(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1472(.a(gate151inter0), .b(s_132), .O(gate151inter1));
  and2  gate1473(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1474(.a(s_132), .O(gate151inter3));
  inv1  gate1475(.a(s_133), .O(gate151inter4));
  nand2 gate1476(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1477(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1478(.a(G510), .O(gate151inter7));
  inv1  gate1479(.a(G513), .O(gate151inter8));
  nand2 gate1480(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1481(.a(s_133), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1482(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1483(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1484(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1919(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1920(.a(gate156inter0), .b(s_196), .O(gate156inter1));
  and2  gate1921(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1922(.a(s_196), .O(gate156inter3));
  inv1  gate1923(.a(s_197), .O(gate156inter4));
  nand2 gate1924(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1925(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1926(.a(G435), .O(gate156inter7));
  inv1  gate1927(.a(G525), .O(gate156inter8));
  nand2 gate1928(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1929(.a(s_197), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1930(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1931(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1932(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1905(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1906(.a(gate158inter0), .b(s_194), .O(gate158inter1));
  and2  gate1907(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1908(.a(s_194), .O(gate158inter3));
  inv1  gate1909(.a(s_195), .O(gate158inter4));
  nand2 gate1910(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1911(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1912(.a(G441), .O(gate158inter7));
  inv1  gate1913(.a(G528), .O(gate158inter8));
  nand2 gate1914(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1915(.a(s_195), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1916(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1917(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1918(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate841(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate842(.a(gate163inter0), .b(s_42), .O(gate163inter1));
  and2  gate843(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate844(.a(s_42), .O(gate163inter3));
  inv1  gate845(.a(s_43), .O(gate163inter4));
  nand2 gate846(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate847(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate848(.a(G456), .O(gate163inter7));
  inv1  gate849(.a(G537), .O(gate163inter8));
  nand2 gate850(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate851(.a(s_43), .b(gate163inter3), .O(gate163inter10));
  nor2  gate852(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate853(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate854(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1219(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1220(.a(gate165inter0), .b(s_96), .O(gate165inter1));
  and2  gate1221(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1222(.a(s_96), .O(gate165inter3));
  inv1  gate1223(.a(s_97), .O(gate165inter4));
  nand2 gate1224(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1225(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1226(.a(G462), .O(gate165inter7));
  inv1  gate1227(.a(G540), .O(gate165inter8));
  nand2 gate1228(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1229(.a(s_97), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1230(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1231(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1232(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1877(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1878(.a(gate166inter0), .b(s_190), .O(gate166inter1));
  and2  gate1879(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1880(.a(s_190), .O(gate166inter3));
  inv1  gate1881(.a(s_191), .O(gate166inter4));
  nand2 gate1882(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1883(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1884(.a(G465), .O(gate166inter7));
  inv1  gate1885(.a(G540), .O(gate166inter8));
  nand2 gate1886(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1887(.a(s_191), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1888(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1889(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1890(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1751(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1752(.a(gate167inter0), .b(s_172), .O(gate167inter1));
  and2  gate1753(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1754(.a(s_172), .O(gate167inter3));
  inv1  gate1755(.a(s_173), .O(gate167inter4));
  nand2 gate1756(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1757(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1758(.a(G468), .O(gate167inter7));
  inv1  gate1759(.a(G543), .O(gate167inter8));
  nand2 gate1760(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1761(.a(s_173), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1762(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1763(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1764(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1359(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1360(.a(gate170inter0), .b(s_116), .O(gate170inter1));
  and2  gate1361(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1362(.a(s_116), .O(gate170inter3));
  inv1  gate1363(.a(s_117), .O(gate170inter4));
  nand2 gate1364(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1365(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1366(.a(G477), .O(gate170inter7));
  inv1  gate1367(.a(G546), .O(gate170inter8));
  nand2 gate1368(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1369(.a(s_117), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1370(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1371(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1372(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1275(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1276(.a(gate171inter0), .b(s_104), .O(gate171inter1));
  and2  gate1277(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1278(.a(s_104), .O(gate171inter3));
  inv1  gate1279(.a(s_105), .O(gate171inter4));
  nand2 gate1280(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1281(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1282(.a(G480), .O(gate171inter7));
  inv1  gate1283(.a(G549), .O(gate171inter8));
  nand2 gate1284(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1285(.a(s_105), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1286(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1287(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1288(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1079(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1080(.a(gate173inter0), .b(s_76), .O(gate173inter1));
  and2  gate1081(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1082(.a(s_76), .O(gate173inter3));
  inv1  gate1083(.a(s_77), .O(gate173inter4));
  nand2 gate1084(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1085(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1086(.a(G486), .O(gate173inter7));
  inv1  gate1087(.a(G552), .O(gate173inter8));
  nand2 gate1088(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1089(.a(s_77), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1090(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1091(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1092(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate995(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate996(.a(gate175inter0), .b(s_64), .O(gate175inter1));
  and2  gate997(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate998(.a(s_64), .O(gate175inter3));
  inv1  gate999(.a(s_65), .O(gate175inter4));
  nand2 gate1000(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1001(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1002(.a(G492), .O(gate175inter7));
  inv1  gate1003(.a(G555), .O(gate175inter8));
  nand2 gate1004(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1005(.a(s_65), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1006(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1007(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1008(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate631(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate632(.a(gate177inter0), .b(s_12), .O(gate177inter1));
  and2  gate633(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate634(.a(s_12), .O(gate177inter3));
  inv1  gate635(.a(s_13), .O(gate177inter4));
  nand2 gate636(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate637(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate638(.a(G498), .O(gate177inter7));
  inv1  gate639(.a(G558), .O(gate177inter8));
  nand2 gate640(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate641(.a(s_13), .b(gate177inter3), .O(gate177inter10));
  nor2  gate642(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate643(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate644(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1023(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1024(.a(gate182inter0), .b(s_68), .O(gate182inter1));
  and2  gate1025(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1026(.a(s_68), .O(gate182inter3));
  inv1  gate1027(.a(s_69), .O(gate182inter4));
  nand2 gate1028(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1029(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1030(.a(G513), .O(gate182inter7));
  inv1  gate1031(.a(G564), .O(gate182inter8));
  nand2 gate1032(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1033(.a(s_69), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1034(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1035(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1036(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate925(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate926(.a(gate184inter0), .b(s_54), .O(gate184inter1));
  and2  gate927(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate928(.a(s_54), .O(gate184inter3));
  inv1  gate929(.a(s_55), .O(gate184inter4));
  nand2 gate930(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate931(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate932(.a(G519), .O(gate184inter7));
  inv1  gate933(.a(G567), .O(gate184inter8));
  nand2 gate934(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate935(.a(s_55), .b(gate184inter3), .O(gate184inter10));
  nor2  gate936(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate937(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate938(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1415(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1416(.a(gate188inter0), .b(s_124), .O(gate188inter1));
  and2  gate1417(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1418(.a(s_124), .O(gate188inter3));
  inv1  gate1419(.a(s_125), .O(gate188inter4));
  nand2 gate1420(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1421(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1422(.a(G576), .O(gate188inter7));
  inv1  gate1423(.a(G577), .O(gate188inter8));
  nand2 gate1424(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1425(.a(s_125), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1426(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1427(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1428(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1863(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1864(.a(gate191inter0), .b(s_188), .O(gate191inter1));
  and2  gate1865(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1866(.a(s_188), .O(gate191inter3));
  inv1  gate1867(.a(s_189), .O(gate191inter4));
  nand2 gate1868(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1869(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1870(.a(G582), .O(gate191inter7));
  inv1  gate1871(.a(G583), .O(gate191inter8));
  nand2 gate1872(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1873(.a(s_189), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1874(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1875(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1876(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1933(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1934(.a(gate194inter0), .b(s_198), .O(gate194inter1));
  and2  gate1935(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1936(.a(s_198), .O(gate194inter3));
  inv1  gate1937(.a(s_199), .O(gate194inter4));
  nand2 gate1938(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1939(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1940(.a(G588), .O(gate194inter7));
  inv1  gate1941(.a(G589), .O(gate194inter8));
  nand2 gate1942(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1943(.a(s_199), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1944(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1945(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1946(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate785(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate786(.a(gate195inter0), .b(s_34), .O(gate195inter1));
  and2  gate787(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate788(.a(s_34), .O(gate195inter3));
  inv1  gate789(.a(s_35), .O(gate195inter4));
  nand2 gate790(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate791(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate792(.a(G590), .O(gate195inter7));
  inv1  gate793(.a(G591), .O(gate195inter8));
  nand2 gate794(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate795(.a(s_35), .b(gate195inter3), .O(gate195inter10));
  nor2  gate796(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate797(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate798(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1429(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1430(.a(gate205inter0), .b(s_126), .O(gate205inter1));
  and2  gate1431(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1432(.a(s_126), .O(gate205inter3));
  inv1  gate1433(.a(s_127), .O(gate205inter4));
  nand2 gate1434(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1435(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1436(.a(G622), .O(gate205inter7));
  inv1  gate1437(.a(G627), .O(gate205inter8));
  nand2 gate1438(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1439(.a(s_127), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1440(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1441(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1442(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1345(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1346(.a(gate226inter0), .b(s_114), .O(gate226inter1));
  and2  gate1347(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1348(.a(s_114), .O(gate226inter3));
  inv1  gate1349(.a(s_115), .O(gate226inter4));
  nand2 gate1350(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1351(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1352(.a(G692), .O(gate226inter7));
  inv1  gate1353(.a(G693), .O(gate226inter8));
  nand2 gate1354(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1355(.a(s_115), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1356(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1357(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1358(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1695(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1696(.a(gate230inter0), .b(s_164), .O(gate230inter1));
  and2  gate1697(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1698(.a(s_164), .O(gate230inter3));
  inv1  gate1699(.a(s_165), .O(gate230inter4));
  nand2 gate1700(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1701(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1702(.a(G700), .O(gate230inter7));
  inv1  gate1703(.a(G701), .O(gate230inter8));
  nand2 gate1704(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1705(.a(s_165), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1706(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1707(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1708(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1233(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1234(.a(gate233inter0), .b(s_98), .O(gate233inter1));
  and2  gate1235(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1236(.a(s_98), .O(gate233inter3));
  inv1  gate1237(.a(s_99), .O(gate233inter4));
  nand2 gate1238(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1239(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1240(.a(G242), .O(gate233inter7));
  inv1  gate1241(.a(G718), .O(gate233inter8));
  nand2 gate1242(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1243(.a(s_99), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1244(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1245(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1246(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1149(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1150(.a(gate236inter0), .b(s_86), .O(gate236inter1));
  and2  gate1151(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1152(.a(s_86), .O(gate236inter3));
  inv1  gate1153(.a(s_87), .O(gate236inter4));
  nand2 gate1154(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1155(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1156(.a(G251), .O(gate236inter7));
  inv1  gate1157(.a(G727), .O(gate236inter8));
  nand2 gate1158(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1159(.a(s_87), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1160(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1161(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1162(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate897(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate898(.a(gate247inter0), .b(s_50), .O(gate247inter1));
  and2  gate899(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate900(.a(s_50), .O(gate247inter3));
  inv1  gate901(.a(s_51), .O(gate247inter4));
  nand2 gate902(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate903(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate904(.a(G251), .O(gate247inter7));
  inv1  gate905(.a(G739), .O(gate247inter8));
  nand2 gate906(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate907(.a(s_51), .b(gate247inter3), .O(gate247inter10));
  nor2  gate908(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate909(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate910(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate547(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate548(.a(gate250inter0), .b(s_0), .O(gate250inter1));
  and2  gate549(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate550(.a(s_0), .O(gate250inter3));
  inv1  gate551(.a(s_1), .O(gate250inter4));
  nand2 gate552(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate553(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate554(.a(G706), .O(gate250inter7));
  inv1  gate555(.a(G742), .O(gate250inter8));
  nand2 gate556(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate557(.a(s_1), .b(gate250inter3), .O(gate250inter10));
  nor2  gate558(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate559(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate560(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1387(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1388(.a(gate252inter0), .b(s_120), .O(gate252inter1));
  and2  gate1389(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1390(.a(s_120), .O(gate252inter3));
  inv1  gate1391(.a(s_121), .O(gate252inter4));
  nand2 gate1392(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1393(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1394(.a(G709), .O(gate252inter7));
  inv1  gate1395(.a(G745), .O(gate252inter8));
  nand2 gate1396(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1397(.a(s_121), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1398(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1399(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1400(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate687(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate688(.a(gate254inter0), .b(s_20), .O(gate254inter1));
  and2  gate689(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate690(.a(s_20), .O(gate254inter3));
  inv1  gate691(.a(s_21), .O(gate254inter4));
  nand2 gate692(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate693(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate694(.a(G712), .O(gate254inter7));
  inv1  gate695(.a(G748), .O(gate254inter8));
  nand2 gate696(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate697(.a(s_21), .b(gate254inter3), .O(gate254inter10));
  nor2  gate698(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate699(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate700(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1261(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1262(.a(gate256inter0), .b(s_102), .O(gate256inter1));
  and2  gate1263(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1264(.a(s_102), .O(gate256inter3));
  inv1  gate1265(.a(s_103), .O(gate256inter4));
  nand2 gate1266(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1267(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1268(.a(G715), .O(gate256inter7));
  inv1  gate1269(.a(G751), .O(gate256inter8));
  nand2 gate1270(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1271(.a(s_103), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1272(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1273(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1274(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1667(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1668(.a(gate262inter0), .b(s_160), .O(gate262inter1));
  and2  gate1669(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1670(.a(s_160), .O(gate262inter3));
  inv1  gate1671(.a(s_161), .O(gate262inter4));
  nand2 gate1672(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1673(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1674(.a(G764), .O(gate262inter7));
  inv1  gate1675(.a(G765), .O(gate262inter8));
  nand2 gate1676(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1677(.a(s_161), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1678(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1679(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1680(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate911(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate912(.a(gate265inter0), .b(s_52), .O(gate265inter1));
  and2  gate913(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate914(.a(s_52), .O(gate265inter3));
  inv1  gate915(.a(s_53), .O(gate265inter4));
  nand2 gate916(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate917(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate918(.a(G642), .O(gate265inter7));
  inv1  gate919(.a(G770), .O(gate265inter8));
  nand2 gate920(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate921(.a(s_53), .b(gate265inter3), .O(gate265inter10));
  nor2  gate922(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate923(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate924(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1065(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1066(.a(gate267inter0), .b(s_74), .O(gate267inter1));
  and2  gate1067(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1068(.a(s_74), .O(gate267inter3));
  inv1  gate1069(.a(s_75), .O(gate267inter4));
  nand2 gate1070(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1071(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1072(.a(G648), .O(gate267inter7));
  inv1  gate1073(.a(G776), .O(gate267inter8));
  nand2 gate1074(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1075(.a(s_75), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1076(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1077(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1078(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1205(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1206(.a(gate270inter0), .b(s_94), .O(gate270inter1));
  and2  gate1207(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1208(.a(s_94), .O(gate270inter3));
  inv1  gate1209(.a(s_95), .O(gate270inter4));
  nand2 gate1210(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1211(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1212(.a(G657), .O(gate270inter7));
  inv1  gate1213(.a(G785), .O(gate270inter8));
  nand2 gate1214(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1215(.a(s_95), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1216(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1217(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1218(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1793(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1794(.a(gate272inter0), .b(s_178), .O(gate272inter1));
  and2  gate1795(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1796(.a(s_178), .O(gate272inter3));
  inv1  gate1797(.a(s_179), .O(gate272inter4));
  nand2 gate1798(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1799(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1800(.a(G663), .O(gate272inter7));
  inv1  gate1801(.a(G791), .O(gate272inter8));
  nand2 gate1802(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1803(.a(s_179), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1804(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1805(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1806(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1485(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1486(.a(gate273inter0), .b(s_134), .O(gate273inter1));
  and2  gate1487(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1488(.a(s_134), .O(gate273inter3));
  inv1  gate1489(.a(s_135), .O(gate273inter4));
  nand2 gate1490(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1491(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1492(.a(G642), .O(gate273inter7));
  inv1  gate1493(.a(G794), .O(gate273inter8));
  nand2 gate1494(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1495(.a(s_135), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1496(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1497(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1498(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1303(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1304(.a(gate283inter0), .b(s_108), .O(gate283inter1));
  and2  gate1305(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1306(.a(s_108), .O(gate283inter3));
  inv1  gate1307(.a(s_109), .O(gate283inter4));
  nand2 gate1308(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1309(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1310(.a(G657), .O(gate283inter7));
  inv1  gate1311(.a(G809), .O(gate283inter8));
  nand2 gate1312(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1313(.a(s_109), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1314(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1315(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1316(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1555(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1556(.a(gate286inter0), .b(s_144), .O(gate286inter1));
  and2  gate1557(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1558(.a(s_144), .O(gate286inter3));
  inv1  gate1559(.a(s_145), .O(gate286inter4));
  nand2 gate1560(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1561(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1562(.a(G788), .O(gate286inter7));
  inv1  gate1563(.a(G812), .O(gate286inter8));
  nand2 gate1564(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1565(.a(s_145), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1566(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1567(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1568(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1625(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1626(.a(gate296inter0), .b(s_154), .O(gate296inter1));
  and2  gate1627(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1628(.a(s_154), .O(gate296inter3));
  inv1  gate1629(.a(s_155), .O(gate296inter4));
  nand2 gate1630(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1631(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1632(.a(G826), .O(gate296inter7));
  inv1  gate1633(.a(G827), .O(gate296inter8));
  nand2 gate1634(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1635(.a(s_155), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1636(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1637(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1638(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate967(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate968(.a(gate390inter0), .b(s_60), .O(gate390inter1));
  and2  gate969(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate970(.a(s_60), .O(gate390inter3));
  inv1  gate971(.a(s_61), .O(gate390inter4));
  nand2 gate972(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate973(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate974(.a(G4), .O(gate390inter7));
  inv1  gate975(.a(G1045), .O(gate390inter8));
  nand2 gate976(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate977(.a(s_61), .b(gate390inter3), .O(gate390inter10));
  nor2  gate978(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate979(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate980(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1331(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1332(.a(gate397inter0), .b(s_112), .O(gate397inter1));
  and2  gate1333(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1334(.a(s_112), .O(gate397inter3));
  inv1  gate1335(.a(s_113), .O(gate397inter4));
  nand2 gate1336(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1337(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1338(.a(G11), .O(gate397inter7));
  inv1  gate1339(.a(G1066), .O(gate397inter8));
  nand2 gate1340(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1341(.a(s_113), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1342(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1343(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1344(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1289(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1290(.a(gate406inter0), .b(s_106), .O(gate406inter1));
  and2  gate1291(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1292(.a(s_106), .O(gate406inter3));
  inv1  gate1293(.a(s_107), .O(gate406inter4));
  nand2 gate1294(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1295(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1296(.a(G20), .O(gate406inter7));
  inv1  gate1297(.a(G1093), .O(gate406inter8));
  nand2 gate1298(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1299(.a(s_107), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1300(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1301(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1302(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1443(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1444(.a(gate415inter0), .b(s_128), .O(gate415inter1));
  and2  gate1445(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1446(.a(s_128), .O(gate415inter3));
  inv1  gate1447(.a(s_129), .O(gate415inter4));
  nand2 gate1448(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1449(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1450(.a(G29), .O(gate415inter7));
  inv1  gate1451(.a(G1120), .O(gate415inter8));
  nand2 gate1452(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1453(.a(s_129), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1454(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1455(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1456(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate673(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate674(.a(gate420inter0), .b(s_18), .O(gate420inter1));
  and2  gate675(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate676(.a(s_18), .O(gate420inter3));
  inv1  gate677(.a(s_19), .O(gate420inter4));
  nand2 gate678(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate679(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate680(.a(G1036), .O(gate420inter7));
  inv1  gate681(.a(G1132), .O(gate420inter8));
  nand2 gate682(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate683(.a(s_19), .b(gate420inter3), .O(gate420inter10));
  nor2  gate684(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate685(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate686(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate827(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate828(.a(gate423inter0), .b(s_40), .O(gate423inter1));
  and2  gate829(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate830(.a(s_40), .O(gate423inter3));
  inv1  gate831(.a(s_41), .O(gate423inter4));
  nand2 gate832(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate833(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate834(.a(G3), .O(gate423inter7));
  inv1  gate835(.a(G1138), .O(gate423inter8));
  nand2 gate836(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate837(.a(s_41), .b(gate423inter3), .O(gate423inter10));
  nor2  gate838(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate839(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate840(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1821(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1822(.a(gate431inter0), .b(s_182), .O(gate431inter1));
  and2  gate1823(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1824(.a(s_182), .O(gate431inter3));
  inv1  gate1825(.a(s_183), .O(gate431inter4));
  nand2 gate1826(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1827(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1828(.a(G7), .O(gate431inter7));
  inv1  gate1829(.a(G1150), .O(gate431inter8));
  nand2 gate1830(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1831(.a(s_183), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1832(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1833(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1834(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1639(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1640(.a(gate435inter0), .b(s_156), .O(gate435inter1));
  and2  gate1641(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1642(.a(s_156), .O(gate435inter3));
  inv1  gate1643(.a(s_157), .O(gate435inter4));
  nand2 gate1644(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1645(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1646(.a(G9), .O(gate435inter7));
  inv1  gate1647(.a(G1156), .O(gate435inter8));
  nand2 gate1648(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1649(.a(s_157), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1650(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1651(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1652(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate883(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate884(.a(gate440inter0), .b(s_48), .O(gate440inter1));
  and2  gate885(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate886(.a(s_48), .O(gate440inter3));
  inv1  gate887(.a(s_49), .O(gate440inter4));
  nand2 gate888(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate889(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate890(.a(G1066), .O(gate440inter7));
  inv1  gate891(.a(G1162), .O(gate440inter8));
  nand2 gate892(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate893(.a(s_49), .b(gate440inter3), .O(gate440inter10));
  nor2  gate894(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate895(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate896(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1597(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1598(.a(gate443inter0), .b(s_150), .O(gate443inter1));
  and2  gate1599(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1600(.a(s_150), .O(gate443inter3));
  inv1  gate1601(.a(s_151), .O(gate443inter4));
  nand2 gate1602(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1603(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1604(.a(G13), .O(gate443inter7));
  inv1  gate1605(.a(G1168), .O(gate443inter8));
  nand2 gate1606(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1607(.a(s_151), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1608(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1609(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1610(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1891(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1892(.a(gate444inter0), .b(s_192), .O(gate444inter1));
  and2  gate1893(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1894(.a(s_192), .O(gate444inter3));
  inv1  gate1895(.a(s_193), .O(gate444inter4));
  nand2 gate1896(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1897(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1898(.a(G1072), .O(gate444inter7));
  inv1  gate1899(.a(G1168), .O(gate444inter8));
  nand2 gate1900(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1901(.a(s_193), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1902(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1903(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1904(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1611(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1612(.a(gate448inter0), .b(s_152), .O(gate448inter1));
  and2  gate1613(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1614(.a(s_152), .O(gate448inter3));
  inv1  gate1615(.a(s_153), .O(gate448inter4));
  nand2 gate1616(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1617(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1618(.a(G1078), .O(gate448inter7));
  inv1  gate1619(.a(G1174), .O(gate448inter8));
  nand2 gate1620(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1621(.a(s_153), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1622(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1623(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1624(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1947(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1948(.a(gate458inter0), .b(s_200), .O(gate458inter1));
  and2  gate1949(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1950(.a(s_200), .O(gate458inter3));
  inv1  gate1951(.a(s_201), .O(gate458inter4));
  nand2 gate1952(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1953(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1954(.a(G1093), .O(gate458inter7));
  inv1  gate1955(.a(G1189), .O(gate458inter8));
  nand2 gate1956(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1957(.a(s_201), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1958(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1959(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1960(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1737(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1738(.a(gate460inter0), .b(s_170), .O(gate460inter1));
  and2  gate1739(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1740(.a(s_170), .O(gate460inter3));
  inv1  gate1741(.a(s_171), .O(gate460inter4));
  nand2 gate1742(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1743(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1744(.a(G1096), .O(gate460inter7));
  inv1  gate1745(.a(G1192), .O(gate460inter8));
  nand2 gate1746(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1747(.a(s_171), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1748(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1749(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1750(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate561(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate562(.a(gate462inter0), .b(s_2), .O(gate462inter1));
  and2  gate563(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate564(.a(s_2), .O(gate462inter3));
  inv1  gate565(.a(s_3), .O(gate462inter4));
  nand2 gate566(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate567(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate568(.a(G1099), .O(gate462inter7));
  inv1  gate569(.a(G1195), .O(gate462inter8));
  nand2 gate570(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate571(.a(s_3), .b(gate462inter3), .O(gate462inter10));
  nor2  gate572(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate573(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate574(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1009(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1010(.a(gate463inter0), .b(s_66), .O(gate463inter1));
  and2  gate1011(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1012(.a(s_66), .O(gate463inter3));
  inv1  gate1013(.a(s_67), .O(gate463inter4));
  nand2 gate1014(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1015(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1016(.a(G23), .O(gate463inter7));
  inv1  gate1017(.a(G1198), .O(gate463inter8));
  nand2 gate1018(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1019(.a(s_67), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1020(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1021(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1022(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1807(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1808(.a(gate464inter0), .b(s_180), .O(gate464inter1));
  and2  gate1809(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1810(.a(s_180), .O(gate464inter3));
  inv1  gate1811(.a(s_181), .O(gate464inter4));
  nand2 gate1812(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1813(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1814(.a(G1102), .O(gate464inter7));
  inv1  gate1815(.a(G1198), .O(gate464inter8));
  nand2 gate1816(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1817(.a(s_181), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1818(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1819(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1820(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate743(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate744(.a(gate467inter0), .b(s_28), .O(gate467inter1));
  and2  gate745(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate746(.a(s_28), .O(gate467inter3));
  inv1  gate747(.a(s_29), .O(gate467inter4));
  nand2 gate748(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate749(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate750(.a(G25), .O(gate467inter7));
  inv1  gate751(.a(G1204), .O(gate467inter8));
  nand2 gate752(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate753(.a(s_29), .b(gate467inter3), .O(gate467inter10));
  nor2  gate754(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate755(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate756(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1401(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1402(.a(gate469inter0), .b(s_122), .O(gate469inter1));
  and2  gate1403(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1404(.a(s_122), .O(gate469inter3));
  inv1  gate1405(.a(s_123), .O(gate469inter4));
  nand2 gate1406(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1407(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1408(.a(G26), .O(gate469inter7));
  inv1  gate1409(.a(G1207), .O(gate469inter8));
  nand2 gate1410(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1411(.a(s_123), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1412(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1413(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1414(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate603(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate604(.a(gate470inter0), .b(s_8), .O(gate470inter1));
  and2  gate605(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate606(.a(s_8), .O(gate470inter3));
  inv1  gate607(.a(s_9), .O(gate470inter4));
  nand2 gate608(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate609(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate610(.a(G1111), .O(gate470inter7));
  inv1  gate611(.a(G1207), .O(gate470inter8));
  nand2 gate612(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate613(.a(s_9), .b(gate470inter3), .O(gate470inter10));
  nor2  gate614(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate615(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate616(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate589(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate590(.a(gate476inter0), .b(s_6), .O(gate476inter1));
  and2  gate591(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate592(.a(s_6), .O(gate476inter3));
  inv1  gate593(.a(s_7), .O(gate476inter4));
  nand2 gate594(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate595(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate596(.a(G1120), .O(gate476inter7));
  inv1  gate597(.a(G1216), .O(gate476inter8));
  nand2 gate598(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate599(.a(s_7), .b(gate476inter3), .O(gate476inter10));
  nor2  gate600(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate601(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate602(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1765(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1766(.a(gate477inter0), .b(s_174), .O(gate477inter1));
  and2  gate1767(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1768(.a(s_174), .O(gate477inter3));
  inv1  gate1769(.a(s_175), .O(gate477inter4));
  nand2 gate1770(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1771(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1772(.a(G30), .O(gate477inter7));
  inv1  gate1773(.a(G1219), .O(gate477inter8));
  nand2 gate1774(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1775(.a(s_175), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1776(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1777(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1778(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate799(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate800(.a(gate482inter0), .b(s_36), .O(gate482inter1));
  and2  gate801(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate802(.a(s_36), .O(gate482inter3));
  inv1  gate803(.a(s_37), .O(gate482inter4));
  nand2 gate804(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate805(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate806(.a(G1129), .O(gate482inter7));
  inv1  gate807(.a(G1225), .O(gate482inter8));
  nand2 gate808(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate809(.a(s_37), .b(gate482inter3), .O(gate482inter10));
  nor2  gate810(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate811(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate812(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate939(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate940(.a(gate489inter0), .b(s_56), .O(gate489inter1));
  and2  gate941(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate942(.a(s_56), .O(gate489inter3));
  inv1  gate943(.a(s_57), .O(gate489inter4));
  nand2 gate944(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate945(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate946(.a(G1240), .O(gate489inter7));
  inv1  gate947(.a(G1241), .O(gate489inter8));
  nand2 gate948(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate949(.a(s_57), .b(gate489inter3), .O(gate489inter10));
  nor2  gate950(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate951(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate952(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate617(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate618(.a(gate491inter0), .b(s_10), .O(gate491inter1));
  and2  gate619(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate620(.a(s_10), .O(gate491inter3));
  inv1  gate621(.a(s_11), .O(gate491inter4));
  nand2 gate622(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate623(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate624(.a(G1244), .O(gate491inter7));
  inv1  gate625(.a(G1245), .O(gate491inter8));
  nand2 gate626(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate627(.a(s_11), .b(gate491inter3), .O(gate491inter10));
  nor2  gate628(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate629(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate630(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate855(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate856(.a(gate493inter0), .b(s_44), .O(gate493inter1));
  and2  gate857(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate858(.a(s_44), .O(gate493inter3));
  inv1  gate859(.a(s_45), .O(gate493inter4));
  nand2 gate860(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate861(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate862(.a(G1248), .O(gate493inter7));
  inv1  gate863(.a(G1249), .O(gate493inter8));
  nand2 gate864(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate865(.a(s_45), .b(gate493inter3), .O(gate493inter10));
  nor2  gate866(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate867(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate868(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1513(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1514(.a(gate497inter0), .b(s_138), .O(gate497inter1));
  and2  gate1515(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1516(.a(s_138), .O(gate497inter3));
  inv1  gate1517(.a(s_139), .O(gate497inter4));
  nand2 gate1518(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1519(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1520(.a(G1256), .O(gate497inter7));
  inv1  gate1521(.a(G1257), .O(gate497inter8));
  nand2 gate1522(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1523(.a(s_139), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1524(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1525(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1526(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate659(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate660(.a(gate499inter0), .b(s_16), .O(gate499inter1));
  and2  gate661(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate662(.a(s_16), .O(gate499inter3));
  inv1  gate663(.a(s_17), .O(gate499inter4));
  nand2 gate664(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate665(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate666(.a(G1260), .O(gate499inter7));
  inv1  gate667(.a(G1261), .O(gate499inter8));
  nand2 gate668(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate669(.a(s_17), .b(gate499inter3), .O(gate499inter10));
  nor2  gate670(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate671(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate672(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate729(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate730(.a(gate500inter0), .b(s_26), .O(gate500inter1));
  and2  gate731(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate732(.a(s_26), .O(gate500inter3));
  inv1  gate733(.a(s_27), .O(gate500inter4));
  nand2 gate734(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate735(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate736(.a(G1262), .O(gate500inter7));
  inv1  gate737(.a(G1263), .O(gate500inter8));
  nand2 gate738(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate739(.a(s_27), .b(gate500inter3), .O(gate500inter10));
  nor2  gate740(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate741(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate742(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate575(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate576(.a(gate501inter0), .b(s_4), .O(gate501inter1));
  and2  gate577(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate578(.a(s_4), .O(gate501inter3));
  inv1  gate579(.a(s_5), .O(gate501inter4));
  nand2 gate580(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate581(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate582(.a(G1264), .O(gate501inter7));
  inv1  gate583(.a(G1265), .O(gate501inter8));
  nand2 gate584(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate585(.a(s_5), .b(gate501inter3), .O(gate501inter10));
  nor2  gate586(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate587(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate588(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1569(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1570(.a(gate502inter0), .b(s_146), .O(gate502inter1));
  and2  gate1571(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1572(.a(s_146), .O(gate502inter3));
  inv1  gate1573(.a(s_147), .O(gate502inter4));
  nand2 gate1574(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1575(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1576(.a(G1266), .O(gate502inter7));
  inv1  gate1577(.a(G1267), .O(gate502inter8));
  nand2 gate1578(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1579(.a(s_147), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1580(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1581(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1582(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1317(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1318(.a(gate506inter0), .b(s_110), .O(gate506inter1));
  and2  gate1319(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1320(.a(s_110), .O(gate506inter3));
  inv1  gate1321(.a(s_111), .O(gate506inter4));
  nand2 gate1322(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1323(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1324(.a(G1274), .O(gate506inter7));
  inv1  gate1325(.a(G1275), .O(gate506inter8));
  nand2 gate1326(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1327(.a(s_111), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1328(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1329(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1330(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1163(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1164(.a(gate510inter0), .b(s_88), .O(gate510inter1));
  and2  gate1165(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1166(.a(s_88), .O(gate510inter3));
  inv1  gate1167(.a(s_89), .O(gate510inter4));
  nand2 gate1168(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1169(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1170(.a(G1282), .O(gate510inter7));
  inv1  gate1171(.a(G1283), .O(gate510inter8));
  nand2 gate1172(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1173(.a(s_89), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1174(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1175(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1176(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule