module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
input s_382,s_383;//RE__ALLOW(00,01,10,11);
input s_384,s_385;//RE__ALLOW(00,01,10,11);
input s_386,s_387;//RE__ALLOW(00,01,10,11);
input s_388,s_389;//RE__ALLOW(00,01,10,11);
input s_390,s_391;//RE__ALLOW(00,01,10,11);
input s_392,s_393;//RE__ALLOW(00,01,10,11);
input s_394,s_395;//RE__ALLOW(00,01,10,11);
input s_396,s_397;//RE__ALLOW(00,01,10,11);
input s_398,s_399;//RE__ALLOW(00,01,10,11);
input s_400,s_401;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2395(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2396(.a(gate10inter0), .b(s_264), .O(gate10inter1));
  and2  gate2397(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2398(.a(s_264), .O(gate10inter3));
  inv1  gate2399(.a(s_265), .O(gate10inter4));
  nand2 gate2400(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2401(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2402(.a(G3), .O(gate10inter7));
  inv1  gate2403(.a(G4), .O(gate10inter8));
  nand2 gate2404(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2405(.a(s_265), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2406(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2407(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2408(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2311(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2312(.a(gate14inter0), .b(s_252), .O(gate14inter1));
  and2  gate2313(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2314(.a(s_252), .O(gate14inter3));
  inv1  gate2315(.a(s_253), .O(gate14inter4));
  nand2 gate2316(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2317(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2318(.a(G11), .O(gate14inter7));
  inv1  gate2319(.a(G12), .O(gate14inter8));
  nand2 gate2320(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2321(.a(s_253), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2322(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2323(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2324(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2031(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2032(.a(gate16inter0), .b(s_212), .O(gate16inter1));
  and2  gate2033(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2034(.a(s_212), .O(gate16inter3));
  inv1  gate2035(.a(s_213), .O(gate16inter4));
  nand2 gate2036(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2037(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2038(.a(G15), .O(gate16inter7));
  inv1  gate2039(.a(G16), .O(gate16inter8));
  nand2 gate2040(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2041(.a(s_213), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2042(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2043(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2044(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2829(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2830(.a(gate17inter0), .b(s_326), .O(gate17inter1));
  and2  gate2831(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2832(.a(s_326), .O(gate17inter3));
  inv1  gate2833(.a(s_327), .O(gate17inter4));
  nand2 gate2834(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2835(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2836(.a(G17), .O(gate17inter7));
  inv1  gate2837(.a(G18), .O(gate17inter8));
  nand2 gate2838(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2839(.a(s_327), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2840(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2841(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2842(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate2815(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2816(.a(gate18inter0), .b(s_324), .O(gate18inter1));
  and2  gate2817(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2818(.a(s_324), .O(gate18inter3));
  inv1  gate2819(.a(s_325), .O(gate18inter4));
  nand2 gate2820(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2821(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2822(.a(G19), .O(gate18inter7));
  inv1  gate2823(.a(G20), .O(gate18inter8));
  nand2 gate2824(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2825(.a(s_325), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2826(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2827(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2828(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2059(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2060(.a(gate19inter0), .b(s_216), .O(gate19inter1));
  and2  gate2061(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2062(.a(s_216), .O(gate19inter3));
  inv1  gate2063(.a(s_217), .O(gate19inter4));
  nand2 gate2064(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2065(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2066(.a(G21), .O(gate19inter7));
  inv1  gate2067(.a(G22), .O(gate19inter8));
  nand2 gate2068(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2069(.a(s_217), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2070(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2071(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2072(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2661(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2662(.a(gate20inter0), .b(s_302), .O(gate20inter1));
  and2  gate2663(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2664(.a(s_302), .O(gate20inter3));
  inv1  gate2665(.a(s_303), .O(gate20inter4));
  nand2 gate2666(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2667(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2668(.a(G23), .O(gate20inter7));
  inv1  gate2669(.a(G24), .O(gate20inter8));
  nand2 gate2670(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2671(.a(s_303), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2672(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2673(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2674(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1583(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1584(.a(gate21inter0), .b(s_148), .O(gate21inter1));
  and2  gate1585(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1586(.a(s_148), .O(gate21inter3));
  inv1  gate1587(.a(s_149), .O(gate21inter4));
  nand2 gate1588(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1589(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1590(.a(G25), .O(gate21inter7));
  inv1  gate1591(.a(G26), .O(gate21inter8));
  nand2 gate1592(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1593(.a(s_149), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1594(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1595(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1596(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2731(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2732(.a(gate24inter0), .b(s_312), .O(gate24inter1));
  and2  gate2733(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2734(.a(s_312), .O(gate24inter3));
  inv1  gate2735(.a(s_313), .O(gate24inter4));
  nand2 gate2736(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2737(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2738(.a(G31), .O(gate24inter7));
  inv1  gate2739(.a(G32), .O(gate24inter8));
  nand2 gate2740(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2741(.a(s_313), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2742(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2743(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2744(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2899(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2900(.a(gate26inter0), .b(s_336), .O(gate26inter1));
  and2  gate2901(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2902(.a(s_336), .O(gate26inter3));
  inv1  gate2903(.a(s_337), .O(gate26inter4));
  nand2 gate2904(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2905(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2906(.a(G9), .O(gate26inter7));
  inv1  gate2907(.a(G13), .O(gate26inter8));
  nand2 gate2908(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2909(.a(s_337), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2910(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2911(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2912(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate2171(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2172(.a(gate27inter0), .b(s_232), .O(gate27inter1));
  and2  gate2173(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2174(.a(s_232), .O(gate27inter3));
  inv1  gate2175(.a(s_233), .O(gate27inter4));
  nand2 gate2176(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2177(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2178(.a(G2), .O(gate27inter7));
  inv1  gate2179(.a(G6), .O(gate27inter8));
  nand2 gate2180(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2181(.a(s_233), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2182(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2183(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2184(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate2017(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2018(.a(gate28inter0), .b(s_210), .O(gate28inter1));
  and2  gate2019(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2020(.a(s_210), .O(gate28inter3));
  inv1  gate2021(.a(s_211), .O(gate28inter4));
  nand2 gate2022(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2023(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2024(.a(G10), .O(gate28inter7));
  inv1  gate2025(.a(G14), .O(gate28inter8));
  nand2 gate2026(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2027(.a(s_211), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2028(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2029(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2030(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2941(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2942(.a(gate29inter0), .b(s_342), .O(gate29inter1));
  and2  gate2943(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2944(.a(s_342), .O(gate29inter3));
  inv1  gate2945(.a(s_343), .O(gate29inter4));
  nand2 gate2946(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2947(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2948(.a(G3), .O(gate29inter7));
  inv1  gate2949(.a(G7), .O(gate29inter8));
  nand2 gate2950(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2951(.a(s_343), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2952(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2953(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2954(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate3109(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate3110(.a(gate31inter0), .b(s_366), .O(gate31inter1));
  and2  gate3111(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate3112(.a(s_366), .O(gate31inter3));
  inv1  gate3113(.a(s_367), .O(gate31inter4));
  nand2 gate3114(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate3115(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate3116(.a(G4), .O(gate31inter7));
  inv1  gate3117(.a(G8), .O(gate31inter8));
  nand2 gate3118(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate3119(.a(s_367), .b(gate31inter3), .O(gate31inter10));
  nor2  gate3120(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate3121(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate3122(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1611(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1612(.a(gate32inter0), .b(s_152), .O(gate32inter1));
  and2  gate1613(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1614(.a(s_152), .O(gate32inter3));
  inv1  gate1615(.a(s_153), .O(gate32inter4));
  nand2 gate1616(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1617(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1618(.a(G12), .O(gate32inter7));
  inv1  gate1619(.a(G16), .O(gate32inter8));
  nand2 gate1620(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1621(.a(s_153), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1622(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1623(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1624(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate2703(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2704(.a(gate33inter0), .b(s_308), .O(gate33inter1));
  and2  gate2705(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2706(.a(s_308), .O(gate33inter3));
  inv1  gate2707(.a(s_309), .O(gate33inter4));
  nand2 gate2708(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2709(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2710(.a(G17), .O(gate33inter7));
  inv1  gate2711(.a(G21), .O(gate33inter8));
  nand2 gate2712(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2713(.a(s_309), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2714(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2715(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2716(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1443(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1444(.a(gate34inter0), .b(s_128), .O(gate34inter1));
  and2  gate1445(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1446(.a(s_128), .O(gate34inter3));
  inv1  gate1447(.a(s_129), .O(gate34inter4));
  nand2 gate1448(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1449(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1450(.a(G25), .O(gate34inter7));
  inv1  gate1451(.a(G29), .O(gate34inter8));
  nand2 gate1452(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1453(.a(s_129), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1454(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1455(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1456(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1849(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1850(.a(gate35inter0), .b(s_186), .O(gate35inter1));
  and2  gate1851(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1852(.a(s_186), .O(gate35inter3));
  inv1  gate1853(.a(s_187), .O(gate35inter4));
  nand2 gate1854(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1855(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1856(.a(G18), .O(gate35inter7));
  inv1  gate1857(.a(G22), .O(gate35inter8));
  nand2 gate1858(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1859(.a(s_187), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1860(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1861(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1862(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2773(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2774(.a(gate40inter0), .b(s_318), .O(gate40inter1));
  and2  gate2775(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2776(.a(s_318), .O(gate40inter3));
  inv1  gate2777(.a(s_319), .O(gate40inter4));
  nand2 gate2778(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2779(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2780(.a(G28), .O(gate40inter7));
  inv1  gate2781(.a(G32), .O(gate40inter8));
  nand2 gate2782(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2783(.a(s_319), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2784(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2785(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2786(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2549(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2550(.a(gate46inter0), .b(s_286), .O(gate46inter1));
  and2  gate2551(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2552(.a(s_286), .O(gate46inter3));
  inv1  gate2553(.a(s_287), .O(gate46inter4));
  nand2 gate2554(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2555(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2556(.a(G6), .O(gate46inter7));
  inv1  gate2557(.a(G272), .O(gate46inter8));
  nand2 gate2558(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2559(.a(s_287), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2560(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2561(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2562(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2297(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2298(.a(gate50inter0), .b(s_250), .O(gate50inter1));
  and2  gate2299(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2300(.a(s_250), .O(gate50inter3));
  inv1  gate2301(.a(s_251), .O(gate50inter4));
  nand2 gate2302(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2303(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2304(.a(G10), .O(gate50inter7));
  inv1  gate2305(.a(G278), .O(gate50inter8));
  nand2 gate2306(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2307(.a(s_251), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2308(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2309(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2310(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1023(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1024(.a(gate52inter0), .b(s_68), .O(gate52inter1));
  and2  gate1025(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1026(.a(s_68), .O(gate52inter3));
  inv1  gate1027(.a(s_69), .O(gate52inter4));
  nand2 gate1028(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1029(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1030(.a(G12), .O(gate52inter7));
  inv1  gate1031(.a(G281), .O(gate52inter8));
  nand2 gate1032(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1033(.a(s_69), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1034(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1035(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1036(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1947(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1948(.a(gate54inter0), .b(s_200), .O(gate54inter1));
  and2  gate1949(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1950(.a(s_200), .O(gate54inter3));
  inv1  gate1951(.a(s_201), .O(gate54inter4));
  nand2 gate1952(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1953(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1954(.a(G14), .O(gate54inter7));
  inv1  gate1955(.a(G284), .O(gate54inter8));
  nand2 gate1956(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1957(.a(s_201), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1958(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1959(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1960(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2997(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2998(.a(gate56inter0), .b(s_350), .O(gate56inter1));
  and2  gate2999(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate3000(.a(s_350), .O(gate56inter3));
  inv1  gate3001(.a(s_351), .O(gate56inter4));
  nand2 gate3002(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate3003(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate3004(.a(G16), .O(gate56inter7));
  inv1  gate3005(.a(G287), .O(gate56inter8));
  nand2 gate3006(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate3007(.a(s_351), .b(gate56inter3), .O(gate56inter10));
  nor2  gate3008(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate3009(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate3010(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate3305(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate3306(.a(gate58inter0), .b(s_394), .O(gate58inter1));
  and2  gate3307(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate3308(.a(s_394), .O(gate58inter3));
  inv1  gate3309(.a(s_395), .O(gate58inter4));
  nand2 gate3310(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate3311(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate3312(.a(G18), .O(gate58inter7));
  inv1  gate3313(.a(G290), .O(gate58inter8));
  nand2 gate3314(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate3315(.a(s_395), .b(gate58inter3), .O(gate58inter10));
  nor2  gate3316(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate3317(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate3318(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate785(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate786(.a(gate59inter0), .b(s_34), .O(gate59inter1));
  and2  gate787(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate788(.a(s_34), .O(gate59inter3));
  inv1  gate789(.a(s_35), .O(gate59inter4));
  nand2 gate790(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate791(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate792(.a(G19), .O(gate59inter7));
  inv1  gate793(.a(G293), .O(gate59inter8));
  nand2 gate794(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate795(.a(s_35), .b(gate59inter3), .O(gate59inter10));
  nor2  gate796(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate797(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate798(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1359(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1360(.a(gate60inter0), .b(s_116), .O(gate60inter1));
  and2  gate1361(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1362(.a(s_116), .O(gate60inter3));
  inv1  gate1363(.a(s_117), .O(gate60inter4));
  nand2 gate1364(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1365(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1366(.a(G20), .O(gate60inter7));
  inv1  gate1367(.a(G293), .O(gate60inter8));
  nand2 gate1368(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1369(.a(s_117), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1370(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1371(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1372(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate3235(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate3236(.a(gate61inter0), .b(s_384), .O(gate61inter1));
  and2  gate3237(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate3238(.a(s_384), .O(gate61inter3));
  inv1  gate3239(.a(s_385), .O(gate61inter4));
  nand2 gate3240(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate3241(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate3242(.a(G21), .O(gate61inter7));
  inv1  gate3243(.a(G296), .O(gate61inter8));
  nand2 gate3244(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate3245(.a(s_385), .b(gate61inter3), .O(gate61inter10));
  nor2  gate3246(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate3247(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate3248(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1387(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1388(.a(gate68inter0), .b(s_120), .O(gate68inter1));
  and2  gate1389(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1390(.a(s_120), .O(gate68inter3));
  inv1  gate1391(.a(s_121), .O(gate68inter4));
  nand2 gate1392(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1393(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1394(.a(G28), .O(gate68inter7));
  inv1  gate1395(.a(G305), .O(gate68inter8));
  nand2 gate1396(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1397(.a(s_121), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1398(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1399(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1400(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate3025(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate3026(.a(gate69inter0), .b(s_354), .O(gate69inter1));
  and2  gate3027(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate3028(.a(s_354), .O(gate69inter3));
  inv1  gate3029(.a(s_355), .O(gate69inter4));
  nand2 gate3030(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate3031(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate3032(.a(G29), .O(gate69inter7));
  inv1  gate3033(.a(G308), .O(gate69inter8));
  nand2 gate3034(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate3035(.a(s_355), .b(gate69inter3), .O(gate69inter10));
  nor2  gate3036(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate3037(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate3038(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate841(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate842(.a(gate71inter0), .b(s_42), .O(gate71inter1));
  and2  gate843(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate844(.a(s_42), .O(gate71inter3));
  inv1  gate845(.a(s_43), .O(gate71inter4));
  nand2 gate846(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate847(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate848(.a(G31), .O(gate71inter7));
  inv1  gate849(.a(G311), .O(gate71inter8));
  nand2 gate850(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate851(.a(s_43), .b(gate71inter3), .O(gate71inter10));
  nor2  gate852(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate853(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate854(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate827(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate828(.a(gate73inter0), .b(s_40), .O(gate73inter1));
  and2  gate829(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate830(.a(s_40), .O(gate73inter3));
  inv1  gate831(.a(s_41), .O(gate73inter4));
  nand2 gate832(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate833(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate834(.a(G1), .O(gate73inter7));
  inv1  gate835(.a(G314), .O(gate73inter8));
  nand2 gate836(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate837(.a(s_41), .b(gate73inter3), .O(gate73inter10));
  nor2  gate838(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate839(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate840(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1695(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1696(.a(gate74inter0), .b(s_164), .O(gate74inter1));
  and2  gate1697(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1698(.a(s_164), .O(gate74inter3));
  inv1  gate1699(.a(s_165), .O(gate74inter4));
  nand2 gate1700(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1701(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1702(.a(G5), .O(gate74inter7));
  inv1  gate1703(.a(G314), .O(gate74inter8));
  nand2 gate1704(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1705(.a(s_165), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1706(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1707(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1708(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate729(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate730(.a(gate75inter0), .b(s_26), .O(gate75inter1));
  and2  gate731(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate732(.a(s_26), .O(gate75inter3));
  inv1  gate733(.a(s_27), .O(gate75inter4));
  nand2 gate734(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate735(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate736(.a(G9), .O(gate75inter7));
  inv1  gate737(.a(G317), .O(gate75inter8));
  nand2 gate738(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate739(.a(s_27), .b(gate75inter3), .O(gate75inter10));
  nor2  gate740(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate741(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate742(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1051(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1052(.a(gate77inter0), .b(s_72), .O(gate77inter1));
  and2  gate1053(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1054(.a(s_72), .O(gate77inter3));
  inv1  gate1055(.a(s_73), .O(gate77inter4));
  nand2 gate1056(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1057(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1058(.a(G2), .O(gate77inter7));
  inv1  gate1059(.a(G320), .O(gate77inter8));
  nand2 gate1060(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1061(.a(s_73), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1062(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1063(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1064(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate3053(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate3054(.a(gate78inter0), .b(s_358), .O(gate78inter1));
  and2  gate3055(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate3056(.a(s_358), .O(gate78inter3));
  inv1  gate3057(.a(s_359), .O(gate78inter4));
  nand2 gate3058(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate3059(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate3060(.a(G6), .O(gate78inter7));
  inv1  gate3061(.a(G320), .O(gate78inter8));
  nand2 gate3062(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate3063(.a(s_359), .b(gate78inter3), .O(gate78inter10));
  nor2  gate3064(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate3065(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate3066(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate925(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate926(.a(gate79inter0), .b(s_54), .O(gate79inter1));
  and2  gate927(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate928(.a(s_54), .O(gate79inter3));
  inv1  gate929(.a(s_55), .O(gate79inter4));
  nand2 gate930(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate931(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate932(.a(G10), .O(gate79inter7));
  inv1  gate933(.a(G323), .O(gate79inter8));
  nand2 gate934(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate935(.a(s_55), .b(gate79inter3), .O(gate79inter10));
  nor2  gate936(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate937(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate938(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate2437(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2438(.a(gate80inter0), .b(s_270), .O(gate80inter1));
  and2  gate2439(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2440(.a(s_270), .O(gate80inter3));
  inv1  gate2441(.a(s_271), .O(gate80inter4));
  nand2 gate2442(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2443(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2444(.a(G14), .O(gate80inter7));
  inv1  gate2445(.a(G323), .O(gate80inter8));
  nand2 gate2446(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2447(.a(s_271), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2448(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2449(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2450(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate3151(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate3152(.a(gate84inter0), .b(s_372), .O(gate84inter1));
  and2  gate3153(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate3154(.a(s_372), .O(gate84inter3));
  inv1  gate3155(.a(s_373), .O(gate84inter4));
  nand2 gate3156(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate3157(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate3158(.a(G15), .O(gate84inter7));
  inv1  gate3159(.a(G329), .O(gate84inter8));
  nand2 gate3160(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate3161(.a(s_373), .b(gate84inter3), .O(gate84inter10));
  nor2  gate3162(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate3163(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate3164(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1793(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1794(.a(gate89inter0), .b(s_178), .O(gate89inter1));
  and2  gate1795(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1796(.a(s_178), .O(gate89inter3));
  inv1  gate1797(.a(s_179), .O(gate89inter4));
  nand2 gate1798(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1799(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1800(.a(G17), .O(gate89inter7));
  inv1  gate1801(.a(G338), .O(gate89inter8));
  nand2 gate1802(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1803(.a(s_179), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1804(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1805(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1806(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate589(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate590(.a(gate91inter0), .b(s_6), .O(gate91inter1));
  and2  gate591(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate592(.a(s_6), .O(gate91inter3));
  inv1  gate593(.a(s_7), .O(gate91inter4));
  nand2 gate594(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate595(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate596(.a(G25), .O(gate91inter7));
  inv1  gate597(.a(G341), .O(gate91inter8));
  nand2 gate598(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate599(.a(s_7), .b(gate91inter3), .O(gate91inter10));
  nor2  gate600(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate601(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate602(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate3277(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate3278(.a(gate95inter0), .b(s_390), .O(gate95inter1));
  and2  gate3279(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate3280(.a(s_390), .O(gate95inter3));
  inv1  gate3281(.a(s_391), .O(gate95inter4));
  nand2 gate3282(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate3283(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate3284(.a(G26), .O(gate95inter7));
  inv1  gate3285(.a(G347), .O(gate95inter8));
  nand2 gate3286(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate3287(.a(s_391), .b(gate95inter3), .O(gate95inter10));
  nor2  gate3288(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate3289(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate3290(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2535(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2536(.a(gate97inter0), .b(s_284), .O(gate97inter1));
  and2  gate2537(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2538(.a(s_284), .O(gate97inter3));
  inv1  gate2539(.a(s_285), .O(gate97inter4));
  nand2 gate2540(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2541(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2542(.a(G19), .O(gate97inter7));
  inv1  gate2543(.a(G350), .O(gate97inter8));
  nand2 gate2544(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2545(.a(s_285), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2546(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2547(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2548(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2927(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2928(.a(gate99inter0), .b(s_340), .O(gate99inter1));
  and2  gate2929(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2930(.a(s_340), .O(gate99inter3));
  inv1  gate2931(.a(s_341), .O(gate99inter4));
  nand2 gate2932(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2933(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2934(.a(G27), .O(gate99inter7));
  inv1  gate2935(.a(G353), .O(gate99inter8));
  nand2 gate2936(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2937(.a(s_341), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2938(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2939(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2940(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate687(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate688(.a(gate101inter0), .b(s_20), .O(gate101inter1));
  and2  gate689(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate690(.a(s_20), .O(gate101inter3));
  inv1  gate691(.a(s_21), .O(gate101inter4));
  nand2 gate692(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate693(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate694(.a(G20), .O(gate101inter7));
  inv1  gate695(.a(G356), .O(gate101inter8));
  nand2 gate696(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate697(.a(s_21), .b(gate101inter3), .O(gate101inter10));
  nor2  gate698(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate699(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate700(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate2199(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2200(.a(gate103inter0), .b(s_236), .O(gate103inter1));
  and2  gate2201(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2202(.a(s_236), .O(gate103inter3));
  inv1  gate2203(.a(s_237), .O(gate103inter4));
  nand2 gate2204(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2205(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2206(.a(G28), .O(gate103inter7));
  inv1  gate2207(.a(G359), .O(gate103inter8));
  nand2 gate2208(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2209(.a(s_237), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2210(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2211(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2212(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1317(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1318(.a(gate105inter0), .b(s_110), .O(gate105inter1));
  and2  gate1319(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1320(.a(s_110), .O(gate105inter3));
  inv1  gate1321(.a(s_111), .O(gate105inter4));
  nand2 gate1322(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1323(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1324(.a(G362), .O(gate105inter7));
  inv1  gate1325(.a(G363), .O(gate105inter8));
  nand2 gate1326(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1327(.a(s_111), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1328(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1329(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1330(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate2745(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2746(.a(gate106inter0), .b(s_314), .O(gate106inter1));
  and2  gate2747(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2748(.a(s_314), .O(gate106inter3));
  inv1  gate2749(.a(s_315), .O(gate106inter4));
  nand2 gate2750(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2751(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2752(.a(G364), .O(gate106inter7));
  inv1  gate2753(.a(G365), .O(gate106inter8));
  nand2 gate2754(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2755(.a(s_315), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2756(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2757(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2758(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate3263(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate3264(.a(gate107inter0), .b(s_388), .O(gate107inter1));
  and2  gate3265(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate3266(.a(s_388), .O(gate107inter3));
  inv1  gate3267(.a(s_389), .O(gate107inter4));
  nand2 gate3268(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate3269(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate3270(.a(G366), .O(gate107inter7));
  inv1  gate3271(.a(G367), .O(gate107inter8));
  nand2 gate3272(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate3273(.a(s_389), .b(gate107inter3), .O(gate107inter10));
  nor2  gate3274(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate3275(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate3276(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1933(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1934(.a(gate109inter0), .b(s_198), .O(gate109inter1));
  and2  gate1935(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1936(.a(s_198), .O(gate109inter3));
  inv1  gate1937(.a(s_199), .O(gate109inter4));
  nand2 gate1938(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1939(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1940(.a(G370), .O(gate109inter7));
  inv1  gate1941(.a(G371), .O(gate109inter8));
  nand2 gate1942(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1943(.a(s_199), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1944(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1945(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1946(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1541(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1542(.a(gate111inter0), .b(s_142), .O(gate111inter1));
  and2  gate1543(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1544(.a(s_142), .O(gate111inter3));
  inv1  gate1545(.a(s_143), .O(gate111inter4));
  nand2 gate1546(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1547(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1548(.a(G374), .O(gate111inter7));
  inv1  gate1549(.a(G375), .O(gate111inter8));
  nand2 gate1550(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1551(.a(s_143), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1552(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1553(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1554(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1821(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1822(.a(gate112inter0), .b(s_182), .O(gate112inter1));
  and2  gate1823(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1824(.a(s_182), .O(gate112inter3));
  inv1  gate1825(.a(s_183), .O(gate112inter4));
  nand2 gate1826(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1827(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1828(.a(G376), .O(gate112inter7));
  inv1  gate1829(.a(G377), .O(gate112inter8));
  nand2 gate1830(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1831(.a(s_183), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1832(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1833(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1834(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1079(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1080(.a(gate115inter0), .b(s_76), .O(gate115inter1));
  and2  gate1081(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1082(.a(s_76), .O(gate115inter3));
  inv1  gate1083(.a(s_77), .O(gate115inter4));
  nand2 gate1084(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1085(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1086(.a(G382), .O(gate115inter7));
  inv1  gate1087(.a(G383), .O(gate115inter8));
  nand2 gate1088(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1089(.a(s_77), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1090(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1091(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1092(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1247(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1248(.a(gate117inter0), .b(s_100), .O(gate117inter1));
  and2  gate1249(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1250(.a(s_100), .O(gate117inter3));
  inv1  gate1251(.a(s_101), .O(gate117inter4));
  nand2 gate1252(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1253(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1254(.a(G386), .O(gate117inter7));
  inv1  gate1255(.a(G387), .O(gate117inter8));
  nand2 gate1256(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1257(.a(s_101), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1258(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1259(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1260(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate631(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate632(.a(gate120inter0), .b(s_12), .O(gate120inter1));
  and2  gate633(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate634(.a(s_12), .O(gate120inter3));
  inv1  gate635(.a(s_13), .O(gate120inter4));
  nand2 gate636(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate637(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate638(.a(G392), .O(gate120inter7));
  inv1  gate639(.a(G393), .O(gate120inter8));
  nand2 gate640(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate641(.a(s_13), .b(gate120inter3), .O(gate120inter10));
  nor2  gate642(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate643(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate644(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate673(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate674(.a(gate125inter0), .b(s_18), .O(gate125inter1));
  and2  gate675(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate676(.a(s_18), .O(gate125inter3));
  inv1  gate677(.a(s_19), .O(gate125inter4));
  nand2 gate678(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate679(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate680(.a(G402), .O(gate125inter7));
  inv1  gate681(.a(G403), .O(gate125inter8));
  nand2 gate682(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate683(.a(s_19), .b(gate125inter3), .O(gate125inter10));
  nor2  gate684(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate685(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate686(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1779(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1780(.a(gate126inter0), .b(s_176), .O(gate126inter1));
  and2  gate1781(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1782(.a(s_176), .O(gate126inter3));
  inv1  gate1783(.a(s_177), .O(gate126inter4));
  nand2 gate1784(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1785(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1786(.a(G404), .O(gate126inter7));
  inv1  gate1787(.a(G405), .O(gate126inter8));
  nand2 gate1788(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1789(.a(s_177), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1790(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1791(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1792(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate939(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate940(.a(gate128inter0), .b(s_56), .O(gate128inter1));
  and2  gate941(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate942(.a(s_56), .O(gate128inter3));
  inv1  gate943(.a(s_57), .O(gate128inter4));
  nand2 gate944(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate945(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate946(.a(G408), .O(gate128inter7));
  inv1  gate947(.a(G409), .O(gate128inter8));
  nand2 gate948(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate949(.a(s_57), .b(gate128inter3), .O(gate128inter10));
  nor2  gate950(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate951(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate952(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate3347(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate3348(.a(gate132inter0), .b(s_400), .O(gate132inter1));
  and2  gate3349(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate3350(.a(s_400), .O(gate132inter3));
  inv1  gate3351(.a(s_401), .O(gate132inter4));
  nand2 gate3352(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate3353(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate3354(.a(G416), .O(gate132inter7));
  inv1  gate3355(.a(G417), .O(gate132inter8));
  nand2 gate3356(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate3357(.a(s_401), .b(gate132inter3), .O(gate132inter10));
  nor2  gate3358(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate3359(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate3360(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate967(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate968(.a(gate134inter0), .b(s_60), .O(gate134inter1));
  and2  gate969(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate970(.a(s_60), .O(gate134inter3));
  inv1  gate971(.a(s_61), .O(gate134inter4));
  nand2 gate972(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate973(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate974(.a(G420), .O(gate134inter7));
  inv1  gate975(.a(G421), .O(gate134inter8));
  nand2 gate976(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate977(.a(s_61), .b(gate134inter3), .O(gate134inter10));
  nor2  gate978(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate979(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate980(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate757(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate758(.a(gate138inter0), .b(s_30), .O(gate138inter1));
  and2  gate759(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate760(.a(s_30), .O(gate138inter3));
  inv1  gate761(.a(s_31), .O(gate138inter4));
  nand2 gate762(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate763(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate764(.a(G432), .O(gate138inter7));
  inv1  gate765(.a(G435), .O(gate138inter8));
  nand2 gate766(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate767(.a(s_31), .b(gate138inter3), .O(gate138inter10));
  nor2  gate768(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate769(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate770(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1597(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1598(.a(gate140inter0), .b(s_150), .O(gate140inter1));
  and2  gate1599(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1600(.a(s_150), .O(gate140inter3));
  inv1  gate1601(.a(s_151), .O(gate140inter4));
  nand2 gate1602(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1603(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1604(.a(G444), .O(gate140inter7));
  inv1  gate1605(.a(G447), .O(gate140inter8));
  nand2 gate1606(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1607(.a(s_151), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1608(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1609(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1610(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2423(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2424(.a(gate143inter0), .b(s_268), .O(gate143inter1));
  and2  gate2425(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2426(.a(s_268), .O(gate143inter3));
  inv1  gate2427(.a(s_269), .O(gate143inter4));
  nand2 gate2428(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2429(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2430(.a(G462), .O(gate143inter7));
  inv1  gate2431(.a(G465), .O(gate143inter8));
  nand2 gate2432(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2433(.a(s_269), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2434(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2435(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2436(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate3179(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate3180(.a(gate144inter0), .b(s_376), .O(gate144inter1));
  and2  gate3181(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate3182(.a(s_376), .O(gate144inter3));
  inv1  gate3183(.a(s_377), .O(gate144inter4));
  nand2 gate3184(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate3185(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate3186(.a(G468), .O(gate144inter7));
  inv1  gate3187(.a(G471), .O(gate144inter8));
  nand2 gate3188(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate3189(.a(s_377), .b(gate144inter3), .O(gate144inter10));
  nor2  gate3190(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate3191(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate3192(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1233(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1234(.a(gate145inter0), .b(s_98), .O(gate145inter1));
  and2  gate1235(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1236(.a(s_98), .O(gate145inter3));
  inv1  gate1237(.a(s_99), .O(gate145inter4));
  nand2 gate1238(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1239(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1240(.a(G474), .O(gate145inter7));
  inv1  gate1241(.a(G477), .O(gate145inter8));
  nand2 gate1242(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1243(.a(s_99), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1244(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1245(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1246(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1289(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1290(.a(gate146inter0), .b(s_106), .O(gate146inter1));
  and2  gate1291(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1292(.a(s_106), .O(gate146inter3));
  inv1  gate1293(.a(s_107), .O(gate146inter4));
  nand2 gate1294(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1295(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1296(.a(G480), .O(gate146inter7));
  inv1  gate1297(.a(G483), .O(gate146inter8));
  nand2 gate1298(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1299(.a(s_107), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1300(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1301(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1302(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2045(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2046(.a(gate148inter0), .b(s_214), .O(gate148inter1));
  and2  gate2047(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2048(.a(s_214), .O(gate148inter3));
  inv1  gate2049(.a(s_215), .O(gate148inter4));
  nand2 gate2050(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2051(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2052(.a(G492), .O(gate148inter7));
  inv1  gate2053(.a(G495), .O(gate148inter8));
  nand2 gate2054(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2055(.a(s_215), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2056(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2057(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2058(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate2339(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2340(.a(gate149inter0), .b(s_256), .O(gate149inter1));
  and2  gate2341(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2342(.a(s_256), .O(gate149inter3));
  inv1  gate2343(.a(s_257), .O(gate149inter4));
  nand2 gate2344(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2345(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2346(.a(G498), .O(gate149inter7));
  inv1  gate2347(.a(G501), .O(gate149inter8));
  nand2 gate2348(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2349(.a(s_257), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2350(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2351(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2352(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2073(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2074(.a(gate151inter0), .b(s_218), .O(gate151inter1));
  and2  gate2075(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2076(.a(s_218), .O(gate151inter3));
  inv1  gate2077(.a(s_219), .O(gate151inter4));
  nand2 gate2078(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2079(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2080(.a(G510), .O(gate151inter7));
  inv1  gate2081(.a(G513), .O(gate151inter8));
  nand2 gate2082(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2083(.a(s_219), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2084(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2085(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2086(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2157(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2158(.a(gate153inter0), .b(s_230), .O(gate153inter1));
  and2  gate2159(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2160(.a(s_230), .O(gate153inter3));
  inv1  gate2161(.a(s_231), .O(gate153inter4));
  nand2 gate2162(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2163(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2164(.a(G426), .O(gate153inter7));
  inv1  gate2165(.a(G522), .O(gate153inter8));
  nand2 gate2166(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2167(.a(s_231), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2168(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2169(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2170(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2451(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2452(.a(gate154inter0), .b(s_272), .O(gate154inter1));
  and2  gate2453(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2454(.a(s_272), .O(gate154inter3));
  inv1  gate2455(.a(s_273), .O(gate154inter4));
  nand2 gate2456(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2457(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2458(.a(G429), .O(gate154inter7));
  inv1  gate2459(.a(G522), .O(gate154inter8));
  nand2 gate2460(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2461(.a(s_273), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2462(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2463(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2464(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2857(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2858(.a(gate155inter0), .b(s_330), .O(gate155inter1));
  and2  gate2859(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2860(.a(s_330), .O(gate155inter3));
  inv1  gate2861(.a(s_331), .O(gate155inter4));
  nand2 gate2862(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2863(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2864(.a(G432), .O(gate155inter7));
  inv1  gate2865(.a(G525), .O(gate155inter8));
  nand2 gate2866(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2867(.a(s_331), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2868(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2869(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2870(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2255(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2256(.a(gate156inter0), .b(s_244), .O(gate156inter1));
  and2  gate2257(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2258(.a(s_244), .O(gate156inter3));
  inv1  gate2259(.a(s_245), .O(gate156inter4));
  nand2 gate2260(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2261(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2262(.a(G435), .O(gate156inter7));
  inv1  gate2263(.a(G525), .O(gate156inter8));
  nand2 gate2264(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2265(.a(s_245), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2266(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2267(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2268(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2213(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2214(.a(gate160inter0), .b(s_238), .O(gate160inter1));
  and2  gate2215(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2216(.a(s_238), .O(gate160inter3));
  inv1  gate2217(.a(s_239), .O(gate160inter4));
  nand2 gate2218(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2219(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2220(.a(G447), .O(gate160inter7));
  inv1  gate2221(.a(G531), .O(gate160inter8));
  nand2 gate2222(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2223(.a(s_239), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2224(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2225(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2226(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate2843(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2844(.a(gate161inter0), .b(s_328), .O(gate161inter1));
  and2  gate2845(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2846(.a(s_328), .O(gate161inter3));
  inv1  gate2847(.a(s_329), .O(gate161inter4));
  nand2 gate2848(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2849(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2850(.a(G450), .O(gate161inter7));
  inv1  gate2851(.a(G534), .O(gate161inter8));
  nand2 gate2852(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2853(.a(s_329), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2854(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2855(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2856(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate3165(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate3166(.a(gate165inter0), .b(s_374), .O(gate165inter1));
  and2  gate3167(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate3168(.a(s_374), .O(gate165inter3));
  inv1  gate3169(.a(s_375), .O(gate165inter4));
  nand2 gate3170(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate3171(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate3172(.a(G462), .O(gate165inter7));
  inv1  gate3173(.a(G540), .O(gate165inter8));
  nand2 gate3174(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate3175(.a(s_375), .b(gate165inter3), .O(gate165inter10));
  nor2  gate3176(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate3177(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate3178(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1219(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1220(.a(gate167inter0), .b(s_96), .O(gate167inter1));
  and2  gate1221(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1222(.a(s_96), .O(gate167inter3));
  inv1  gate1223(.a(s_97), .O(gate167inter4));
  nand2 gate1224(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1225(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1226(.a(G468), .O(gate167inter7));
  inv1  gate1227(.a(G543), .O(gate167inter8));
  nand2 gate1228(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1229(.a(s_97), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1230(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1231(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1232(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate813(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate814(.a(gate169inter0), .b(s_38), .O(gate169inter1));
  and2  gate815(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate816(.a(s_38), .O(gate169inter3));
  inv1  gate817(.a(s_39), .O(gate169inter4));
  nand2 gate818(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate819(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate820(.a(G474), .O(gate169inter7));
  inv1  gate821(.a(G546), .O(gate169inter8));
  nand2 gate822(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate823(.a(s_39), .b(gate169inter3), .O(gate169inter10));
  nor2  gate824(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate825(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate826(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2367(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2368(.a(gate170inter0), .b(s_260), .O(gate170inter1));
  and2  gate2369(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2370(.a(s_260), .O(gate170inter3));
  inv1  gate2371(.a(s_261), .O(gate170inter4));
  nand2 gate2372(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2373(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2374(.a(G477), .O(gate170inter7));
  inv1  gate2375(.a(G546), .O(gate170inter8));
  nand2 gate2376(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2377(.a(s_261), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2378(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2379(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2380(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate561(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate562(.a(gate171inter0), .b(s_2), .O(gate171inter1));
  and2  gate563(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate564(.a(s_2), .O(gate171inter3));
  inv1  gate565(.a(s_3), .O(gate171inter4));
  nand2 gate566(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate567(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate568(.a(G480), .O(gate171inter7));
  inv1  gate569(.a(G549), .O(gate171inter8));
  nand2 gate570(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate571(.a(s_3), .b(gate171inter3), .O(gate171inter10));
  nor2  gate572(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate573(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate574(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate897(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate898(.a(gate173inter0), .b(s_50), .O(gate173inter1));
  and2  gate899(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate900(.a(s_50), .O(gate173inter3));
  inv1  gate901(.a(s_51), .O(gate173inter4));
  nand2 gate902(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate903(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate904(.a(G486), .O(gate173inter7));
  inv1  gate905(.a(G552), .O(gate173inter8));
  nand2 gate906(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate907(.a(s_51), .b(gate173inter3), .O(gate173inter10));
  nor2  gate908(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate909(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate910(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1499(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1500(.a(gate175inter0), .b(s_136), .O(gate175inter1));
  and2  gate1501(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1502(.a(s_136), .O(gate175inter3));
  inv1  gate1503(.a(s_137), .O(gate175inter4));
  nand2 gate1504(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1505(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1506(.a(G492), .O(gate175inter7));
  inv1  gate1507(.a(G555), .O(gate175inter8));
  nand2 gate1508(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1509(.a(s_137), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1510(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1511(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1512(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate911(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate912(.a(gate180inter0), .b(s_52), .O(gate180inter1));
  and2  gate913(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate914(.a(s_52), .O(gate180inter3));
  inv1  gate915(.a(s_53), .O(gate180inter4));
  nand2 gate916(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate917(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate918(.a(G507), .O(gate180inter7));
  inv1  gate919(.a(G561), .O(gate180inter8));
  nand2 gate920(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate921(.a(s_53), .b(gate180inter3), .O(gate180inter10));
  nor2  gate922(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate923(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate924(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2087(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2088(.a(gate182inter0), .b(s_220), .O(gate182inter1));
  and2  gate2089(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2090(.a(s_220), .O(gate182inter3));
  inv1  gate2091(.a(s_221), .O(gate182inter4));
  nand2 gate2092(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2093(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2094(.a(G513), .O(gate182inter7));
  inv1  gate2095(.a(G564), .O(gate182inter8));
  nand2 gate2096(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2097(.a(s_221), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2098(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2099(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2100(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate953(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate954(.a(gate187inter0), .b(s_58), .O(gate187inter1));
  and2  gate955(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate956(.a(s_58), .O(gate187inter3));
  inv1  gate957(.a(s_59), .O(gate187inter4));
  nand2 gate958(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate959(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate960(.a(G574), .O(gate187inter7));
  inv1  gate961(.a(G575), .O(gate187inter8));
  nand2 gate962(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate963(.a(s_59), .b(gate187inter3), .O(gate187inter10));
  nor2  gate964(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate965(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate966(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate617(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate618(.a(gate192inter0), .b(s_10), .O(gate192inter1));
  and2  gate619(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate620(.a(s_10), .O(gate192inter3));
  inv1  gate621(.a(s_11), .O(gate192inter4));
  nand2 gate622(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate623(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate624(.a(G584), .O(gate192inter7));
  inv1  gate625(.a(G585), .O(gate192inter8));
  nand2 gate626(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate627(.a(s_11), .b(gate192inter3), .O(gate192inter10));
  nor2  gate628(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate629(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate630(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate659(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate660(.a(gate193inter0), .b(s_16), .O(gate193inter1));
  and2  gate661(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate662(.a(s_16), .O(gate193inter3));
  inv1  gate663(.a(s_17), .O(gate193inter4));
  nand2 gate664(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate665(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate666(.a(G586), .O(gate193inter7));
  inv1  gate667(.a(G587), .O(gate193inter8));
  nand2 gate668(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate669(.a(s_17), .b(gate193inter3), .O(gate193inter10));
  nor2  gate670(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate671(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate672(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate3333(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate3334(.a(gate196inter0), .b(s_398), .O(gate196inter1));
  and2  gate3335(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate3336(.a(s_398), .O(gate196inter3));
  inv1  gate3337(.a(s_399), .O(gate196inter4));
  nand2 gate3338(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate3339(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate3340(.a(G592), .O(gate196inter7));
  inv1  gate3341(.a(G593), .O(gate196inter8));
  nand2 gate3342(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate3343(.a(s_399), .b(gate196inter3), .O(gate196inter10));
  nor2  gate3344(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate3345(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate3346(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate771(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate772(.a(gate198inter0), .b(s_32), .O(gate198inter1));
  and2  gate773(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate774(.a(s_32), .O(gate198inter3));
  inv1  gate775(.a(s_33), .O(gate198inter4));
  nand2 gate776(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate777(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate778(.a(G596), .O(gate198inter7));
  inv1  gate779(.a(G597), .O(gate198inter8));
  nand2 gate780(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate781(.a(s_33), .b(gate198inter3), .O(gate198inter10));
  nor2  gate782(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate783(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate784(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2325(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2326(.a(gate199inter0), .b(s_254), .O(gate199inter1));
  and2  gate2327(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2328(.a(s_254), .O(gate199inter3));
  inv1  gate2329(.a(s_255), .O(gate199inter4));
  nand2 gate2330(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2331(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2332(.a(G598), .O(gate199inter7));
  inv1  gate2333(.a(G599), .O(gate199inter8));
  nand2 gate2334(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2335(.a(s_255), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2336(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2337(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2338(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1961(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1962(.a(gate200inter0), .b(s_202), .O(gate200inter1));
  and2  gate1963(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1964(.a(s_202), .O(gate200inter3));
  inv1  gate1965(.a(s_203), .O(gate200inter4));
  nand2 gate1966(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1967(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1968(.a(G600), .O(gate200inter7));
  inv1  gate1969(.a(G601), .O(gate200inter8));
  nand2 gate1970(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1971(.a(s_203), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1972(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1973(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1974(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1471(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1472(.a(gate201inter0), .b(s_132), .O(gate201inter1));
  and2  gate1473(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1474(.a(s_132), .O(gate201inter3));
  inv1  gate1475(.a(s_133), .O(gate201inter4));
  nand2 gate1476(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1477(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1478(.a(G602), .O(gate201inter7));
  inv1  gate1479(.a(G607), .O(gate201inter8));
  nand2 gate1480(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1481(.a(s_133), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1482(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1483(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1484(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1555(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1556(.a(gate203inter0), .b(s_144), .O(gate203inter1));
  and2  gate1557(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1558(.a(s_144), .O(gate203inter3));
  inv1  gate1559(.a(s_145), .O(gate203inter4));
  nand2 gate1560(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1561(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1562(.a(G602), .O(gate203inter7));
  inv1  gate1563(.a(G612), .O(gate203inter8));
  nand2 gate1564(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1565(.a(s_145), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1566(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1567(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1568(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate2465(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2466(.a(gate204inter0), .b(s_274), .O(gate204inter1));
  and2  gate2467(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2468(.a(s_274), .O(gate204inter3));
  inv1  gate2469(.a(s_275), .O(gate204inter4));
  nand2 gate2470(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2471(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2472(.a(G607), .O(gate204inter7));
  inv1  gate2473(.a(G617), .O(gate204inter8));
  nand2 gate2474(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2475(.a(s_275), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2476(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2477(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2478(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate981(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate982(.a(gate206inter0), .b(s_62), .O(gate206inter1));
  and2  gate983(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate984(.a(s_62), .O(gate206inter3));
  inv1  gate985(.a(s_63), .O(gate206inter4));
  nand2 gate986(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate987(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate988(.a(G632), .O(gate206inter7));
  inv1  gate989(.a(G637), .O(gate206inter8));
  nand2 gate990(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate991(.a(s_63), .b(gate206inter3), .O(gate206inter10));
  nor2  gate992(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate993(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate994(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1303(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1304(.a(gate208inter0), .b(s_108), .O(gate208inter1));
  and2  gate1305(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1306(.a(s_108), .O(gate208inter3));
  inv1  gate1307(.a(s_109), .O(gate208inter4));
  nand2 gate1308(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1309(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1310(.a(G627), .O(gate208inter7));
  inv1  gate1311(.a(G637), .O(gate208inter8));
  nand2 gate1312(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1313(.a(s_109), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1314(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1315(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1316(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate3137(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate3138(.a(gate209inter0), .b(s_370), .O(gate209inter1));
  and2  gate3139(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate3140(.a(s_370), .O(gate209inter3));
  inv1  gate3141(.a(s_371), .O(gate209inter4));
  nand2 gate3142(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate3143(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate3144(.a(G602), .O(gate209inter7));
  inv1  gate3145(.a(G666), .O(gate209inter8));
  nand2 gate3146(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate3147(.a(s_371), .b(gate209inter3), .O(gate209inter10));
  nor2  gate3148(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate3149(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate3150(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate3319(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate3320(.a(gate210inter0), .b(s_396), .O(gate210inter1));
  and2  gate3321(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate3322(.a(s_396), .O(gate210inter3));
  inv1  gate3323(.a(s_397), .O(gate210inter4));
  nand2 gate3324(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate3325(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate3326(.a(G607), .O(gate210inter7));
  inv1  gate3327(.a(G666), .O(gate210inter8));
  nand2 gate3328(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate3329(.a(s_397), .b(gate210inter3), .O(gate210inter10));
  nor2  gate3330(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate3331(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate3332(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate2129(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2130(.a(gate211inter0), .b(s_226), .O(gate211inter1));
  and2  gate2131(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2132(.a(s_226), .O(gate211inter3));
  inv1  gate2133(.a(s_227), .O(gate211inter4));
  nand2 gate2134(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2135(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2136(.a(G612), .O(gate211inter7));
  inv1  gate2137(.a(G669), .O(gate211inter8));
  nand2 gate2138(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2139(.a(s_227), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2140(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2141(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2142(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate3081(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate3082(.a(gate213inter0), .b(s_362), .O(gate213inter1));
  and2  gate3083(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate3084(.a(s_362), .O(gate213inter3));
  inv1  gate3085(.a(s_363), .O(gate213inter4));
  nand2 gate3086(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate3087(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate3088(.a(G602), .O(gate213inter7));
  inv1  gate3089(.a(G672), .O(gate213inter8));
  nand2 gate3090(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate3091(.a(s_363), .b(gate213inter3), .O(gate213inter10));
  nor2  gate3092(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate3093(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate3094(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1625(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1626(.a(gate215inter0), .b(s_154), .O(gate215inter1));
  and2  gate1627(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1628(.a(s_154), .O(gate215inter3));
  inv1  gate1629(.a(s_155), .O(gate215inter4));
  nand2 gate1630(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1631(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1632(.a(G607), .O(gate215inter7));
  inv1  gate1633(.a(G675), .O(gate215inter8));
  nand2 gate1634(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1635(.a(s_155), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1636(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1637(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1638(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate701(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate702(.a(gate216inter0), .b(s_22), .O(gate216inter1));
  and2  gate703(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate704(.a(s_22), .O(gate216inter3));
  inv1  gate705(.a(s_23), .O(gate216inter4));
  nand2 gate706(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate707(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate708(.a(G617), .O(gate216inter7));
  inv1  gate709(.a(G675), .O(gate216inter8));
  nand2 gate710(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate711(.a(s_23), .b(gate216inter3), .O(gate216inter10));
  nor2  gate712(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate713(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate714(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2227(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2228(.a(gate219inter0), .b(s_240), .O(gate219inter1));
  and2  gate2229(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2230(.a(s_240), .O(gate219inter3));
  inv1  gate2231(.a(s_241), .O(gate219inter4));
  nand2 gate2232(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2233(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2234(.a(G632), .O(gate219inter7));
  inv1  gate2235(.a(G681), .O(gate219inter8));
  nand2 gate2236(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2237(.a(s_241), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2238(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2239(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2240(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1891(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1892(.a(gate220inter0), .b(s_192), .O(gate220inter1));
  and2  gate1893(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1894(.a(s_192), .O(gate220inter3));
  inv1  gate1895(.a(s_193), .O(gate220inter4));
  nand2 gate1896(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1897(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1898(.a(G637), .O(gate220inter7));
  inv1  gate1899(.a(G681), .O(gate220inter8));
  nand2 gate1900(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1901(.a(s_193), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1902(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1903(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1904(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate3207(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate3208(.a(gate221inter0), .b(s_380), .O(gate221inter1));
  and2  gate3209(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate3210(.a(s_380), .O(gate221inter3));
  inv1  gate3211(.a(s_381), .O(gate221inter4));
  nand2 gate3212(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate3213(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate3214(.a(G622), .O(gate221inter7));
  inv1  gate3215(.a(G684), .O(gate221inter8));
  nand2 gate3216(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate3217(.a(s_381), .b(gate221inter3), .O(gate221inter10));
  nor2  gate3218(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate3219(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate3220(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate2521(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2522(.a(gate222inter0), .b(s_282), .O(gate222inter1));
  and2  gate2523(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2524(.a(s_282), .O(gate222inter3));
  inv1  gate2525(.a(s_283), .O(gate222inter4));
  nand2 gate2526(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2527(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2528(.a(G632), .O(gate222inter7));
  inv1  gate2529(.a(G684), .O(gate222inter8));
  nand2 gate2530(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2531(.a(s_283), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2532(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2533(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2534(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1667(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1668(.a(gate223inter0), .b(s_160), .O(gate223inter1));
  and2  gate1669(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1670(.a(s_160), .O(gate223inter3));
  inv1  gate1671(.a(s_161), .O(gate223inter4));
  nand2 gate1672(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1673(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1674(.a(G627), .O(gate223inter7));
  inv1  gate1675(.a(G687), .O(gate223inter8));
  nand2 gate1676(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1677(.a(s_161), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1678(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1679(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1680(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate2115(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2116(.a(gate224inter0), .b(s_224), .O(gate224inter1));
  and2  gate2117(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2118(.a(s_224), .O(gate224inter3));
  inv1  gate2119(.a(s_225), .O(gate224inter4));
  nand2 gate2120(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2121(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2122(.a(G637), .O(gate224inter7));
  inv1  gate2123(.a(G687), .O(gate224inter8));
  nand2 gate2124(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2125(.a(s_225), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2126(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2127(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2128(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate3011(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate3012(.a(gate225inter0), .b(s_352), .O(gate225inter1));
  and2  gate3013(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate3014(.a(s_352), .O(gate225inter3));
  inv1  gate3015(.a(s_353), .O(gate225inter4));
  nand2 gate3016(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate3017(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate3018(.a(G690), .O(gate225inter7));
  inv1  gate3019(.a(G691), .O(gate225inter8));
  nand2 gate3020(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate3021(.a(s_353), .b(gate225inter3), .O(gate225inter10));
  nor2  gate3022(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate3023(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate3024(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1765(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1766(.a(gate226inter0), .b(s_174), .O(gate226inter1));
  and2  gate1767(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1768(.a(s_174), .O(gate226inter3));
  inv1  gate1769(.a(s_175), .O(gate226inter4));
  nand2 gate1770(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1771(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1772(.a(G692), .O(gate226inter7));
  inv1  gate1773(.a(G693), .O(gate226inter8));
  nand2 gate1774(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1775(.a(s_175), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1776(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1777(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1778(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1415(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1416(.a(gate227inter0), .b(s_124), .O(gate227inter1));
  and2  gate1417(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1418(.a(s_124), .O(gate227inter3));
  inv1  gate1419(.a(s_125), .O(gate227inter4));
  nand2 gate1420(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1421(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1422(.a(G694), .O(gate227inter7));
  inv1  gate1423(.a(G695), .O(gate227inter8));
  nand2 gate1424(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1425(.a(s_125), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1426(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1427(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1428(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate3067(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate3068(.a(gate228inter0), .b(s_360), .O(gate228inter1));
  and2  gate3069(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate3070(.a(s_360), .O(gate228inter3));
  inv1  gate3071(.a(s_361), .O(gate228inter4));
  nand2 gate3072(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate3073(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate3074(.a(G696), .O(gate228inter7));
  inv1  gate3075(.a(G697), .O(gate228inter8));
  nand2 gate3076(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate3077(.a(s_361), .b(gate228inter3), .O(gate228inter10));
  nor2  gate3078(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate3079(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate3080(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2381(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2382(.a(gate230inter0), .b(s_262), .O(gate230inter1));
  and2  gate2383(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2384(.a(s_262), .O(gate230inter3));
  inv1  gate2385(.a(s_263), .O(gate230inter4));
  nand2 gate2386(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2387(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2388(.a(G700), .O(gate230inter7));
  inv1  gate2389(.a(G701), .O(gate230inter8));
  nand2 gate2390(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2391(.a(s_263), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2392(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2393(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2394(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2493(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2494(.a(gate231inter0), .b(s_278), .O(gate231inter1));
  and2  gate2495(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2496(.a(s_278), .O(gate231inter3));
  inv1  gate2497(.a(s_279), .O(gate231inter4));
  nand2 gate2498(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2499(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2500(.a(G702), .O(gate231inter7));
  inv1  gate2501(.a(G703), .O(gate231inter8));
  nand2 gate2502(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2503(.a(s_279), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2504(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2505(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2506(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1723(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1724(.a(gate237inter0), .b(s_168), .O(gate237inter1));
  and2  gate1725(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1726(.a(s_168), .O(gate237inter3));
  inv1  gate1727(.a(s_169), .O(gate237inter4));
  nand2 gate1728(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1729(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1730(.a(G254), .O(gate237inter7));
  inv1  gate1731(.a(G706), .O(gate237inter8));
  nand2 gate1732(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1733(.a(s_169), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1734(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1735(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1736(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2283(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2284(.a(gate241inter0), .b(s_248), .O(gate241inter1));
  and2  gate2285(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2286(.a(s_248), .O(gate241inter3));
  inv1  gate2287(.a(s_249), .O(gate241inter4));
  nand2 gate2288(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2289(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2290(.a(G242), .O(gate241inter7));
  inv1  gate2291(.a(G730), .O(gate241inter8));
  nand2 gate2292(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2293(.a(s_249), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2294(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2295(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2296(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate2143(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2144(.a(gate242inter0), .b(s_228), .O(gate242inter1));
  and2  gate2145(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2146(.a(s_228), .O(gate242inter3));
  inv1  gate2147(.a(s_229), .O(gate242inter4));
  nand2 gate2148(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2149(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2150(.a(G718), .O(gate242inter7));
  inv1  gate2151(.a(G730), .O(gate242inter8));
  nand2 gate2152(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2153(.a(s_229), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2154(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2155(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2156(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1037(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1038(.a(gate244inter0), .b(s_70), .O(gate244inter1));
  and2  gate1039(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1040(.a(s_70), .O(gate244inter3));
  inv1  gate1041(.a(s_71), .O(gate244inter4));
  nand2 gate1042(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1043(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1044(.a(G721), .O(gate244inter7));
  inv1  gate1045(.a(G733), .O(gate244inter8));
  nand2 gate1046(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1047(.a(s_71), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1048(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1049(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1050(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1569(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1570(.a(gate245inter0), .b(s_146), .O(gate245inter1));
  and2  gate1571(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1572(.a(s_146), .O(gate245inter3));
  inv1  gate1573(.a(s_147), .O(gate245inter4));
  nand2 gate1574(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1575(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1576(.a(G248), .O(gate245inter7));
  inv1  gate1577(.a(G736), .O(gate245inter8));
  nand2 gate1578(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1579(.a(s_147), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1580(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1581(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1582(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2577(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2578(.a(gate248inter0), .b(s_290), .O(gate248inter1));
  and2  gate2579(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2580(.a(s_290), .O(gate248inter3));
  inv1  gate2581(.a(s_291), .O(gate248inter4));
  nand2 gate2582(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2583(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2584(.a(G727), .O(gate248inter7));
  inv1  gate2585(.a(G739), .O(gate248inter8));
  nand2 gate2586(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2587(.a(s_291), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2588(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2589(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2590(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1639(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1640(.a(gate252inter0), .b(s_156), .O(gate252inter1));
  and2  gate1641(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1642(.a(s_156), .O(gate252inter3));
  inv1  gate1643(.a(s_157), .O(gate252inter4));
  nand2 gate1644(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1645(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1646(.a(G709), .O(gate252inter7));
  inv1  gate1647(.a(G745), .O(gate252inter8));
  nand2 gate1648(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1649(.a(s_157), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1650(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1651(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1652(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2353(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2354(.a(gate254inter0), .b(s_258), .O(gate254inter1));
  and2  gate2355(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2356(.a(s_258), .O(gate254inter3));
  inv1  gate2357(.a(s_259), .O(gate254inter4));
  nand2 gate2358(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2359(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2360(.a(G712), .O(gate254inter7));
  inv1  gate2361(.a(G748), .O(gate254inter8));
  nand2 gate2362(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2363(.a(s_259), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2364(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2365(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2366(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate3095(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate3096(.a(gate255inter0), .b(s_364), .O(gate255inter1));
  and2  gate3097(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate3098(.a(s_364), .O(gate255inter3));
  inv1  gate3099(.a(s_365), .O(gate255inter4));
  nand2 gate3100(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate3101(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate3102(.a(G263), .O(gate255inter7));
  inv1  gate3103(.a(G751), .O(gate255inter8));
  nand2 gate3104(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate3105(.a(s_365), .b(gate255inter3), .O(gate255inter10));
  nor2  gate3106(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate3107(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate3108(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2885(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2886(.a(gate258inter0), .b(s_334), .O(gate258inter1));
  and2  gate2887(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2888(.a(s_334), .O(gate258inter3));
  inv1  gate2889(.a(s_335), .O(gate258inter4));
  nand2 gate2890(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2891(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2892(.a(G756), .O(gate258inter7));
  inv1  gate2893(.a(G757), .O(gate258inter8));
  nand2 gate2894(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2895(.a(s_335), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2896(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2897(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2898(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1485(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1486(.a(gate259inter0), .b(s_134), .O(gate259inter1));
  and2  gate1487(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1488(.a(s_134), .O(gate259inter3));
  inv1  gate1489(.a(s_135), .O(gate259inter4));
  nand2 gate1490(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1491(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1492(.a(G758), .O(gate259inter7));
  inv1  gate1493(.a(G759), .O(gate259inter8));
  nand2 gate1494(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1495(.a(s_135), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1496(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1497(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1498(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1205(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1206(.a(gate261inter0), .b(s_94), .O(gate261inter1));
  and2  gate1207(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1208(.a(s_94), .O(gate261inter3));
  inv1  gate1209(.a(s_95), .O(gate261inter4));
  nand2 gate1210(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1211(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1212(.a(G762), .O(gate261inter7));
  inv1  gate1213(.a(G763), .O(gate261inter8));
  nand2 gate1214(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1215(.a(s_95), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1216(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1217(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1218(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1975(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1976(.a(gate263inter0), .b(s_204), .O(gate263inter1));
  and2  gate1977(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1978(.a(s_204), .O(gate263inter3));
  inv1  gate1979(.a(s_205), .O(gate263inter4));
  nand2 gate1980(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1981(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1982(.a(G766), .O(gate263inter7));
  inv1  gate1983(.a(G767), .O(gate263inter8));
  nand2 gate1984(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1985(.a(s_205), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1986(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1987(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1988(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1527(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1528(.a(gate266inter0), .b(s_140), .O(gate266inter1));
  and2  gate1529(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1530(.a(s_140), .O(gate266inter3));
  inv1  gate1531(.a(s_141), .O(gate266inter4));
  nand2 gate1532(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1533(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1534(.a(G645), .O(gate266inter7));
  inv1  gate1535(.a(G773), .O(gate266inter8));
  nand2 gate1536(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1537(.a(s_141), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1538(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1539(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1540(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2801(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2802(.a(gate268inter0), .b(s_322), .O(gate268inter1));
  and2  gate2803(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2804(.a(s_322), .O(gate268inter3));
  inv1  gate2805(.a(s_323), .O(gate268inter4));
  nand2 gate2806(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2807(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2808(.a(G651), .O(gate268inter7));
  inv1  gate2809(.a(G779), .O(gate268inter8));
  nand2 gate2810(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2811(.a(s_323), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2812(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2813(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2814(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate603(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate604(.a(gate270inter0), .b(s_8), .O(gate270inter1));
  and2  gate605(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate606(.a(s_8), .O(gate270inter3));
  inv1  gate607(.a(s_9), .O(gate270inter4));
  nand2 gate608(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate609(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate610(.a(G657), .O(gate270inter7));
  inv1  gate611(.a(G785), .O(gate270inter8));
  nand2 gate612(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate613(.a(s_9), .b(gate270inter3), .O(gate270inter10));
  nor2  gate614(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate615(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate616(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2913(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2914(.a(gate271inter0), .b(s_338), .O(gate271inter1));
  and2  gate2915(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2916(.a(s_338), .O(gate271inter3));
  inv1  gate2917(.a(s_339), .O(gate271inter4));
  nand2 gate2918(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2919(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2920(.a(G660), .O(gate271inter7));
  inv1  gate2921(.a(G788), .O(gate271inter8));
  nand2 gate2922(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2923(.a(s_339), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2924(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2925(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2926(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2185(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2186(.a(gate272inter0), .b(s_234), .O(gate272inter1));
  and2  gate2187(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2188(.a(s_234), .O(gate272inter3));
  inv1  gate2189(.a(s_235), .O(gate272inter4));
  nand2 gate2190(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2191(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2192(.a(G663), .O(gate272inter7));
  inv1  gate2193(.a(G791), .O(gate272inter8));
  nand2 gate2194(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2195(.a(s_235), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2196(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2197(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2198(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate2003(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2004(.a(gate273inter0), .b(s_208), .O(gate273inter1));
  and2  gate2005(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2006(.a(s_208), .O(gate273inter3));
  inv1  gate2007(.a(s_209), .O(gate273inter4));
  nand2 gate2008(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2009(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2010(.a(G642), .O(gate273inter7));
  inv1  gate2011(.a(G794), .O(gate273inter8));
  nand2 gate2012(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2013(.a(s_209), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2014(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2015(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2016(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2605(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2606(.a(gate276inter0), .b(s_294), .O(gate276inter1));
  and2  gate2607(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2608(.a(s_294), .O(gate276inter3));
  inv1  gate2609(.a(s_295), .O(gate276inter4));
  nand2 gate2610(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2611(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2612(.a(G773), .O(gate276inter7));
  inv1  gate2613(.a(G797), .O(gate276inter8));
  nand2 gate2614(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2615(.a(s_295), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2616(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2617(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2618(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate715(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate716(.a(gate279inter0), .b(s_24), .O(gate279inter1));
  and2  gate717(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate718(.a(s_24), .O(gate279inter3));
  inv1  gate719(.a(s_25), .O(gate279inter4));
  nand2 gate720(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate721(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate722(.a(G651), .O(gate279inter7));
  inv1  gate723(.a(G803), .O(gate279inter8));
  nand2 gate724(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate725(.a(s_25), .b(gate279inter3), .O(gate279inter10));
  nor2  gate726(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate727(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate728(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate3039(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate3040(.a(gate281inter0), .b(s_356), .O(gate281inter1));
  and2  gate3041(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate3042(.a(s_356), .O(gate281inter3));
  inv1  gate3043(.a(s_357), .O(gate281inter4));
  nand2 gate3044(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate3045(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate3046(.a(G654), .O(gate281inter7));
  inv1  gate3047(.a(G806), .O(gate281inter8));
  nand2 gate3048(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate3049(.a(s_357), .b(gate281inter3), .O(gate281inter10));
  nor2  gate3050(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate3051(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate3052(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate799(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate800(.a(gate283inter0), .b(s_36), .O(gate283inter1));
  and2  gate801(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate802(.a(s_36), .O(gate283inter3));
  inv1  gate803(.a(s_37), .O(gate283inter4));
  nand2 gate804(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate805(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate806(.a(G657), .O(gate283inter7));
  inv1  gate807(.a(G809), .O(gate283inter8));
  nand2 gate808(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate809(.a(s_37), .b(gate283inter3), .O(gate283inter10));
  nor2  gate810(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate811(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate812(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2689(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2690(.a(gate285inter0), .b(s_306), .O(gate285inter1));
  and2  gate2691(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2692(.a(s_306), .O(gate285inter3));
  inv1  gate2693(.a(s_307), .O(gate285inter4));
  nand2 gate2694(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2695(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2696(.a(G660), .O(gate285inter7));
  inv1  gate2697(.a(G812), .O(gate285inter8));
  nand2 gate2698(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2699(.a(s_307), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2700(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2701(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2702(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1751(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1752(.a(gate286inter0), .b(s_172), .O(gate286inter1));
  and2  gate1753(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1754(.a(s_172), .O(gate286inter3));
  inv1  gate1755(.a(s_173), .O(gate286inter4));
  nand2 gate1756(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1757(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1758(.a(G788), .O(gate286inter7));
  inv1  gate1759(.a(G812), .O(gate286inter8));
  nand2 gate1760(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1761(.a(s_173), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1762(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1763(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1764(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1331(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1332(.a(gate289inter0), .b(s_112), .O(gate289inter1));
  and2  gate1333(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1334(.a(s_112), .O(gate289inter3));
  inv1  gate1335(.a(s_113), .O(gate289inter4));
  nand2 gate1336(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1337(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1338(.a(G818), .O(gate289inter7));
  inv1  gate1339(.a(G819), .O(gate289inter8));
  nand2 gate1340(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1341(.a(s_113), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1342(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1343(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1344(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1709(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1710(.a(gate291inter0), .b(s_166), .O(gate291inter1));
  and2  gate1711(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1712(.a(s_166), .O(gate291inter3));
  inv1  gate1713(.a(s_167), .O(gate291inter4));
  nand2 gate1714(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1715(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1716(.a(G822), .O(gate291inter7));
  inv1  gate1717(.a(G823), .O(gate291inter8));
  nand2 gate1718(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1719(.a(s_167), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1720(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1721(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1722(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2507(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2508(.a(gate293inter0), .b(s_280), .O(gate293inter1));
  and2  gate2509(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2510(.a(s_280), .O(gate293inter3));
  inv1  gate2511(.a(s_281), .O(gate293inter4));
  nand2 gate2512(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2513(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2514(.a(G828), .O(gate293inter7));
  inv1  gate2515(.a(G829), .O(gate293inter8));
  nand2 gate2516(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2517(.a(s_281), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2518(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2519(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2520(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2479(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2480(.a(gate295inter0), .b(s_276), .O(gate295inter1));
  and2  gate2481(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2482(.a(s_276), .O(gate295inter3));
  inv1  gate2483(.a(s_277), .O(gate295inter4));
  nand2 gate2484(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2485(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2486(.a(G830), .O(gate295inter7));
  inv1  gate2487(.a(G831), .O(gate295inter8));
  nand2 gate2488(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2489(.a(s_277), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2490(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2491(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2492(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate3123(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate3124(.a(gate296inter0), .b(s_368), .O(gate296inter1));
  and2  gate3125(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate3126(.a(s_368), .O(gate296inter3));
  inv1  gate3127(.a(s_369), .O(gate296inter4));
  nand2 gate3128(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate3129(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate3130(.a(G826), .O(gate296inter7));
  inv1  gate3131(.a(G827), .O(gate296inter8));
  nand2 gate3132(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate3133(.a(s_369), .b(gate296inter3), .O(gate296inter10));
  nor2  gate3134(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate3135(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate3136(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1807(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1808(.a(gate387inter0), .b(s_180), .O(gate387inter1));
  and2  gate1809(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1810(.a(s_180), .O(gate387inter3));
  inv1  gate1811(.a(s_181), .O(gate387inter4));
  nand2 gate1812(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1813(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1814(.a(G1), .O(gate387inter7));
  inv1  gate1815(.a(G1036), .O(gate387inter8));
  nand2 gate1816(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1817(.a(s_181), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1818(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1819(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1820(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2633(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2634(.a(gate391inter0), .b(s_298), .O(gate391inter1));
  and2  gate2635(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2636(.a(s_298), .O(gate391inter3));
  inv1  gate2637(.a(s_299), .O(gate391inter4));
  nand2 gate2638(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2639(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2640(.a(G5), .O(gate391inter7));
  inv1  gate2641(.a(G1048), .O(gate391inter8));
  nand2 gate2642(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2643(.a(s_299), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2644(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2645(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2646(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate2759(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2760(.a(gate392inter0), .b(s_316), .O(gate392inter1));
  and2  gate2761(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2762(.a(s_316), .O(gate392inter3));
  inv1  gate2763(.a(s_317), .O(gate392inter4));
  nand2 gate2764(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2765(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2766(.a(G6), .O(gate392inter7));
  inv1  gate2767(.a(G1051), .O(gate392inter8));
  nand2 gate2768(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2769(.a(s_317), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2770(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2771(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2772(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1457(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1458(.a(gate396inter0), .b(s_130), .O(gate396inter1));
  and2  gate1459(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1460(.a(s_130), .O(gate396inter3));
  inv1  gate1461(.a(s_131), .O(gate396inter4));
  nand2 gate1462(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1463(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1464(.a(G10), .O(gate396inter7));
  inv1  gate1465(.a(G1063), .O(gate396inter8));
  nand2 gate1466(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1467(.a(s_131), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1468(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1469(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1470(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate883(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate884(.a(gate397inter0), .b(s_48), .O(gate397inter1));
  and2  gate885(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate886(.a(s_48), .O(gate397inter3));
  inv1  gate887(.a(s_49), .O(gate397inter4));
  nand2 gate888(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate889(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate890(.a(G11), .O(gate397inter7));
  inv1  gate891(.a(G1066), .O(gate397inter8));
  nand2 gate892(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate893(.a(s_49), .b(gate397inter3), .O(gate397inter10));
  nor2  gate894(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate895(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate896(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2787(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2788(.a(gate398inter0), .b(s_320), .O(gate398inter1));
  and2  gate2789(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2790(.a(s_320), .O(gate398inter3));
  inv1  gate2791(.a(s_321), .O(gate398inter4));
  nand2 gate2792(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2793(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2794(.a(G12), .O(gate398inter7));
  inv1  gate2795(.a(G1069), .O(gate398inter8));
  nand2 gate2796(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2797(.a(s_321), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2798(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2799(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2800(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1261(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1262(.a(gate400inter0), .b(s_102), .O(gate400inter1));
  and2  gate1263(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1264(.a(s_102), .O(gate400inter3));
  inv1  gate1265(.a(s_103), .O(gate400inter4));
  nand2 gate1266(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1267(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1268(.a(G14), .O(gate400inter7));
  inv1  gate1269(.a(G1075), .O(gate400inter8));
  nand2 gate1270(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1271(.a(s_103), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1272(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1273(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1274(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2591(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2592(.a(gate406inter0), .b(s_292), .O(gate406inter1));
  and2  gate2593(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2594(.a(s_292), .O(gate406inter3));
  inv1  gate2595(.a(s_293), .O(gate406inter4));
  nand2 gate2596(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2597(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2598(.a(G20), .O(gate406inter7));
  inv1  gate2599(.a(G1093), .O(gate406inter8));
  nand2 gate2600(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2601(.a(s_293), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2602(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2603(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2604(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1345(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1346(.a(gate413inter0), .b(s_114), .O(gate413inter1));
  and2  gate1347(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1348(.a(s_114), .O(gate413inter3));
  inv1  gate1349(.a(s_115), .O(gate413inter4));
  nand2 gate1350(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1351(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1352(.a(G27), .O(gate413inter7));
  inv1  gate1353(.a(G1114), .O(gate413inter8));
  nand2 gate1354(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1355(.a(s_115), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1356(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1357(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1358(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate869(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate870(.a(gate414inter0), .b(s_46), .O(gate414inter1));
  and2  gate871(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate872(.a(s_46), .O(gate414inter3));
  inv1  gate873(.a(s_47), .O(gate414inter4));
  nand2 gate874(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate875(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate876(.a(G28), .O(gate414inter7));
  inv1  gate877(.a(G1117), .O(gate414inter8));
  nand2 gate878(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate879(.a(s_47), .b(gate414inter3), .O(gate414inter10));
  nor2  gate880(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate881(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate882(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate3221(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate3222(.a(gate415inter0), .b(s_382), .O(gate415inter1));
  and2  gate3223(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate3224(.a(s_382), .O(gate415inter3));
  inv1  gate3225(.a(s_383), .O(gate415inter4));
  nand2 gate3226(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate3227(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate3228(.a(G29), .O(gate415inter7));
  inv1  gate3229(.a(G1120), .O(gate415inter8));
  nand2 gate3230(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate3231(.a(s_383), .b(gate415inter3), .O(gate415inter10));
  nor2  gate3232(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate3233(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate3234(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate3291(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate3292(.a(gate417inter0), .b(s_392), .O(gate417inter1));
  and2  gate3293(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate3294(.a(s_392), .O(gate417inter3));
  inv1  gate3295(.a(s_393), .O(gate417inter4));
  nand2 gate3296(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate3297(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate3298(.a(G31), .O(gate417inter7));
  inv1  gate3299(.a(G1126), .O(gate417inter8));
  nand2 gate3300(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate3301(.a(s_393), .b(gate417inter3), .O(gate417inter10));
  nor2  gate3302(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate3303(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate3304(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1275(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1276(.a(gate418inter0), .b(s_104), .O(gate418inter1));
  and2  gate1277(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1278(.a(s_104), .O(gate418inter3));
  inv1  gate1279(.a(s_105), .O(gate418inter4));
  nand2 gate1280(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1281(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1282(.a(G32), .O(gate418inter7));
  inv1  gate1283(.a(G1129), .O(gate418inter8));
  nand2 gate1284(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1285(.a(s_105), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1286(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1287(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1288(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1107(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1108(.a(gate419inter0), .b(s_80), .O(gate419inter1));
  and2  gate1109(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1110(.a(s_80), .O(gate419inter3));
  inv1  gate1111(.a(s_81), .O(gate419inter4));
  nand2 gate1112(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1113(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1114(.a(G1), .O(gate419inter7));
  inv1  gate1115(.a(G1132), .O(gate419inter8));
  nand2 gate1116(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1117(.a(s_81), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1118(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1119(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1120(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1163(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1164(.a(gate420inter0), .b(s_88), .O(gate420inter1));
  and2  gate1165(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1166(.a(s_88), .O(gate420inter3));
  inv1  gate1167(.a(s_89), .O(gate420inter4));
  nand2 gate1168(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1169(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1170(.a(G1036), .O(gate420inter7));
  inv1  gate1171(.a(G1132), .O(gate420inter8));
  nand2 gate1172(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1173(.a(s_89), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1174(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1175(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1176(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2969(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2970(.a(gate422inter0), .b(s_346), .O(gate422inter1));
  and2  gate2971(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2972(.a(s_346), .O(gate422inter3));
  inv1  gate2973(.a(s_347), .O(gate422inter4));
  nand2 gate2974(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2975(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2976(.a(G1039), .O(gate422inter7));
  inv1  gate2977(.a(G1135), .O(gate422inter8));
  nand2 gate2978(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2979(.a(s_347), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2980(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2981(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2982(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1835(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1836(.a(gate429inter0), .b(s_184), .O(gate429inter1));
  and2  gate1837(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1838(.a(s_184), .O(gate429inter3));
  inv1  gate1839(.a(s_185), .O(gate429inter4));
  nand2 gate1840(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1841(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1842(.a(G6), .O(gate429inter7));
  inv1  gate1843(.a(G1147), .O(gate429inter8));
  nand2 gate1844(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1845(.a(s_185), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1846(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1847(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1848(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate2717(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2718(.a(gate430inter0), .b(s_310), .O(gate430inter1));
  and2  gate2719(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2720(.a(s_310), .O(gate430inter3));
  inv1  gate2721(.a(s_311), .O(gate430inter4));
  nand2 gate2722(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2723(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2724(.a(G1051), .O(gate430inter7));
  inv1  gate2725(.a(G1147), .O(gate430inter8));
  nand2 gate2726(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2727(.a(s_311), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2728(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2729(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2730(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1149(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1150(.a(gate432inter0), .b(s_86), .O(gate432inter1));
  and2  gate1151(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1152(.a(s_86), .O(gate432inter3));
  inv1  gate1153(.a(s_87), .O(gate432inter4));
  nand2 gate1154(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1155(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1156(.a(G1054), .O(gate432inter7));
  inv1  gate1157(.a(G1150), .O(gate432inter8));
  nand2 gate1158(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1159(.a(s_87), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1160(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1161(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1162(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2983(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2984(.a(gate433inter0), .b(s_348), .O(gate433inter1));
  and2  gate2985(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2986(.a(s_348), .O(gate433inter3));
  inv1  gate2987(.a(s_349), .O(gate433inter4));
  nand2 gate2988(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2989(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2990(.a(G8), .O(gate433inter7));
  inv1  gate2991(.a(G1153), .O(gate433inter8));
  nand2 gate2992(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2993(.a(s_349), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2994(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2995(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2996(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2955(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2956(.a(gate435inter0), .b(s_344), .O(gate435inter1));
  and2  gate2957(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2958(.a(s_344), .O(gate435inter3));
  inv1  gate2959(.a(s_345), .O(gate435inter4));
  nand2 gate2960(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2961(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2962(.a(G9), .O(gate435inter7));
  inv1  gate2963(.a(G1156), .O(gate435inter8));
  nand2 gate2964(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2965(.a(s_345), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2966(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2967(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2968(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1191(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1192(.a(gate437inter0), .b(s_92), .O(gate437inter1));
  and2  gate1193(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1194(.a(s_92), .O(gate437inter3));
  inv1  gate1195(.a(s_93), .O(gate437inter4));
  nand2 gate1196(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1197(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1198(.a(G10), .O(gate437inter7));
  inv1  gate1199(.a(G1159), .O(gate437inter8));
  nand2 gate1200(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1201(.a(s_93), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1202(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1203(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1204(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1653(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1654(.a(gate441inter0), .b(s_158), .O(gate441inter1));
  and2  gate1655(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1656(.a(s_158), .O(gate441inter3));
  inv1  gate1657(.a(s_159), .O(gate441inter4));
  nand2 gate1658(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1659(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1660(.a(G12), .O(gate441inter7));
  inv1  gate1661(.a(G1165), .O(gate441inter8));
  nand2 gate1662(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1663(.a(s_159), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1664(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1665(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1666(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2675(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2676(.a(gate442inter0), .b(s_304), .O(gate442inter1));
  and2  gate2677(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2678(.a(s_304), .O(gate442inter3));
  inv1  gate2679(.a(s_305), .O(gate442inter4));
  nand2 gate2680(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2681(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2682(.a(G1069), .O(gate442inter7));
  inv1  gate2683(.a(G1165), .O(gate442inter8));
  nand2 gate2684(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2685(.a(s_305), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2686(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2687(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2688(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1009(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1010(.a(gate443inter0), .b(s_66), .O(gate443inter1));
  and2  gate1011(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1012(.a(s_66), .O(gate443inter3));
  inv1  gate1013(.a(s_67), .O(gate443inter4));
  nand2 gate1014(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1015(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1016(.a(G13), .O(gate443inter7));
  inv1  gate1017(.a(G1168), .O(gate443inter8));
  nand2 gate1018(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1019(.a(s_67), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1020(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1021(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1022(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2563(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2564(.a(gate445inter0), .b(s_288), .O(gate445inter1));
  and2  gate2565(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2566(.a(s_288), .O(gate445inter3));
  inv1  gate2567(.a(s_289), .O(gate445inter4));
  nand2 gate2568(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2569(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2570(.a(G14), .O(gate445inter7));
  inv1  gate2571(.a(G1171), .O(gate445inter8));
  nand2 gate2572(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2573(.a(s_289), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2574(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2575(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2576(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2241(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2242(.a(gate448inter0), .b(s_242), .O(gate448inter1));
  and2  gate2243(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2244(.a(s_242), .O(gate448inter3));
  inv1  gate2245(.a(s_243), .O(gate448inter4));
  nand2 gate2246(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2247(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2248(.a(G1078), .O(gate448inter7));
  inv1  gate2249(.a(G1174), .O(gate448inter8));
  nand2 gate2250(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2251(.a(s_243), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2252(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2253(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2254(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1877(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1878(.a(gate450inter0), .b(s_190), .O(gate450inter1));
  and2  gate1879(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1880(.a(s_190), .O(gate450inter3));
  inv1  gate1881(.a(s_191), .O(gate450inter4));
  nand2 gate1882(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1883(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1884(.a(G1081), .O(gate450inter7));
  inv1  gate1885(.a(G1177), .O(gate450inter8));
  nand2 gate1886(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1887(.a(s_191), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1888(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1889(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1890(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate547(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate548(.a(gate453inter0), .b(s_0), .O(gate453inter1));
  and2  gate549(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate550(.a(s_0), .O(gate453inter3));
  inv1  gate551(.a(s_1), .O(gate453inter4));
  nand2 gate552(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate553(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate554(.a(G18), .O(gate453inter7));
  inv1  gate555(.a(G1183), .O(gate453inter8));
  nand2 gate556(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate557(.a(s_1), .b(gate453inter3), .O(gate453inter10));
  nor2  gate558(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate559(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate560(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1989(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1990(.a(gate454inter0), .b(s_206), .O(gate454inter1));
  and2  gate1991(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1992(.a(s_206), .O(gate454inter3));
  inv1  gate1993(.a(s_207), .O(gate454inter4));
  nand2 gate1994(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1995(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1996(.a(G1087), .O(gate454inter7));
  inv1  gate1997(.a(G1183), .O(gate454inter8));
  nand2 gate1998(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1999(.a(s_207), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2000(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2001(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2002(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate743(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate744(.a(gate455inter0), .b(s_28), .O(gate455inter1));
  and2  gate745(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate746(.a(s_28), .O(gate455inter3));
  inv1  gate747(.a(s_29), .O(gate455inter4));
  nand2 gate748(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate749(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate750(.a(G19), .O(gate455inter7));
  inv1  gate751(.a(G1186), .O(gate455inter8));
  nand2 gate752(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate753(.a(s_29), .b(gate455inter3), .O(gate455inter10));
  nor2  gate754(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate755(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate756(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1121(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1122(.a(gate456inter0), .b(s_82), .O(gate456inter1));
  and2  gate1123(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1124(.a(s_82), .O(gate456inter3));
  inv1  gate1125(.a(s_83), .O(gate456inter4));
  nand2 gate1126(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1127(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1128(.a(G1090), .O(gate456inter7));
  inv1  gate1129(.a(G1186), .O(gate456inter8));
  nand2 gate1130(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1131(.a(s_83), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1132(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1133(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1134(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1401(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1402(.a(gate458inter0), .b(s_122), .O(gate458inter1));
  and2  gate1403(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1404(.a(s_122), .O(gate458inter3));
  inv1  gate1405(.a(s_123), .O(gate458inter4));
  nand2 gate1406(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1407(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1408(.a(G1093), .O(gate458inter7));
  inv1  gate1409(.a(G1189), .O(gate458inter8));
  nand2 gate1410(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1411(.a(s_123), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1412(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1413(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1414(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1093(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1094(.a(gate461inter0), .b(s_78), .O(gate461inter1));
  and2  gate1095(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1096(.a(s_78), .O(gate461inter3));
  inv1  gate1097(.a(s_79), .O(gate461inter4));
  nand2 gate1098(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1099(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1100(.a(G22), .O(gate461inter7));
  inv1  gate1101(.a(G1195), .O(gate461inter8));
  nand2 gate1102(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1103(.a(s_79), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1104(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1105(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1106(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2619(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2620(.a(gate462inter0), .b(s_296), .O(gate462inter1));
  and2  gate2621(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2622(.a(s_296), .O(gate462inter3));
  inv1  gate2623(.a(s_297), .O(gate462inter4));
  nand2 gate2624(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2625(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2626(.a(G1099), .O(gate462inter7));
  inv1  gate2627(.a(G1195), .O(gate462inter8));
  nand2 gate2628(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2629(.a(s_297), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2630(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2631(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2632(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate3193(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate3194(.a(gate464inter0), .b(s_378), .O(gate464inter1));
  and2  gate3195(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate3196(.a(s_378), .O(gate464inter3));
  inv1  gate3197(.a(s_379), .O(gate464inter4));
  nand2 gate3198(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate3199(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate3200(.a(G1102), .O(gate464inter7));
  inv1  gate3201(.a(G1198), .O(gate464inter8));
  nand2 gate3202(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate3203(.a(s_379), .b(gate464inter3), .O(gate464inter10));
  nor2  gate3204(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate3205(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate3206(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1065(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1066(.a(gate465inter0), .b(s_74), .O(gate465inter1));
  and2  gate1067(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1068(.a(s_74), .O(gate465inter3));
  inv1  gate1069(.a(s_75), .O(gate465inter4));
  nand2 gate1070(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1071(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1072(.a(G24), .O(gate465inter7));
  inv1  gate1073(.a(G1201), .O(gate465inter8));
  nand2 gate1074(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1075(.a(s_75), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1076(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1077(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1078(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1905(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1906(.a(gate469inter0), .b(s_194), .O(gate469inter1));
  and2  gate1907(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1908(.a(s_194), .O(gate469inter3));
  inv1  gate1909(.a(s_195), .O(gate469inter4));
  nand2 gate1910(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1911(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1912(.a(G26), .O(gate469inter7));
  inv1  gate1913(.a(G1207), .O(gate469inter8));
  nand2 gate1914(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1915(.a(s_195), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1916(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1917(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1918(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate575(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate576(.a(gate471inter0), .b(s_4), .O(gate471inter1));
  and2  gate577(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate578(.a(s_4), .O(gate471inter3));
  inv1  gate579(.a(s_5), .O(gate471inter4));
  nand2 gate580(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate581(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate582(.a(G27), .O(gate471inter7));
  inv1  gate583(.a(G1210), .O(gate471inter8));
  nand2 gate584(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate585(.a(s_5), .b(gate471inter3), .O(gate471inter10));
  nor2  gate586(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate587(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate588(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1681(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1682(.a(gate476inter0), .b(s_162), .O(gate476inter1));
  and2  gate1683(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1684(.a(s_162), .O(gate476inter3));
  inv1  gate1685(.a(s_163), .O(gate476inter4));
  nand2 gate1686(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1687(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1688(.a(G1120), .O(gate476inter7));
  inv1  gate1689(.a(G1216), .O(gate476inter8));
  nand2 gate1690(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1691(.a(s_163), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1692(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1693(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1694(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1737(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1738(.a(gate479inter0), .b(s_170), .O(gate479inter1));
  and2  gate1739(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1740(.a(s_170), .O(gate479inter3));
  inv1  gate1741(.a(s_171), .O(gate479inter4));
  nand2 gate1742(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1743(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1744(.a(G31), .O(gate479inter7));
  inv1  gate1745(.a(G1222), .O(gate479inter8));
  nand2 gate1746(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1747(.a(s_171), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1748(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1749(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1750(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1863(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1864(.a(gate482inter0), .b(s_188), .O(gate482inter1));
  and2  gate1865(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1866(.a(s_188), .O(gate482inter3));
  inv1  gate1867(.a(s_189), .O(gate482inter4));
  nand2 gate1868(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1869(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1870(.a(G1129), .O(gate482inter7));
  inv1  gate1871(.a(G1225), .O(gate482inter8));
  nand2 gate1872(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1873(.a(s_189), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1874(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1875(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1876(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate645(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate646(.a(gate485inter0), .b(s_14), .O(gate485inter1));
  and2  gate647(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate648(.a(s_14), .O(gate485inter3));
  inv1  gate649(.a(s_15), .O(gate485inter4));
  nand2 gate650(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate651(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate652(.a(G1232), .O(gate485inter7));
  inv1  gate653(.a(G1233), .O(gate485inter8));
  nand2 gate654(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate655(.a(s_15), .b(gate485inter3), .O(gate485inter10));
  nor2  gate656(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate657(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate658(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2269(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2270(.a(gate490inter0), .b(s_246), .O(gate490inter1));
  and2  gate2271(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2272(.a(s_246), .O(gate490inter3));
  inv1  gate2273(.a(s_247), .O(gate490inter4));
  nand2 gate2274(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2275(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2276(.a(G1242), .O(gate490inter7));
  inv1  gate2277(.a(G1243), .O(gate490inter8));
  nand2 gate2278(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2279(.a(s_247), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2280(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2281(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2282(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2101(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2102(.a(gate492inter0), .b(s_222), .O(gate492inter1));
  and2  gate2103(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2104(.a(s_222), .O(gate492inter3));
  inv1  gate2105(.a(s_223), .O(gate492inter4));
  nand2 gate2106(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2107(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2108(.a(G1246), .O(gate492inter7));
  inv1  gate2109(.a(G1247), .O(gate492inter8));
  nand2 gate2110(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2111(.a(s_223), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2112(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2113(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2114(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate855(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate856(.a(gate493inter0), .b(s_44), .O(gate493inter1));
  and2  gate857(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate858(.a(s_44), .O(gate493inter3));
  inv1  gate859(.a(s_45), .O(gate493inter4));
  nand2 gate860(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate861(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate862(.a(G1248), .O(gate493inter7));
  inv1  gate863(.a(G1249), .O(gate493inter8));
  nand2 gate864(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate865(.a(s_45), .b(gate493inter3), .O(gate493inter10));
  nor2  gate866(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate867(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate868(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1429(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1430(.a(gate494inter0), .b(s_126), .O(gate494inter1));
  and2  gate1431(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1432(.a(s_126), .O(gate494inter3));
  inv1  gate1433(.a(s_127), .O(gate494inter4));
  nand2 gate1434(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1435(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1436(.a(G1250), .O(gate494inter7));
  inv1  gate1437(.a(G1251), .O(gate494inter8));
  nand2 gate1438(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1439(.a(s_127), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1440(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1441(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1442(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2409(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2410(.a(gate497inter0), .b(s_266), .O(gate497inter1));
  and2  gate2411(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2412(.a(s_266), .O(gate497inter3));
  inv1  gate2413(.a(s_267), .O(gate497inter4));
  nand2 gate2414(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2415(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2416(.a(G1256), .O(gate497inter7));
  inv1  gate2417(.a(G1257), .O(gate497inter8));
  nand2 gate2418(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2419(.a(s_267), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2420(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2421(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2422(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1919(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1920(.a(gate500inter0), .b(s_196), .O(gate500inter1));
  and2  gate1921(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1922(.a(s_196), .O(gate500inter3));
  inv1  gate1923(.a(s_197), .O(gate500inter4));
  nand2 gate1924(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1925(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1926(.a(G1262), .O(gate500inter7));
  inv1  gate1927(.a(G1263), .O(gate500inter8));
  nand2 gate1928(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1929(.a(s_197), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1930(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1931(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1932(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1135(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1136(.a(gate501inter0), .b(s_84), .O(gate501inter1));
  and2  gate1137(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1138(.a(s_84), .O(gate501inter3));
  inv1  gate1139(.a(s_85), .O(gate501inter4));
  nand2 gate1140(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1141(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1142(.a(G1264), .O(gate501inter7));
  inv1  gate1143(.a(G1265), .O(gate501inter8));
  nand2 gate1144(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1145(.a(s_85), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1146(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1147(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1148(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1513(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1514(.a(gate502inter0), .b(s_138), .O(gate502inter1));
  and2  gate1515(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1516(.a(s_138), .O(gate502inter3));
  inv1  gate1517(.a(s_139), .O(gate502inter4));
  nand2 gate1518(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1519(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1520(.a(G1266), .O(gate502inter7));
  inv1  gate1521(.a(G1267), .O(gate502inter8));
  nand2 gate1522(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1523(.a(s_139), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1524(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1525(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1526(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1373(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1374(.a(gate503inter0), .b(s_118), .O(gate503inter1));
  and2  gate1375(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1376(.a(s_118), .O(gate503inter3));
  inv1  gate1377(.a(s_119), .O(gate503inter4));
  nand2 gate1378(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1379(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1380(.a(G1268), .O(gate503inter7));
  inv1  gate1381(.a(G1269), .O(gate503inter8));
  nand2 gate1382(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1383(.a(s_119), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1384(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1385(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1386(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2647(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2648(.a(gate504inter0), .b(s_300), .O(gate504inter1));
  and2  gate2649(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2650(.a(s_300), .O(gate504inter3));
  inv1  gate2651(.a(s_301), .O(gate504inter4));
  nand2 gate2652(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2653(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2654(.a(G1270), .O(gate504inter7));
  inv1  gate2655(.a(G1271), .O(gate504inter8));
  nand2 gate2656(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2657(.a(s_301), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2658(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2659(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2660(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1177(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1178(.a(gate506inter0), .b(s_90), .O(gate506inter1));
  and2  gate1179(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1180(.a(s_90), .O(gate506inter3));
  inv1  gate1181(.a(s_91), .O(gate506inter4));
  nand2 gate1182(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1183(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1184(.a(G1274), .O(gate506inter7));
  inv1  gate1185(.a(G1275), .O(gate506inter8));
  nand2 gate1186(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1187(.a(s_91), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1188(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1189(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1190(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2871(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2872(.a(gate509inter0), .b(s_332), .O(gate509inter1));
  and2  gate2873(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2874(.a(s_332), .O(gate509inter3));
  inv1  gate2875(.a(s_333), .O(gate509inter4));
  nand2 gate2876(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2877(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2878(.a(G1280), .O(gate509inter7));
  inv1  gate2879(.a(G1281), .O(gate509inter8));
  nand2 gate2880(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2881(.a(s_333), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2882(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2883(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2884(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate3249(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate3250(.a(gate511inter0), .b(s_386), .O(gate511inter1));
  and2  gate3251(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate3252(.a(s_386), .O(gate511inter3));
  inv1  gate3253(.a(s_387), .O(gate511inter4));
  nand2 gate3254(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate3255(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate3256(.a(G1284), .O(gate511inter7));
  inv1  gate3257(.a(G1285), .O(gate511inter8));
  nand2 gate3258(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate3259(.a(s_387), .b(gate511inter3), .O(gate511inter10));
  nor2  gate3260(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate3261(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate3262(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate995(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate996(.a(gate513inter0), .b(s_64), .O(gate513inter1));
  and2  gate997(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate998(.a(s_64), .O(gate513inter3));
  inv1  gate999(.a(s_65), .O(gate513inter4));
  nand2 gate1000(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1001(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1002(.a(G1288), .O(gate513inter7));
  inv1  gate1003(.a(G1289), .O(gate513inter8));
  nand2 gate1004(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1005(.a(s_65), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1006(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1007(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1008(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule