module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate7inter0, gate7inter1, gate7inter2, gate7inter3, gate7inter4, gate7inter5, gate7inter6, gate7inter7, gate7inter8, gate7inter9, gate7inter10, gate7inter11, gate7inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate231(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate232(.a(gate3inter0), .b(s_4), .O(gate3inter1));
  and2  gate233(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate234(.a(s_4), .O(gate3inter3));
  inv1  gate235(.a(s_5), .O(gate3inter4));
  nand2 gate236(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate237(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate238(.a(N17), .O(gate3inter7));
  inv1  gate239(.a(N21), .O(gate3inter8));
  nand2 gate240(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate241(.a(s_5), .b(gate3inter3), .O(gate3inter10));
  nor2  gate242(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate243(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate244(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate329(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate330(.a(gate6inter0), .b(s_18), .O(gate6inter1));
  and2  gate331(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate332(.a(s_18), .O(gate6inter3));
  inv1  gate333(.a(s_19), .O(gate6inter4));
  nand2 gate334(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate335(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate336(.a(N41), .O(gate6inter7));
  inv1  gate337(.a(N45), .O(gate6inter8));
  nand2 gate338(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate339(.a(s_19), .b(gate6inter3), .O(gate6inter10));
  nor2  gate340(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate341(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate342(.a(gate6inter12), .b(gate6inter1), .O(N255));

  xor2  gate413(.a(N53), .b(N49), .O(gate7inter0));
  nand2 gate414(.a(gate7inter0), .b(s_30), .O(gate7inter1));
  and2  gate415(.a(N53), .b(N49), .O(gate7inter2));
  inv1  gate416(.a(s_30), .O(gate7inter3));
  inv1  gate417(.a(s_31), .O(gate7inter4));
  nand2 gate418(.a(gate7inter4), .b(gate7inter3), .O(gate7inter5));
  nor2  gate419(.a(gate7inter5), .b(gate7inter2), .O(gate7inter6));
  inv1  gate420(.a(N49), .O(gate7inter7));
  inv1  gate421(.a(N53), .O(gate7inter8));
  nand2 gate422(.a(gate7inter8), .b(gate7inter7), .O(gate7inter9));
  nand2 gate423(.a(s_31), .b(gate7inter3), .O(gate7inter10));
  nor2  gate424(.a(gate7inter10), .b(gate7inter9), .O(gate7inter11));
  nor2  gate425(.a(gate7inter11), .b(gate7inter6), .O(gate7inter12));
  nand2 gate426(.a(gate7inter12), .b(gate7inter1), .O(N256));
xor2 gate8( .a(N57), .b(N61), .O(N257) );

  xor2  gate287(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate288(.a(gate9inter0), .b(s_12), .O(gate9inter1));
  and2  gate289(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate290(.a(s_12), .O(gate9inter3));
  inv1  gate291(.a(s_13), .O(gate9inter4));
  nand2 gate292(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate293(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate294(.a(N65), .O(gate9inter7));
  inv1  gate295(.a(N69), .O(gate9inter8));
  nand2 gate296(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate297(.a(s_13), .b(gate9inter3), .O(gate9inter10));
  nor2  gate298(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate299(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate300(.a(gate9inter12), .b(gate9inter1), .O(N258));
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );

  xor2  gate217(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate218(.a(gate13inter0), .b(s_2), .O(gate13inter1));
  and2  gate219(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate220(.a(s_2), .O(gate13inter3));
  inv1  gate221(.a(s_3), .O(gate13inter4));
  nand2 gate222(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate223(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate224(.a(N97), .O(gate13inter7));
  inv1  gate225(.a(N101), .O(gate13inter8));
  nand2 gate226(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate227(.a(s_3), .b(gate13inter3), .O(gate13inter10));
  nor2  gate228(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate229(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate230(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );

  xor2  gate371(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate372(.a(gate15inter0), .b(s_24), .O(gate15inter1));
  and2  gate373(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate374(.a(s_24), .O(gate15inter3));
  inv1  gate375(.a(s_25), .O(gate15inter4));
  nand2 gate376(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate377(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate378(.a(N113), .O(gate15inter7));
  inv1  gate379(.a(N117), .O(gate15inter8));
  nand2 gate380(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate381(.a(s_25), .b(gate15inter3), .O(gate15inter10));
  nor2  gate382(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate383(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate384(.a(gate15inter12), .b(gate15inter1), .O(N264));
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate301(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate302(.a(gate25inter0), .b(s_14), .O(gate25inter1));
  and2  gate303(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate304(.a(s_14), .O(gate25inter3));
  inv1  gate305(.a(s_15), .O(gate25inter4));
  nand2 gate306(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate307(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate308(.a(N1), .O(gate25inter7));
  inv1  gate309(.a(N17), .O(gate25inter8));
  nand2 gate310(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate311(.a(s_15), .b(gate25inter3), .O(gate25inter10));
  nor2  gate312(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate313(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate314(.a(gate25inter12), .b(gate25inter1), .O(N274));

  xor2  gate259(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate260(.a(gate26inter0), .b(s_8), .O(gate26inter1));
  and2  gate261(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate262(.a(s_8), .O(gate26inter3));
  inv1  gate263(.a(s_9), .O(gate26inter4));
  nand2 gate264(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate265(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate266(.a(N33), .O(gate26inter7));
  inv1  gate267(.a(N49), .O(gate26inter8));
  nand2 gate268(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate269(.a(s_9), .b(gate26inter3), .O(gate26inter10));
  nor2  gate270(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate271(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate272(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate315(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate316(.a(gate55inter0), .b(s_16), .O(gate55inter1));
  and2  gate317(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate318(.a(s_16), .O(gate55inter3));
  inv1  gate319(.a(s_17), .O(gate55inter4));
  nand2 gate320(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate321(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate322(.a(N286), .O(gate55inter7));
  inv1  gate323(.a(N287), .O(gate55inter8));
  nand2 gate324(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate325(.a(s_17), .b(gate55inter3), .O(gate55inter10));
  nor2  gate326(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate327(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate328(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate385(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate386(.a(gate59inter0), .b(s_26), .O(gate59inter1));
  and2  gate387(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate388(.a(s_26), .O(gate59inter3));
  inv1  gate389(.a(s_27), .O(gate59inter4));
  nand2 gate390(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate391(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate392(.a(N290), .O(gate59inter7));
  inv1  gate393(.a(N296), .O(gate59inter8));
  nand2 gate394(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate395(.a(s_27), .b(gate59inter3), .O(gate59inter10));
  nor2  gate396(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate397(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate398(.a(gate59inter12), .b(gate59inter1), .O(N340));
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );

  xor2  gate399(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate400(.a(gate63inter0), .b(s_28), .O(gate63inter1));
  and2  gate401(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate402(.a(s_28), .O(gate63inter3));
  inv1  gate403(.a(s_29), .O(gate63inter4));
  nand2 gate404(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate405(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate406(.a(N302), .O(gate63inter7));
  inv1  gate407(.a(N308), .O(gate63inter8));
  nand2 gate408(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate409(.a(s_29), .b(gate63inter3), .O(gate63inter10));
  nor2  gate410(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate411(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate412(.a(gate63inter12), .b(gate63inter1), .O(N344));
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );

  xor2  gate273(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate274(.a(gate66inter0), .b(s_10), .O(gate66inter1));
  and2  gate275(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate276(.a(s_10), .O(gate66inter3));
  inv1  gate277(.a(s_11), .O(gate66inter4));
  nand2 gate278(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate279(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate280(.a(N267), .O(gate66inter7));
  inv1  gate281(.a(N343), .O(gate66inter8));
  nand2 gate282(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate283(.a(s_11), .b(gate66inter3), .O(gate66inter10));
  nor2  gate284(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate285(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate286(.a(gate66inter12), .b(gate66inter1), .O(N347));
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate245(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate246(.a(gate176inter0), .b(s_6), .O(gate176inter1));
  and2  gate247(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate248(.a(s_6), .O(gate176inter3));
  inv1  gate249(.a(s_7), .O(gate176inter4));
  nand2 gate250(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate251(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate252(.a(N21), .O(gate176inter7));
  inv1  gate253(.a(N697), .O(gate176inter8));
  nand2 gate254(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate255(.a(s_7), .b(gate176inter3), .O(gate176inter10));
  nor2  gate256(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate257(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate258(.a(gate176inter12), .b(gate176inter1), .O(N729));
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );

  xor2  gate357(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate358(.a(gate181inter0), .b(s_22), .O(gate181inter1));
  and2  gate359(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate360(.a(s_22), .O(gate181inter3));
  inv1  gate361(.a(s_23), .O(gate181inter4));
  nand2 gate362(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate363(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate364(.a(N41), .O(gate181inter7));
  inv1  gate365(.a(N702), .O(gate181inter8));
  nand2 gate366(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate367(.a(s_23), .b(gate181inter3), .O(gate181inter10));
  nor2  gate368(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate369(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate370(.a(gate181inter12), .b(gate181inter1), .O(N734));
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );

  xor2  gate203(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate204(.a(gate190inter0), .b(s_0), .O(gate190inter1));
  and2  gate205(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate206(.a(s_0), .O(gate190inter3));
  inv1  gate207(.a(s_1), .O(gate190inter4));
  nand2 gate208(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate209(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate210(.a(N77), .O(gate190inter7));
  inv1  gate211(.a(N711), .O(gate190inter8));
  nand2 gate212(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate213(.a(s_1), .b(gate190inter3), .O(gate190inter10));
  nor2  gate214(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate215(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate216(.a(gate190inter12), .b(gate190inter1), .O(N743));
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate343(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate344(.a(gate201inter0), .b(s_20), .O(gate201inter1));
  and2  gate345(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate346(.a(s_20), .O(gate201inter3));
  inv1  gate347(.a(s_21), .O(gate201inter4));
  nand2 gate348(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate349(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate350(.a(N121), .O(gate201inter7));
  inv1  gate351(.a(N722), .O(gate201inter8));
  nand2 gate352(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate353(.a(s_21), .b(gate201inter3), .O(gate201inter10));
  nor2  gate354(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate355(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate356(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule