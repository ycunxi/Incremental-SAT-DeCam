module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1261(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1262(.a(gate9inter0), .b(s_102), .O(gate9inter1));
  and2  gate1263(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1264(.a(s_102), .O(gate9inter3));
  inv1  gate1265(.a(s_103), .O(gate9inter4));
  nand2 gate1266(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1267(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1268(.a(G1), .O(gate9inter7));
  inv1  gate1269(.a(G2), .O(gate9inter8));
  nand2 gate1270(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1271(.a(s_103), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1272(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1273(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1274(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1163(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1164(.a(gate12inter0), .b(s_88), .O(gate12inter1));
  and2  gate1165(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1166(.a(s_88), .O(gate12inter3));
  inv1  gate1167(.a(s_89), .O(gate12inter4));
  nand2 gate1168(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1169(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1170(.a(G7), .O(gate12inter7));
  inv1  gate1171(.a(G8), .O(gate12inter8));
  nand2 gate1172(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1173(.a(s_89), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1174(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1175(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1176(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1611(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1612(.a(gate13inter0), .b(s_152), .O(gate13inter1));
  and2  gate1613(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1614(.a(s_152), .O(gate13inter3));
  inv1  gate1615(.a(s_153), .O(gate13inter4));
  nand2 gate1616(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1617(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1618(.a(G9), .O(gate13inter7));
  inv1  gate1619(.a(G10), .O(gate13inter8));
  nand2 gate1620(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1621(.a(s_153), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1622(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1623(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1624(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1513(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1514(.a(gate15inter0), .b(s_138), .O(gate15inter1));
  and2  gate1515(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1516(.a(s_138), .O(gate15inter3));
  inv1  gate1517(.a(s_139), .O(gate15inter4));
  nand2 gate1518(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1519(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1520(.a(G13), .O(gate15inter7));
  inv1  gate1521(.a(G14), .O(gate15inter8));
  nand2 gate1522(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1523(.a(s_139), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1524(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1525(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1526(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate995(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate996(.a(gate17inter0), .b(s_64), .O(gate17inter1));
  and2  gate997(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate998(.a(s_64), .O(gate17inter3));
  inv1  gate999(.a(s_65), .O(gate17inter4));
  nand2 gate1000(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1001(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1002(.a(G17), .O(gate17inter7));
  inv1  gate1003(.a(G18), .O(gate17inter8));
  nand2 gate1004(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1005(.a(s_65), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1006(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1007(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1008(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1723(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1724(.a(gate19inter0), .b(s_168), .O(gate19inter1));
  and2  gate1725(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1726(.a(s_168), .O(gate19inter3));
  inv1  gate1727(.a(s_169), .O(gate19inter4));
  nand2 gate1728(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1729(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1730(.a(G21), .O(gate19inter7));
  inv1  gate1731(.a(G22), .O(gate19inter8));
  nand2 gate1732(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1733(.a(s_169), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1734(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1735(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1736(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate617(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate618(.a(gate30inter0), .b(s_10), .O(gate30inter1));
  and2  gate619(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate620(.a(s_10), .O(gate30inter3));
  inv1  gate621(.a(s_11), .O(gate30inter4));
  nand2 gate622(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate623(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate624(.a(G11), .O(gate30inter7));
  inv1  gate625(.a(G15), .O(gate30inter8));
  nand2 gate626(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate627(.a(s_11), .b(gate30inter3), .O(gate30inter10));
  nor2  gate628(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate629(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate630(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate603(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate604(.a(gate31inter0), .b(s_8), .O(gate31inter1));
  and2  gate605(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate606(.a(s_8), .O(gate31inter3));
  inv1  gate607(.a(s_9), .O(gate31inter4));
  nand2 gate608(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate609(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate610(.a(G4), .O(gate31inter7));
  inv1  gate611(.a(G8), .O(gate31inter8));
  nand2 gate612(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate613(.a(s_9), .b(gate31inter3), .O(gate31inter10));
  nor2  gate614(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate615(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate616(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate659(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate660(.a(gate32inter0), .b(s_16), .O(gate32inter1));
  and2  gate661(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate662(.a(s_16), .O(gate32inter3));
  inv1  gate663(.a(s_17), .O(gate32inter4));
  nand2 gate664(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate665(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate666(.a(G12), .O(gate32inter7));
  inv1  gate667(.a(G16), .O(gate32inter8));
  nand2 gate668(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate669(.a(s_17), .b(gate32inter3), .O(gate32inter10));
  nor2  gate670(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate671(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate672(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate715(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate716(.a(gate36inter0), .b(s_24), .O(gate36inter1));
  and2  gate717(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate718(.a(s_24), .O(gate36inter3));
  inv1  gate719(.a(s_25), .O(gate36inter4));
  nand2 gate720(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate721(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate722(.a(G26), .O(gate36inter7));
  inv1  gate723(.a(G30), .O(gate36inter8));
  nand2 gate724(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate725(.a(s_25), .b(gate36inter3), .O(gate36inter10));
  nor2  gate726(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate727(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate728(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1359(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1360(.a(gate38inter0), .b(s_116), .O(gate38inter1));
  and2  gate1361(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1362(.a(s_116), .O(gate38inter3));
  inv1  gate1363(.a(s_117), .O(gate38inter4));
  nand2 gate1364(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1365(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1366(.a(G27), .O(gate38inter7));
  inv1  gate1367(.a(G31), .O(gate38inter8));
  nand2 gate1368(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1369(.a(s_117), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1370(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1371(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1372(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1443(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1444(.a(gate42inter0), .b(s_128), .O(gate42inter1));
  and2  gate1445(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1446(.a(s_128), .O(gate42inter3));
  inv1  gate1447(.a(s_129), .O(gate42inter4));
  nand2 gate1448(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1449(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1450(.a(G2), .O(gate42inter7));
  inv1  gate1451(.a(G266), .O(gate42inter8));
  nand2 gate1452(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1453(.a(s_129), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1454(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1455(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1456(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate813(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate814(.a(gate50inter0), .b(s_38), .O(gate50inter1));
  and2  gate815(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate816(.a(s_38), .O(gate50inter3));
  inv1  gate817(.a(s_39), .O(gate50inter4));
  nand2 gate818(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate819(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate820(.a(G10), .O(gate50inter7));
  inv1  gate821(.a(G278), .O(gate50inter8));
  nand2 gate822(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate823(.a(s_39), .b(gate50inter3), .O(gate50inter10));
  nor2  gate824(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate825(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate826(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate771(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate772(.a(gate51inter0), .b(s_32), .O(gate51inter1));
  and2  gate773(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate774(.a(s_32), .O(gate51inter3));
  inv1  gate775(.a(s_33), .O(gate51inter4));
  nand2 gate776(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate777(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate778(.a(G11), .O(gate51inter7));
  inv1  gate779(.a(G281), .O(gate51inter8));
  nand2 gate780(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate781(.a(s_33), .b(gate51inter3), .O(gate51inter10));
  nor2  gate782(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate783(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate784(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate981(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate982(.a(gate52inter0), .b(s_62), .O(gate52inter1));
  and2  gate983(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate984(.a(s_62), .O(gate52inter3));
  inv1  gate985(.a(s_63), .O(gate52inter4));
  nand2 gate986(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate987(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate988(.a(G12), .O(gate52inter7));
  inv1  gate989(.a(G281), .O(gate52inter8));
  nand2 gate990(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate991(.a(s_63), .b(gate52inter3), .O(gate52inter10));
  nor2  gate992(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate993(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate994(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1205(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1206(.a(gate58inter0), .b(s_94), .O(gate58inter1));
  and2  gate1207(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1208(.a(s_94), .O(gate58inter3));
  inv1  gate1209(.a(s_95), .O(gate58inter4));
  nand2 gate1210(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1211(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1212(.a(G18), .O(gate58inter7));
  inv1  gate1213(.a(G290), .O(gate58inter8));
  nand2 gate1214(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1215(.a(s_95), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1216(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1217(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1218(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1289(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1290(.a(gate59inter0), .b(s_106), .O(gate59inter1));
  and2  gate1291(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1292(.a(s_106), .O(gate59inter3));
  inv1  gate1293(.a(s_107), .O(gate59inter4));
  nand2 gate1294(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1295(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1296(.a(G19), .O(gate59inter7));
  inv1  gate1297(.a(G293), .O(gate59inter8));
  nand2 gate1298(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1299(.a(s_107), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1300(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1301(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1302(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1695(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1696(.a(gate66inter0), .b(s_164), .O(gate66inter1));
  and2  gate1697(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1698(.a(s_164), .O(gate66inter3));
  inv1  gate1699(.a(s_165), .O(gate66inter4));
  nand2 gate1700(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1701(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1702(.a(G26), .O(gate66inter7));
  inv1  gate1703(.a(G302), .O(gate66inter8));
  nand2 gate1704(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1705(.a(s_165), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1706(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1707(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1708(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1597(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1598(.a(gate69inter0), .b(s_150), .O(gate69inter1));
  and2  gate1599(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1600(.a(s_150), .O(gate69inter3));
  inv1  gate1601(.a(s_151), .O(gate69inter4));
  nand2 gate1602(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1603(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1604(.a(G29), .O(gate69inter7));
  inv1  gate1605(.a(G308), .O(gate69inter8));
  nand2 gate1606(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1607(.a(s_151), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1608(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1609(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1610(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate967(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate968(.a(gate84inter0), .b(s_60), .O(gate84inter1));
  and2  gate969(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate970(.a(s_60), .O(gate84inter3));
  inv1  gate971(.a(s_61), .O(gate84inter4));
  nand2 gate972(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate973(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate974(.a(G15), .O(gate84inter7));
  inv1  gate975(.a(G329), .O(gate84inter8));
  nand2 gate976(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate977(.a(s_61), .b(gate84inter3), .O(gate84inter10));
  nor2  gate978(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate979(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate980(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1751(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1752(.a(gate90inter0), .b(s_172), .O(gate90inter1));
  and2  gate1753(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1754(.a(s_172), .O(gate90inter3));
  inv1  gate1755(.a(s_173), .O(gate90inter4));
  nand2 gate1756(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1757(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1758(.a(G21), .O(gate90inter7));
  inv1  gate1759(.a(G338), .O(gate90inter8));
  nand2 gate1760(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1761(.a(s_173), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1762(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1763(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1764(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate673(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate674(.a(gate91inter0), .b(s_18), .O(gate91inter1));
  and2  gate675(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate676(.a(s_18), .O(gate91inter3));
  inv1  gate677(.a(s_19), .O(gate91inter4));
  nand2 gate678(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate679(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate680(.a(G25), .O(gate91inter7));
  inv1  gate681(.a(G341), .O(gate91inter8));
  nand2 gate682(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate683(.a(s_19), .b(gate91inter3), .O(gate91inter10));
  nor2  gate684(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate685(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate686(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1093(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1094(.a(gate96inter0), .b(s_78), .O(gate96inter1));
  and2  gate1095(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1096(.a(s_78), .O(gate96inter3));
  inv1  gate1097(.a(s_79), .O(gate96inter4));
  nand2 gate1098(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1099(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1100(.a(G30), .O(gate96inter7));
  inv1  gate1101(.a(G347), .O(gate96inter8));
  nand2 gate1102(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1103(.a(s_79), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1104(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1105(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1106(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1345(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1346(.a(gate98inter0), .b(s_114), .O(gate98inter1));
  and2  gate1347(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1348(.a(s_114), .O(gate98inter3));
  inv1  gate1349(.a(s_115), .O(gate98inter4));
  nand2 gate1350(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1351(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1352(.a(G23), .O(gate98inter7));
  inv1  gate1353(.a(G350), .O(gate98inter8));
  nand2 gate1354(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1355(.a(s_115), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1356(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1357(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1358(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1079(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1080(.a(gate104inter0), .b(s_76), .O(gate104inter1));
  and2  gate1081(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1082(.a(s_76), .O(gate104inter3));
  inv1  gate1083(.a(s_77), .O(gate104inter4));
  nand2 gate1084(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1085(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1086(.a(G32), .O(gate104inter7));
  inv1  gate1087(.a(G359), .O(gate104inter8));
  nand2 gate1088(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1089(.a(s_77), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1090(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1091(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1092(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1219(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1220(.a(gate105inter0), .b(s_96), .O(gate105inter1));
  and2  gate1221(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1222(.a(s_96), .O(gate105inter3));
  inv1  gate1223(.a(s_97), .O(gate105inter4));
  nand2 gate1224(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1225(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1226(.a(G362), .O(gate105inter7));
  inv1  gate1227(.a(G363), .O(gate105inter8));
  nand2 gate1228(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1229(.a(s_97), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1230(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1231(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1232(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1681(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1682(.a(gate114inter0), .b(s_162), .O(gate114inter1));
  and2  gate1683(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1684(.a(s_162), .O(gate114inter3));
  inv1  gate1685(.a(s_163), .O(gate114inter4));
  nand2 gate1686(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1687(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1688(.a(G380), .O(gate114inter7));
  inv1  gate1689(.a(G381), .O(gate114inter8));
  nand2 gate1690(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1691(.a(s_163), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1692(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1693(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1694(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate589(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate590(.a(gate116inter0), .b(s_6), .O(gate116inter1));
  and2  gate591(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate592(.a(s_6), .O(gate116inter3));
  inv1  gate593(.a(s_7), .O(gate116inter4));
  nand2 gate594(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate595(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate596(.a(G384), .O(gate116inter7));
  inv1  gate597(.a(G385), .O(gate116inter8));
  nand2 gate598(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate599(.a(s_7), .b(gate116inter3), .O(gate116inter10));
  nor2  gate600(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate601(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate602(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1149(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1150(.a(gate118inter0), .b(s_86), .O(gate118inter1));
  and2  gate1151(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1152(.a(s_86), .O(gate118inter3));
  inv1  gate1153(.a(s_87), .O(gate118inter4));
  nand2 gate1154(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1155(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1156(.a(G388), .O(gate118inter7));
  inv1  gate1157(.a(G389), .O(gate118inter8));
  nand2 gate1158(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1159(.a(s_87), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1160(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1161(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1162(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate897(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate898(.a(gate125inter0), .b(s_50), .O(gate125inter1));
  and2  gate899(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate900(.a(s_50), .O(gate125inter3));
  inv1  gate901(.a(s_51), .O(gate125inter4));
  nand2 gate902(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate903(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate904(.a(G402), .O(gate125inter7));
  inv1  gate905(.a(G403), .O(gate125inter8));
  nand2 gate906(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate907(.a(s_51), .b(gate125inter3), .O(gate125inter10));
  nor2  gate908(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate909(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate910(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1639(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1640(.a(gate126inter0), .b(s_156), .O(gate126inter1));
  and2  gate1641(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1642(.a(s_156), .O(gate126inter3));
  inv1  gate1643(.a(s_157), .O(gate126inter4));
  nand2 gate1644(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1645(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1646(.a(G404), .O(gate126inter7));
  inv1  gate1647(.a(G405), .O(gate126inter8));
  nand2 gate1648(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1649(.a(s_157), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1650(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1651(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1652(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1121(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1122(.a(gate131inter0), .b(s_82), .O(gate131inter1));
  and2  gate1123(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1124(.a(s_82), .O(gate131inter3));
  inv1  gate1125(.a(s_83), .O(gate131inter4));
  nand2 gate1126(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1127(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1128(.a(G414), .O(gate131inter7));
  inv1  gate1129(.a(G415), .O(gate131inter8));
  nand2 gate1130(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1131(.a(s_83), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1132(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1133(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1134(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate855(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate856(.a(gate132inter0), .b(s_44), .O(gate132inter1));
  and2  gate857(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate858(.a(s_44), .O(gate132inter3));
  inv1  gate859(.a(s_45), .O(gate132inter4));
  nand2 gate860(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate861(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate862(.a(G416), .O(gate132inter7));
  inv1  gate863(.a(G417), .O(gate132inter8));
  nand2 gate864(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate865(.a(s_45), .b(gate132inter3), .O(gate132inter10));
  nor2  gate866(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate867(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate868(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1037(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1038(.a(gate147inter0), .b(s_70), .O(gate147inter1));
  and2  gate1039(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1040(.a(s_70), .O(gate147inter3));
  inv1  gate1041(.a(s_71), .O(gate147inter4));
  nand2 gate1042(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1043(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1044(.a(G486), .O(gate147inter7));
  inv1  gate1045(.a(G489), .O(gate147inter8));
  nand2 gate1046(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1047(.a(s_71), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1048(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1049(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1050(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1009(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1010(.a(gate148inter0), .b(s_66), .O(gate148inter1));
  and2  gate1011(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1012(.a(s_66), .O(gate148inter3));
  inv1  gate1013(.a(s_67), .O(gate148inter4));
  nand2 gate1014(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1015(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1016(.a(G492), .O(gate148inter7));
  inv1  gate1017(.a(G495), .O(gate148inter8));
  nand2 gate1018(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1019(.a(s_67), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1020(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1021(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1022(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate645(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate646(.a(gate150inter0), .b(s_14), .O(gate150inter1));
  and2  gate647(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate648(.a(s_14), .O(gate150inter3));
  inv1  gate649(.a(s_15), .O(gate150inter4));
  nand2 gate650(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate651(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate652(.a(G504), .O(gate150inter7));
  inv1  gate653(.a(G507), .O(gate150inter8));
  nand2 gate654(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate655(.a(s_15), .b(gate150inter3), .O(gate150inter10));
  nor2  gate656(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate657(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate658(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1457(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1458(.a(gate154inter0), .b(s_130), .O(gate154inter1));
  and2  gate1459(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1460(.a(s_130), .O(gate154inter3));
  inv1  gate1461(.a(s_131), .O(gate154inter4));
  nand2 gate1462(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1463(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1464(.a(G429), .O(gate154inter7));
  inv1  gate1465(.a(G522), .O(gate154inter8));
  nand2 gate1466(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1467(.a(s_131), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1468(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1469(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1470(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1541(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1542(.a(gate158inter0), .b(s_142), .O(gate158inter1));
  and2  gate1543(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1544(.a(s_142), .O(gate158inter3));
  inv1  gate1545(.a(s_143), .O(gate158inter4));
  nand2 gate1546(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1547(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1548(.a(G441), .O(gate158inter7));
  inv1  gate1549(.a(G528), .O(gate158inter8));
  nand2 gate1550(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1551(.a(s_143), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1552(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1553(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1554(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate841(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate842(.a(gate161inter0), .b(s_42), .O(gate161inter1));
  and2  gate843(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate844(.a(s_42), .O(gate161inter3));
  inv1  gate845(.a(s_43), .O(gate161inter4));
  nand2 gate846(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate847(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate848(.a(G450), .O(gate161inter7));
  inv1  gate849(.a(G534), .O(gate161inter8));
  nand2 gate850(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate851(.a(s_43), .b(gate161inter3), .O(gate161inter10));
  nor2  gate852(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate853(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate854(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate561(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate562(.a(gate165inter0), .b(s_2), .O(gate165inter1));
  and2  gate563(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate564(.a(s_2), .O(gate165inter3));
  inv1  gate565(.a(s_3), .O(gate165inter4));
  nand2 gate566(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate567(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate568(.a(G462), .O(gate165inter7));
  inv1  gate569(.a(G540), .O(gate165inter8));
  nand2 gate570(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate571(.a(s_3), .b(gate165inter3), .O(gate165inter10));
  nor2  gate572(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate573(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate574(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1051(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1052(.a(gate169inter0), .b(s_72), .O(gate169inter1));
  and2  gate1053(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1054(.a(s_72), .O(gate169inter3));
  inv1  gate1055(.a(s_73), .O(gate169inter4));
  nand2 gate1056(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1057(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1058(.a(G474), .O(gate169inter7));
  inv1  gate1059(.a(G546), .O(gate169inter8));
  nand2 gate1060(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1061(.a(s_73), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1062(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1063(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1064(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1667(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1668(.a(gate176inter0), .b(s_160), .O(gate176inter1));
  and2  gate1669(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1670(.a(s_160), .O(gate176inter3));
  inv1  gate1671(.a(s_161), .O(gate176inter4));
  nand2 gate1672(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1673(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1674(.a(G495), .O(gate176inter7));
  inv1  gate1675(.a(G555), .O(gate176inter8));
  nand2 gate1676(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1677(.a(s_161), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1678(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1679(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1680(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1107(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1108(.a(gate179inter0), .b(s_80), .O(gate179inter1));
  and2  gate1109(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1110(.a(s_80), .O(gate179inter3));
  inv1  gate1111(.a(s_81), .O(gate179inter4));
  nand2 gate1112(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1113(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1114(.a(G504), .O(gate179inter7));
  inv1  gate1115(.a(G561), .O(gate179inter8));
  nand2 gate1116(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1117(.a(s_81), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1118(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1119(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1120(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1023(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1024(.a(gate181inter0), .b(s_68), .O(gate181inter1));
  and2  gate1025(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1026(.a(s_68), .O(gate181inter3));
  inv1  gate1027(.a(s_69), .O(gate181inter4));
  nand2 gate1028(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1029(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1030(.a(G510), .O(gate181inter7));
  inv1  gate1031(.a(G564), .O(gate181inter8));
  nand2 gate1032(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1033(.a(s_69), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1034(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1035(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1036(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1401(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1402(.a(gate193inter0), .b(s_122), .O(gate193inter1));
  and2  gate1403(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1404(.a(s_122), .O(gate193inter3));
  inv1  gate1405(.a(s_123), .O(gate193inter4));
  nand2 gate1406(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1407(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1408(.a(G586), .O(gate193inter7));
  inv1  gate1409(.a(G587), .O(gate193inter8));
  nand2 gate1410(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1411(.a(s_123), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1412(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1413(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1414(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1807(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1808(.a(gate196inter0), .b(s_180), .O(gate196inter1));
  and2  gate1809(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1810(.a(s_180), .O(gate196inter3));
  inv1  gate1811(.a(s_181), .O(gate196inter4));
  nand2 gate1812(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1813(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1814(.a(G592), .O(gate196inter7));
  inv1  gate1815(.a(G593), .O(gate196inter8));
  nand2 gate1816(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1817(.a(s_181), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1818(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1819(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1820(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate799(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate800(.a(gate203inter0), .b(s_36), .O(gate203inter1));
  and2  gate801(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate802(.a(s_36), .O(gate203inter3));
  inv1  gate803(.a(s_37), .O(gate203inter4));
  nand2 gate804(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate805(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate806(.a(G602), .O(gate203inter7));
  inv1  gate807(.a(G612), .O(gate203inter8));
  nand2 gate808(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate809(.a(s_37), .b(gate203inter3), .O(gate203inter10));
  nor2  gate810(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate811(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate812(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1765(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1766(.a(gate205inter0), .b(s_174), .O(gate205inter1));
  and2  gate1767(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1768(.a(s_174), .O(gate205inter3));
  inv1  gate1769(.a(s_175), .O(gate205inter4));
  nand2 gate1770(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1771(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1772(.a(G622), .O(gate205inter7));
  inv1  gate1773(.a(G627), .O(gate205inter8));
  nand2 gate1774(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1775(.a(s_175), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1776(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1777(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1778(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate785(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate786(.a(gate206inter0), .b(s_34), .O(gate206inter1));
  and2  gate787(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate788(.a(s_34), .O(gate206inter3));
  inv1  gate789(.a(s_35), .O(gate206inter4));
  nand2 gate790(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate791(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate792(.a(G632), .O(gate206inter7));
  inv1  gate793(.a(G637), .O(gate206inter8));
  nand2 gate794(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate795(.a(s_35), .b(gate206inter3), .O(gate206inter10));
  nor2  gate796(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate797(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate798(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate729(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate730(.a(gate219inter0), .b(s_26), .O(gate219inter1));
  and2  gate731(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate732(.a(s_26), .O(gate219inter3));
  inv1  gate733(.a(s_27), .O(gate219inter4));
  nand2 gate734(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate735(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate736(.a(G632), .O(gate219inter7));
  inv1  gate737(.a(G681), .O(gate219inter8));
  nand2 gate738(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate739(.a(s_27), .b(gate219inter3), .O(gate219inter10));
  nor2  gate740(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate741(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate742(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1191(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1192(.a(gate223inter0), .b(s_92), .O(gate223inter1));
  and2  gate1193(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1194(.a(s_92), .O(gate223inter3));
  inv1  gate1195(.a(s_93), .O(gate223inter4));
  nand2 gate1196(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1197(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1198(.a(G627), .O(gate223inter7));
  inv1  gate1199(.a(G687), .O(gate223inter8));
  nand2 gate1200(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1201(.a(s_93), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1202(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1203(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1204(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1555(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1556(.a(gate227inter0), .b(s_144), .O(gate227inter1));
  and2  gate1557(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1558(.a(s_144), .O(gate227inter3));
  inv1  gate1559(.a(s_145), .O(gate227inter4));
  nand2 gate1560(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1561(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1562(.a(G694), .O(gate227inter7));
  inv1  gate1563(.a(G695), .O(gate227inter8));
  nand2 gate1564(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1565(.a(s_145), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1566(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1567(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1568(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1317(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1318(.a(gate232inter0), .b(s_110), .O(gate232inter1));
  and2  gate1319(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1320(.a(s_110), .O(gate232inter3));
  inv1  gate1321(.a(s_111), .O(gate232inter4));
  nand2 gate1322(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1323(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1324(.a(G704), .O(gate232inter7));
  inv1  gate1325(.a(G705), .O(gate232inter8));
  nand2 gate1326(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1327(.a(s_111), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1328(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1329(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1330(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1569(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1570(.a(gate236inter0), .b(s_146), .O(gate236inter1));
  and2  gate1571(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1572(.a(s_146), .O(gate236inter3));
  inv1  gate1573(.a(s_147), .O(gate236inter4));
  nand2 gate1574(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1575(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1576(.a(G251), .O(gate236inter7));
  inv1  gate1577(.a(G727), .O(gate236inter8));
  nand2 gate1578(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1579(.a(s_147), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1580(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1581(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1582(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1135(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1136(.a(gate246inter0), .b(s_84), .O(gate246inter1));
  and2  gate1137(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1138(.a(s_84), .O(gate246inter3));
  inv1  gate1139(.a(s_85), .O(gate246inter4));
  nand2 gate1140(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1141(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1142(.a(G724), .O(gate246inter7));
  inv1  gate1143(.a(G736), .O(gate246inter8));
  nand2 gate1144(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1145(.a(s_85), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1146(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1147(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1148(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1415(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1416(.a(gate255inter0), .b(s_124), .O(gate255inter1));
  and2  gate1417(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1418(.a(s_124), .O(gate255inter3));
  inv1  gate1419(.a(s_125), .O(gate255inter4));
  nand2 gate1420(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1421(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1422(.a(G263), .O(gate255inter7));
  inv1  gate1423(.a(G751), .O(gate255inter8));
  nand2 gate1424(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1425(.a(s_125), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1426(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1427(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1428(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1275(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1276(.a(gate259inter0), .b(s_104), .O(gate259inter1));
  and2  gate1277(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1278(.a(s_104), .O(gate259inter3));
  inv1  gate1279(.a(s_105), .O(gate259inter4));
  nand2 gate1280(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1281(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1282(.a(G758), .O(gate259inter7));
  inv1  gate1283(.a(G759), .O(gate259inter8));
  nand2 gate1284(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1285(.a(s_105), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1286(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1287(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1288(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1709(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1710(.a(gate260inter0), .b(s_166), .O(gate260inter1));
  and2  gate1711(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1712(.a(s_166), .O(gate260inter3));
  inv1  gate1713(.a(s_167), .O(gate260inter4));
  nand2 gate1714(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1715(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1716(.a(G760), .O(gate260inter7));
  inv1  gate1717(.a(G761), .O(gate260inter8));
  nand2 gate1718(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1719(.a(s_167), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1720(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1721(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1722(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1779(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1780(.a(gate262inter0), .b(s_176), .O(gate262inter1));
  and2  gate1781(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1782(.a(s_176), .O(gate262inter3));
  inv1  gate1783(.a(s_177), .O(gate262inter4));
  nand2 gate1784(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1785(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1786(.a(G764), .O(gate262inter7));
  inv1  gate1787(.a(G765), .O(gate262inter8));
  nand2 gate1788(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1789(.a(s_177), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1790(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1791(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1792(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate953(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate954(.a(gate265inter0), .b(s_58), .O(gate265inter1));
  and2  gate955(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate956(.a(s_58), .O(gate265inter3));
  inv1  gate957(.a(s_59), .O(gate265inter4));
  nand2 gate958(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate959(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate960(.a(G642), .O(gate265inter7));
  inv1  gate961(.a(G770), .O(gate265inter8));
  nand2 gate962(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate963(.a(s_59), .b(gate265inter3), .O(gate265inter10));
  nor2  gate964(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate965(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate966(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate925(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate926(.a(gate279inter0), .b(s_54), .O(gate279inter1));
  and2  gate927(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate928(.a(s_54), .O(gate279inter3));
  inv1  gate929(.a(s_55), .O(gate279inter4));
  nand2 gate930(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate931(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate932(.a(G651), .O(gate279inter7));
  inv1  gate933(.a(G803), .O(gate279inter8));
  nand2 gate934(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate935(.a(s_55), .b(gate279inter3), .O(gate279inter10));
  nor2  gate936(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate937(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate938(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate575(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate576(.a(gate280inter0), .b(s_4), .O(gate280inter1));
  and2  gate577(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate578(.a(s_4), .O(gate280inter3));
  inv1  gate579(.a(s_5), .O(gate280inter4));
  nand2 gate580(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate581(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate582(.a(G779), .O(gate280inter7));
  inv1  gate583(.a(G803), .O(gate280inter8));
  nand2 gate584(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate585(.a(s_5), .b(gate280inter3), .O(gate280inter10));
  nor2  gate586(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate587(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate588(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1583(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1584(.a(gate282inter0), .b(s_148), .O(gate282inter1));
  and2  gate1585(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1586(.a(s_148), .O(gate282inter3));
  inv1  gate1587(.a(s_149), .O(gate282inter4));
  nand2 gate1588(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1589(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1590(.a(G782), .O(gate282inter7));
  inv1  gate1591(.a(G806), .O(gate282inter8));
  nand2 gate1592(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1593(.a(s_149), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1594(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1595(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1596(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1527(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1528(.a(gate288inter0), .b(s_140), .O(gate288inter1));
  and2  gate1529(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1530(.a(s_140), .O(gate288inter3));
  inv1  gate1531(.a(s_141), .O(gate288inter4));
  nand2 gate1532(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1533(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1534(.a(G791), .O(gate288inter7));
  inv1  gate1535(.a(G815), .O(gate288inter8));
  nand2 gate1536(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1537(.a(s_141), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1538(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1539(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1540(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1387(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1388(.a(gate293inter0), .b(s_120), .O(gate293inter1));
  and2  gate1389(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1390(.a(s_120), .O(gate293inter3));
  inv1  gate1391(.a(s_121), .O(gate293inter4));
  nand2 gate1392(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1393(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1394(.a(G828), .O(gate293inter7));
  inv1  gate1395(.a(G829), .O(gate293inter8));
  nand2 gate1396(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1397(.a(s_121), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1398(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1399(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1400(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate743(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate744(.a(gate294inter0), .b(s_28), .O(gate294inter1));
  and2  gate745(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate746(.a(s_28), .O(gate294inter3));
  inv1  gate747(.a(s_29), .O(gate294inter4));
  nand2 gate748(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate749(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate750(.a(G832), .O(gate294inter7));
  inv1  gate751(.a(G833), .O(gate294inter8));
  nand2 gate752(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate753(.a(s_29), .b(gate294inter3), .O(gate294inter10));
  nor2  gate754(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate755(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate756(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1625(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1626(.a(gate387inter0), .b(s_154), .O(gate387inter1));
  and2  gate1627(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1628(.a(s_154), .O(gate387inter3));
  inv1  gate1629(.a(s_155), .O(gate387inter4));
  nand2 gate1630(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1631(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1632(.a(G1), .O(gate387inter7));
  inv1  gate1633(.a(G1036), .O(gate387inter8));
  nand2 gate1634(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1635(.a(s_155), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1636(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1637(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1638(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1429(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1430(.a(gate388inter0), .b(s_126), .O(gate388inter1));
  and2  gate1431(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1432(.a(s_126), .O(gate388inter3));
  inv1  gate1433(.a(s_127), .O(gate388inter4));
  nand2 gate1434(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1435(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1436(.a(G2), .O(gate388inter7));
  inv1  gate1437(.a(G1039), .O(gate388inter8));
  nand2 gate1438(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1439(.a(s_127), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1440(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1441(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1442(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1247(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1248(.a(gate389inter0), .b(s_100), .O(gate389inter1));
  and2  gate1249(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1250(.a(s_100), .O(gate389inter3));
  inv1  gate1251(.a(s_101), .O(gate389inter4));
  nand2 gate1252(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1253(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1254(.a(G3), .O(gate389inter7));
  inv1  gate1255(.a(G1042), .O(gate389inter8));
  nand2 gate1256(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1257(.a(s_101), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1258(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1259(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1260(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1737(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1738(.a(gate400inter0), .b(s_170), .O(gate400inter1));
  and2  gate1739(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1740(.a(s_170), .O(gate400inter3));
  inv1  gate1741(.a(s_171), .O(gate400inter4));
  nand2 gate1742(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1743(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1744(.a(G14), .O(gate400inter7));
  inv1  gate1745(.a(G1075), .O(gate400inter8));
  nand2 gate1746(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1747(.a(s_171), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1748(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1749(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1750(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate701(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate702(.a(gate408inter0), .b(s_22), .O(gate408inter1));
  and2  gate703(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate704(.a(s_22), .O(gate408inter3));
  inv1  gate705(.a(s_23), .O(gate408inter4));
  nand2 gate706(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate707(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate708(.a(G22), .O(gate408inter7));
  inv1  gate709(.a(G1099), .O(gate408inter8));
  nand2 gate710(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate711(.a(s_23), .b(gate408inter3), .O(gate408inter10));
  nor2  gate712(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate713(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate714(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1653(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1654(.a(gate418inter0), .b(s_158), .O(gate418inter1));
  and2  gate1655(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1656(.a(s_158), .O(gate418inter3));
  inv1  gate1657(.a(s_159), .O(gate418inter4));
  nand2 gate1658(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1659(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1660(.a(G32), .O(gate418inter7));
  inv1  gate1661(.a(G1129), .O(gate418inter8));
  nand2 gate1662(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1663(.a(s_159), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1664(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1665(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1666(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1177(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1178(.a(gate420inter0), .b(s_90), .O(gate420inter1));
  and2  gate1179(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1180(.a(s_90), .O(gate420inter3));
  inv1  gate1181(.a(s_91), .O(gate420inter4));
  nand2 gate1182(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1183(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1184(.a(G1036), .O(gate420inter7));
  inv1  gate1185(.a(G1132), .O(gate420inter8));
  nand2 gate1186(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1187(.a(s_91), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1188(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1189(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1190(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate869(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate870(.a(gate422inter0), .b(s_46), .O(gate422inter1));
  and2  gate871(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate872(.a(s_46), .O(gate422inter3));
  inv1  gate873(.a(s_47), .O(gate422inter4));
  nand2 gate874(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate875(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate876(.a(G1039), .O(gate422inter7));
  inv1  gate877(.a(G1135), .O(gate422inter8));
  nand2 gate878(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate879(.a(s_47), .b(gate422inter3), .O(gate422inter10));
  nor2  gate880(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate881(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate882(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1485(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1486(.a(gate435inter0), .b(s_134), .O(gate435inter1));
  and2  gate1487(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1488(.a(s_134), .O(gate435inter3));
  inv1  gate1489(.a(s_135), .O(gate435inter4));
  nand2 gate1490(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1491(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1492(.a(G9), .O(gate435inter7));
  inv1  gate1493(.a(G1156), .O(gate435inter8));
  nand2 gate1494(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1495(.a(s_135), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1496(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1497(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1498(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1303(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1304(.a(gate436inter0), .b(s_108), .O(gate436inter1));
  and2  gate1305(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1306(.a(s_108), .O(gate436inter3));
  inv1  gate1307(.a(s_109), .O(gate436inter4));
  nand2 gate1308(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1309(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1310(.a(G1060), .O(gate436inter7));
  inv1  gate1311(.a(G1156), .O(gate436inter8));
  nand2 gate1312(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1313(.a(s_109), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1314(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1315(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1316(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate827(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate828(.a(gate438inter0), .b(s_40), .O(gate438inter1));
  and2  gate829(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate830(.a(s_40), .O(gate438inter3));
  inv1  gate831(.a(s_41), .O(gate438inter4));
  nand2 gate832(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate833(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate834(.a(G1063), .O(gate438inter7));
  inv1  gate835(.a(G1159), .O(gate438inter8));
  nand2 gate836(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate837(.a(s_41), .b(gate438inter3), .O(gate438inter10));
  nor2  gate838(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate839(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate840(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1065(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1066(.a(gate443inter0), .b(s_74), .O(gate443inter1));
  and2  gate1067(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1068(.a(s_74), .O(gate443inter3));
  inv1  gate1069(.a(s_75), .O(gate443inter4));
  nand2 gate1070(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1071(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1072(.a(G13), .O(gate443inter7));
  inv1  gate1073(.a(G1168), .O(gate443inter8));
  nand2 gate1074(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1075(.a(s_75), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1076(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1077(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1078(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate883(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate884(.a(gate460inter0), .b(s_48), .O(gate460inter1));
  and2  gate885(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate886(.a(s_48), .O(gate460inter3));
  inv1  gate887(.a(s_49), .O(gate460inter4));
  nand2 gate888(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate889(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate890(.a(G1096), .O(gate460inter7));
  inv1  gate891(.a(G1192), .O(gate460inter8));
  nand2 gate892(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate893(.a(s_49), .b(gate460inter3), .O(gate460inter10));
  nor2  gate894(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate895(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate896(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1499(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1500(.a(gate462inter0), .b(s_136), .O(gate462inter1));
  and2  gate1501(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1502(.a(s_136), .O(gate462inter3));
  inv1  gate1503(.a(s_137), .O(gate462inter4));
  nand2 gate1504(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1505(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1506(.a(G1099), .O(gate462inter7));
  inv1  gate1507(.a(G1195), .O(gate462inter8));
  nand2 gate1508(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1509(.a(s_137), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1510(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1511(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1512(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate757(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate758(.a(gate463inter0), .b(s_30), .O(gate463inter1));
  and2  gate759(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate760(.a(s_30), .O(gate463inter3));
  inv1  gate761(.a(s_31), .O(gate463inter4));
  nand2 gate762(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate763(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate764(.a(G23), .O(gate463inter7));
  inv1  gate765(.a(G1198), .O(gate463inter8));
  nand2 gate766(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate767(.a(s_31), .b(gate463inter3), .O(gate463inter10));
  nor2  gate768(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate769(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate770(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1331(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1332(.a(gate464inter0), .b(s_112), .O(gate464inter1));
  and2  gate1333(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1334(.a(s_112), .O(gate464inter3));
  inv1  gate1335(.a(s_113), .O(gate464inter4));
  nand2 gate1336(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1337(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1338(.a(G1102), .O(gate464inter7));
  inv1  gate1339(.a(G1198), .O(gate464inter8));
  nand2 gate1340(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1341(.a(s_113), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1342(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1343(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1344(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1793(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1794(.a(gate466inter0), .b(s_178), .O(gate466inter1));
  and2  gate1795(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1796(.a(s_178), .O(gate466inter3));
  inv1  gate1797(.a(s_179), .O(gate466inter4));
  nand2 gate1798(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1799(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1800(.a(G1105), .O(gate466inter7));
  inv1  gate1801(.a(G1201), .O(gate466inter8));
  nand2 gate1802(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1803(.a(s_179), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1804(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1805(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1806(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1373(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1374(.a(gate467inter0), .b(s_118), .O(gate467inter1));
  and2  gate1375(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1376(.a(s_118), .O(gate467inter3));
  inv1  gate1377(.a(s_119), .O(gate467inter4));
  nand2 gate1378(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1379(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1380(.a(G25), .O(gate467inter7));
  inv1  gate1381(.a(G1204), .O(gate467inter8));
  nand2 gate1382(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1383(.a(s_119), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1384(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1385(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1386(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate547(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate548(.a(gate468inter0), .b(s_0), .O(gate468inter1));
  and2  gate549(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate550(.a(s_0), .O(gate468inter3));
  inv1  gate551(.a(s_1), .O(gate468inter4));
  nand2 gate552(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate553(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate554(.a(G1108), .O(gate468inter7));
  inv1  gate555(.a(G1204), .O(gate468inter8));
  nand2 gate556(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate557(.a(s_1), .b(gate468inter3), .O(gate468inter10));
  nor2  gate558(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate559(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate560(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate939(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate940(.a(gate471inter0), .b(s_56), .O(gate471inter1));
  and2  gate941(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate942(.a(s_56), .O(gate471inter3));
  inv1  gate943(.a(s_57), .O(gate471inter4));
  nand2 gate944(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate945(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate946(.a(G27), .O(gate471inter7));
  inv1  gate947(.a(G1210), .O(gate471inter8));
  nand2 gate948(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate949(.a(s_57), .b(gate471inter3), .O(gate471inter10));
  nor2  gate950(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate951(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate952(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate631(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate632(.a(gate473inter0), .b(s_12), .O(gate473inter1));
  and2  gate633(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate634(.a(s_12), .O(gate473inter3));
  inv1  gate635(.a(s_13), .O(gate473inter4));
  nand2 gate636(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate637(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate638(.a(G28), .O(gate473inter7));
  inv1  gate639(.a(G1213), .O(gate473inter8));
  nand2 gate640(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate641(.a(s_13), .b(gate473inter3), .O(gate473inter10));
  nor2  gate642(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate643(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate644(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate687(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate688(.a(gate486inter0), .b(s_20), .O(gate486inter1));
  and2  gate689(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate690(.a(s_20), .O(gate486inter3));
  inv1  gate691(.a(s_21), .O(gate486inter4));
  nand2 gate692(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate693(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate694(.a(G1234), .O(gate486inter7));
  inv1  gate695(.a(G1235), .O(gate486inter8));
  nand2 gate696(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate697(.a(s_21), .b(gate486inter3), .O(gate486inter10));
  nor2  gate698(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate699(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate700(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1233(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1234(.a(gate505inter0), .b(s_98), .O(gate505inter1));
  and2  gate1235(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1236(.a(s_98), .O(gate505inter3));
  inv1  gate1237(.a(s_99), .O(gate505inter4));
  nand2 gate1238(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1239(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1240(.a(G1272), .O(gate505inter7));
  inv1  gate1241(.a(G1273), .O(gate505inter8));
  nand2 gate1242(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1243(.a(s_99), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1244(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1245(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1246(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1471(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1472(.a(gate506inter0), .b(s_132), .O(gate506inter1));
  and2  gate1473(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1474(.a(s_132), .O(gate506inter3));
  inv1  gate1475(.a(s_133), .O(gate506inter4));
  nand2 gate1476(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1477(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1478(.a(G1274), .O(gate506inter7));
  inv1  gate1479(.a(G1275), .O(gate506inter8));
  nand2 gate1480(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1481(.a(s_133), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1482(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1483(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1484(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate911(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate912(.a(gate512inter0), .b(s_52), .O(gate512inter1));
  and2  gate913(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate914(.a(s_52), .O(gate512inter3));
  inv1  gate915(.a(s_53), .O(gate512inter4));
  nand2 gate916(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate917(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate918(.a(G1286), .O(gate512inter7));
  inv1  gate919(.a(G1287), .O(gate512inter8));
  nand2 gate920(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate921(.a(s_53), .b(gate512inter3), .O(gate512inter10));
  nor2  gate922(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate923(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate924(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule