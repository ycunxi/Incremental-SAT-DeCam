module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate858inter0, gate858inter1, gate858inter2, gate858inter3, gate858inter4, gate858inter5, gate858inter6, gate858inter7, gate858inter8, gate858inter9, gate858inter10, gate858inter11, gate858inter12, gate808inter0, gate808inter1, gate808inter2, gate808inter3, gate808inter4, gate808inter5, gate808inter6, gate808inter7, gate808inter8, gate808inter9, gate808inter10, gate808inter11, gate808inter12, gate340inter0, gate340inter1, gate340inter2, gate340inter3, gate340inter4, gate340inter5, gate340inter6, gate340inter7, gate340inter8, gate340inter9, gate340inter10, gate340inter11, gate340inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate380inter0, gate380inter1, gate380inter2, gate380inter3, gate380inter4, gate380inter5, gate380inter6, gate380inter7, gate380inter8, gate380inter9, gate380inter10, gate380inter11, gate380inter12, gate765inter0, gate765inter1, gate765inter2, gate765inter3, gate765inter4, gate765inter5, gate765inter6, gate765inter7, gate765inter8, gate765inter9, gate765inter10, gate765inter11, gate765inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate527inter0, gate527inter1, gate527inter2, gate527inter3, gate527inter4, gate527inter5, gate527inter6, gate527inter7, gate527inter8, gate527inter9, gate527inter10, gate527inter11, gate527inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate351inter0, gate351inter1, gate351inter2, gate351inter3, gate351inter4, gate351inter5, gate351inter6, gate351inter7, gate351inter8, gate351inter9, gate351inter10, gate351inter11, gate351inter12, gate818inter0, gate818inter1, gate818inter2, gate818inter3, gate818inter4, gate818inter5, gate818inter6, gate818inter7, gate818inter8, gate818inter9, gate818inter10, gate818inter11, gate818inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate329inter0, gate329inter1, gate329inter2, gate329inter3, gate329inter4, gate329inter5, gate329inter6, gate329inter7, gate329inter8, gate329inter9, gate329inter10, gate329inter11, gate329inter12, gate517inter0, gate517inter1, gate517inter2, gate517inter3, gate517inter4, gate517inter5, gate517inter6, gate517inter7, gate517inter8, gate517inter9, gate517inter10, gate517inter11, gate517inter12, gate600inter0, gate600inter1, gate600inter2, gate600inter3, gate600inter4, gate600inter5, gate600inter6, gate600inter7, gate600inter8, gate600inter9, gate600inter10, gate600inter11, gate600inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate802inter0, gate802inter1, gate802inter2, gate802inter3, gate802inter4, gate802inter5, gate802inter6, gate802inter7, gate802inter8, gate802inter9, gate802inter10, gate802inter11, gate802inter12, gate794inter0, gate794inter1, gate794inter2, gate794inter3, gate794inter4, gate794inter5, gate794inter6, gate794inter7, gate794inter8, gate794inter9, gate794inter10, gate794inter11, gate794inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate616inter0, gate616inter1, gate616inter2, gate616inter3, gate616inter4, gate616inter5, gate616inter6, gate616inter7, gate616inter8, gate616inter9, gate616inter10, gate616inter11, gate616inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate649inter0, gate649inter1, gate649inter2, gate649inter3, gate649inter4, gate649inter5, gate649inter6, gate649inter7, gate649inter8, gate649inter9, gate649inter10, gate649inter11, gate649inter12, gate539inter0, gate539inter1, gate539inter2, gate539inter3, gate539inter4, gate539inter5, gate539inter6, gate539inter7, gate539inter8, gate539inter9, gate539inter10, gate539inter11, gate539inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate526inter0, gate526inter1, gate526inter2, gate526inter3, gate526inter4, gate526inter5, gate526inter6, gate526inter7, gate526inter8, gate526inter9, gate526inter10, gate526inter11, gate526inter12, gate582inter0, gate582inter1, gate582inter2, gate582inter3, gate582inter4, gate582inter5, gate582inter6, gate582inter7, gate582inter8, gate582inter9, gate582inter10, gate582inter11, gate582inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate809inter0, gate809inter1, gate809inter2, gate809inter3, gate809inter4, gate809inter5, gate809inter6, gate809inter7, gate809inter8, gate809inter9, gate809inter10, gate809inter11, gate809inter12, gate518inter0, gate518inter1, gate518inter2, gate518inter3, gate518inter4, gate518inter5, gate518inter6, gate518inter7, gate518inter8, gate518inter9, gate518inter10, gate518inter11, gate518inter12, gate530inter0, gate530inter1, gate530inter2, gate530inter3, gate530inter4, gate530inter5, gate530inter6, gate530inter7, gate530inter8, gate530inter9, gate530inter10, gate530inter11, gate530inter12, gate543inter0, gate543inter1, gate543inter2, gate543inter3, gate543inter4, gate543inter5, gate543inter6, gate543inter7, gate543inter8, gate543inter9, gate543inter10, gate543inter11, gate543inter12, gate838inter0, gate838inter1, gate838inter2, gate838inter3, gate838inter4, gate838inter5, gate838inter6, gate838inter7, gate838inter8, gate838inter9, gate838inter10, gate838inter11, gate838inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate786inter0, gate786inter1, gate786inter2, gate786inter3, gate786inter4, gate786inter5, gate786inter6, gate786inter7, gate786inter8, gate786inter9, gate786inter10, gate786inter11, gate786inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate861inter0, gate861inter1, gate861inter2, gate861inter3, gate861inter4, gate861inter5, gate861inter6, gate861inter7, gate861inter8, gate861inter9, gate861inter10, gate861inter11, gate861inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate318inter0, gate318inter1, gate318inter2, gate318inter3, gate318inter4, gate318inter5, gate318inter6, gate318inter7, gate318inter8, gate318inter9, gate318inter10, gate318inter11, gate318inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate752inter0, gate752inter1, gate752inter2, gate752inter3, gate752inter4, gate752inter5, gate752inter6, gate752inter7, gate752inter8, gate752inter9, gate752inter10, gate752inter11, gate752inter12, gate524inter0, gate524inter1, gate524inter2, gate524inter3, gate524inter4, gate524inter5, gate524inter6, gate524inter7, gate524inter8, gate524inter9, gate524inter10, gate524inter11, gate524inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate345inter0, gate345inter1, gate345inter2, gate345inter3, gate345inter4, gate345inter5, gate345inter6, gate345inter7, gate345inter8, gate345inter9, gate345inter10, gate345inter11, gate345inter12, gate637inter0, gate637inter1, gate637inter2, gate637inter3, gate637inter4, gate637inter5, gate637inter6, gate637inter7, gate637inter8, gate637inter9, gate637inter10, gate637inter11, gate637inter12, gate681inter0, gate681inter1, gate681inter2, gate681inter3, gate681inter4, gate681inter5, gate681inter6, gate681inter7, gate681inter8, gate681inter9, gate681inter10, gate681inter11, gate681inter12, gate608inter0, gate608inter1, gate608inter2, gate608inter3, gate608inter4, gate608inter5, gate608inter6, gate608inter7, gate608inter8, gate608inter9, gate608inter10, gate608inter11, gate608inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate363inter0, gate363inter1, gate363inter2, gate363inter3, gate363inter4, gate363inter5, gate363inter6, gate363inter7, gate363inter8, gate363inter9, gate363inter10, gate363inter11, gate363inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate828inter0, gate828inter1, gate828inter2, gate828inter3, gate828inter4, gate828inter5, gate828inter6, gate828inter7, gate828inter8, gate828inter9, gate828inter10, gate828inter11, gate828inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate779inter0, gate779inter1, gate779inter2, gate779inter3, gate779inter4, gate779inter5, gate779inter6, gate779inter7, gate779inter8, gate779inter9, gate779inter10, gate779inter11, gate779inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate663inter0, gate663inter1, gate663inter2, gate663inter3, gate663inter4, gate663inter5, gate663inter6, gate663inter7, gate663inter8, gate663inter9, gate663inter10, gate663inter11, gate663inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate624inter0, gate624inter1, gate624inter2, gate624inter3, gate624inter4, gate624inter5, gate624inter6, gate624inter7, gate624inter8, gate624inter9, gate624inter10, gate624inter11, gate624inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate534inter0, gate534inter1, gate534inter2, gate534inter3, gate534inter4, gate534inter5, gate534inter6, gate534inter7, gate534inter8, gate534inter9, gate534inter10, gate534inter11, gate534inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate771inter0, gate771inter1, gate771inter2, gate771inter3, gate771inter4, gate771inter5, gate771inter6, gate771inter7, gate771inter8, gate771inter9, gate771inter10, gate771inter11, gate771inter12;



inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate1749(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate1750(.a(gate17inter0), .b(s_124), .O(gate17inter1));
  and2  gate1751(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate1752(.a(s_124), .O(gate17inter3));
  inv1  gate1753(.a(s_125), .O(gate17inter4));
  nand2 gate1754(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1755(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1756(.a(N63), .O(gate17inter7));
  inv1  gate1757(.a(N88), .O(gate17inter8));
  nand2 gate1758(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1759(.a(s_125), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1760(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1761(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1762(.a(gate17inter12), .b(gate17inter1), .O(N251));
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );

  xor2  gate965(.a(N331), .b(N306), .O(gate75inter0));
  nand2 gate966(.a(gate75inter0), .b(s_12), .O(gate75inter1));
  and2  gate967(.a(N331), .b(N306), .O(gate75inter2));
  inv1  gate968(.a(s_12), .O(gate75inter3));
  inv1  gate969(.a(s_13), .O(gate75inter4));
  nand2 gate970(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate971(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate972(.a(N306), .O(gate75inter7));
  inv1  gate973(.a(N331), .O(gate75inter8));
  nand2 gate974(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate975(.a(s_13), .b(gate75inter3), .O(gate75inter10));
  nor2  gate976(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate977(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate978(.a(gate75inter12), .b(gate75inter1), .O(N550));
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );

  xor2  gate1259(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate1260(.a(gate79inter0), .b(s_54), .O(gate79inter1));
  and2  gate1261(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate1262(.a(s_54), .O(gate79inter3));
  inv1  gate1263(.a(s_55), .O(gate79inter4));
  nand2 gate1264(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1265(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1266(.a(N306), .O(gate79inter7));
  inv1  gate1267(.a(N331), .O(gate79inter8));
  nand2 gate1268(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1269(.a(s_55), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1270(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1271(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1272(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );

  xor2  gate2267(.a(N280), .b(N326), .O(gate97inter0));
  nand2 gate2268(.a(gate97inter0), .b(s_198), .O(gate97inter1));
  and2  gate2269(.a(N280), .b(N326), .O(gate97inter2));
  inv1  gate2270(.a(s_198), .O(gate97inter3));
  inv1  gate2271(.a(s_199), .O(gate97inter4));
  nand2 gate2272(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2273(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2274(.a(N326), .O(gate97inter7));
  inv1  gate2275(.a(N280), .O(gate97inter8));
  nand2 gate2276(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2277(.a(s_199), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2278(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2279(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2280(.a(gate97inter12), .b(gate97inter1), .O(N602));

  xor2  gate1413(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate1414(.a(gate98inter0), .b(s_76), .O(gate98inter1));
  and2  gate1415(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate1416(.a(s_76), .O(gate98inter3));
  inv1  gate1417(.a(s_77), .O(gate98inter4));
  nand2 gate1418(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1419(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1420(.a(N260), .O(gate98inter7));
  inv1  gate1421(.a(N72), .O(gate98inter8));
  nand2 gate1422(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1423(.a(s_77), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1424(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1425(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1426(.a(gate98inter12), .b(gate98inter1), .O(N603));
nand2 gate99( .a(N260), .b(N300), .O(N608) );

  xor2  gate1385(.a(N300), .b(N256), .O(gate100inter0));
  nand2 gate1386(.a(gate100inter0), .b(s_72), .O(gate100inter1));
  and2  gate1387(.a(N300), .b(N256), .O(gate100inter2));
  inv1  gate1388(.a(s_72), .O(gate100inter3));
  inv1  gate1389(.a(s_73), .O(gate100inter4));
  nand2 gate1390(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1391(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1392(.a(N256), .O(gate100inter7));
  inv1  gate1393(.a(N300), .O(gate100inter8));
  nand2 gate1394(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1395(.a(s_73), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1396(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1397(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1398(.a(gate100inter12), .b(gate100inter1), .O(N612));
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );

  xor2  gate1791(.a(N989), .b(N718), .O(gate240inter0));
  nand2 gate1792(.a(gate240inter0), .b(s_130), .O(gate240inter1));
  and2  gate1793(.a(N989), .b(N718), .O(gate240inter2));
  inv1  gate1794(.a(s_130), .O(gate240inter3));
  inv1  gate1795(.a(s_131), .O(gate240inter4));
  nand2 gate1796(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1797(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1798(.a(N718), .O(gate240inter7));
  inv1  gate1799(.a(N989), .O(gate240inter8));
  nand2 gate1800(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1801(.a(s_131), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1802(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1803(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1804(.a(gate240inter12), .b(gate240inter1), .O(N1120));
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );

  xor2  gate1637(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate1638(.a(gate244inter0), .b(s_108), .O(gate244inter1));
  and2  gate1639(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate1640(.a(s_108), .O(gate244inter3));
  inv1  gate1641(.a(s_109), .O(gate244inter4));
  nand2 gate1642(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1643(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1644(.a(N736), .O(gate244inter7));
  inv1  gate1645(.a(N1003), .O(gate244inter8));
  nand2 gate1646(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1647(.a(s_109), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1648(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1649(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1650(.a(gate244inter12), .b(gate244inter1), .O(N1129));
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate1063(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate1064(.a(gate268inter0), .b(s_26), .O(gate268inter1));
  and2  gate1065(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate1066(.a(s_26), .O(gate268inter3));
  inv1  gate1067(.a(s_27), .O(gate268inter4));
  nand2 gate1068(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1069(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1070(.a(N921), .O(gate268inter7));
  inv1  gate1071(.a(N923), .O(gate268inter8));
  nand2 gate1072(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1073(.a(s_27), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1074(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1075(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1076(.a(gate268inter12), .b(gate268inter1), .O(N1171));

  xor2  gate1105(.a(N923), .b(N922), .O(gate269inter0));
  nand2 gate1106(.a(gate269inter0), .b(s_32), .O(gate269inter1));
  and2  gate1107(.a(N923), .b(N922), .O(gate269inter2));
  inv1  gate1108(.a(s_32), .O(gate269inter3));
  inv1  gate1109(.a(s_33), .O(gate269inter4));
  nand2 gate1110(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1111(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1112(.a(N922), .O(gate269inter7));
  inv1  gate1113(.a(N923), .O(gate269inter8));
  nand2 gate1114(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1115(.a(s_33), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1116(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1117(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1118(.a(gate269inter12), .b(gate269inter1), .O(N1188));
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate1133(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate1134(.a(gate273inter0), .b(s_36), .O(gate273inter1));
  and2  gate1135(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate1136(.a(s_36), .O(gate273inter3));
  inv1  gate1137(.a(s_37), .O(gate273inter4));
  nand2 gate1138(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1139(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1140(.a(N1013), .O(gate273inter7));
  inv1  gate1141(.a(N942), .O(gate273inter8));
  nand2 gate1142(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1143(.a(s_37), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1144(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1145(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1146(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate1077(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate1078(.a(gate275inter0), .b(s_28), .O(gate275inter1));
  and2  gate1079(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate1080(.a(s_28), .O(gate275inter3));
  inv1  gate1081(.a(s_29), .O(gate275inter4));
  nand2 gate1082(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1083(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1084(.a(N1016), .O(gate275inter7));
  inv1  gate1085(.a(N946), .O(gate275inter8));
  nand2 gate1086(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1087(.a(s_29), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1088(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1089(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1090(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate881(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate882(.a(gate277inter0), .b(s_0), .O(gate277inter1));
  and2  gate883(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate884(.a(s_0), .O(gate277inter3));
  inv1  gate885(.a(s_1), .O(gate277inter4));
  nand2 gate886(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate887(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate888(.a(N1019), .O(gate277inter7));
  inv1  gate889(.a(N950), .O(gate277inter8));
  nand2 gate890(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate891(.a(s_1), .b(gate277inter3), .O(gate277inter10));
  nor2  gate892(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate893(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate894(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );

  xor2  gate1595(.a(N954), .b(N1022), .O(gate279inter0));
  nand2 gate1596(.a(gate279inter0), .b(s_102), .O(gate279inter1));
  and2  gate1597(.a(N954), .b(N1022), .O(gate279inter2));
  inv1  gate1598(.a(s_102), .O(gate279inter3));
  inv1  gate1599(.a(s_103), .O(gate279inter4));
  nand2 gate1600(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1601(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1602(.a(N1022), .O(gate279inter7));
  inv1  gate1603(.a(N954), .O(gate279inter8));
  nand2 gate1604(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1605(.a(s_103), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1606(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1607(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1608(.a(gate279inter12), .b(gate279inter1), .O(N1214));
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );

  xor2  gate1721(.a(N976), .b(N1040), .O(gate291inter0));
  nand2 gate1722(.a(gate291inter0), .b(s_120), .O(gate291inter1));
  and2  gate1723(.a(N976), .b(N1040), .O(gate291inter2));
  inv1  gate1724(.a(s_120), .O(gate291inter3));
  inv1  gate1725(.a(s_121), .O(gate291inter4));
  nand2 gate1726(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1727(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1728(.a(N1040), .O(gate291inter7));
  inv1  gate1729(.a(N976), .O(gate291inter8));
  nand2 gate1730(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1731(.a(s_121), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1732(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1733(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1734(.a(gate291inter12), .b(gate291inter1), .O(N1226));
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );

  xor2  gate1623(.a(N984), .b(N981), .O(gate296inter0));
  nand2 gate1624(.a(gate296inter0), .b(s_106), .O(gate296inter1));
  and2  gate1625(.a(N984), .b(N981), .O(gate296inter2));
  inv1  gate1626(.a(s_106), .O(gate296inter3));
  inv1  gate1627(.a(s_107), .O(gate296inter4));
  nand2 gate1628(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1629(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1630(.a(N981), .O(gate296inter7));
  inv1  gate1631(.a(N984), .O(gate296inter8));
  nand2 gate1632(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1633(.a(s_107), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1634(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1635(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1636(.a(gate296inter12), .b(gate296inter1), .O(N1231));

  xor2  gate1315(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate1316(.a(gate297inter0), .b(s_62), .O(gate297inter1));
  and2  gate1317(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate1318(.a(s_62), .O(gate297inter3));
  inv1  gate1319(.a(s_63), .O(gate297inter4));
  nand2 gate1320(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate1321(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate1322(.a(N1119), .O(gate297inter7));
  inv1  gate1323(.a(N1120), .O(gate297inter8));
  nand2 gate1324(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate1325(.a(s_63), .b(gate297inter3), .O(gate297inter10));
  nor2  gate1326(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate1327(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate1328(.a(gate297inter12), .b(gate297inter1), .O(N1232));
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );

  xor2  gate1371(.a(N997), .b(N1046), .O(gate300inter0));
  nand2 gate1372(.a(gate300inter0), .b(s_70), .O(gate300inter1));
  and2  gate1373(.a(N997), .b(N1046), .O(gate300inter2));
  inv1  gate1374(.a(s_70), .O(gate300inter3));
  inv1  gate1375(.a(s_71), .O(gate300inter4));
  nand2 gate1376(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate1377(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate1378(.a(N1046), .O(gate300inter7));
  inv1  gate1379(.a(N997), .O(gate300inter8));
  nand2 gate1380(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate1381(.a(s_71), .b(gate300inter3), .O(gate300inter10));
  nor2  gate1382(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate1383(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate1384(.a(gate300inter12), .b(gate300inter1), .O(N1239));
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );

  xor2  gate1091(.a(N1207), .b(N691), .O(gate314inter0));
  nand2 gate1092(.a(gate314inter0), .b(s_30), .O(gate314inter1));
  and2  gate1093(.a(N1207), .b(N691), .O(gate314inter2));
  inv1  gate1094(.a(s_30), .O(gate314inter3));
  inv1  gate1095(.a(s_31), .O(gate314inter4));
  nand2 gate1096(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate1097(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate1098(.a(N691), .O(gate314inter7));
  inv1  gate1099(.a(N1207), .O(gate314inter8));
  nand2 gate1100(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate1101(.a(s_31), .b(gate314inter3), .O(gate314inter10));
  nor2  gate1102(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate1103(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate1104(.a(gate314inter12), .b(gate314inter1), .O(N1310));
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );

  xor2  gate2323(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate2324(.a(gate316inter0), .b(s_206), .O(gate316inter1));
  and2  gate2325(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate2326(.a(s_206), .O(gate316inter3));
  inv1  gate2327(.a(s_207), .O(gate316inter4));
  nand2 gate2328(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate2329(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate2330(.a(N697), .O(gate316inter7));
  inv1  gate2331(.a(N1211), .O(gate316inter8));
  nand2 gate2332(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate2333(.a(s_207), .b(gate316inter3), .O(gate316inter10));
  nor2  gate2334(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate2335(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate2336(.a(gate316inter12), .b(gate316inter1), .O(N1312));
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );

  xor2  gate1819(.a(N1215), .b(N703), .O(gate318inter0));
  nand2 gate1820(.a(gate318inter0), .b(s_134), .O(gate318inter1));
  and2  gate1821(.a(N1215), .b(N703), .O(gate318inter2));
  inv1  gate1822(.a(s_134), .O(gate318inter3));
  inv1  gate1823(.a(s_135), .O(gate318inter4));
  nand2 gate1824(.a(gate318inter4), .b(gate318inter3), .O(gate318inter5));
  nor2  gate1825(.a(gate318inter5), .b(gate318inter2), .O(gate318inter6));
  inv1  gate1826(.a(N703), .O(gate318inter7));
  inv1  gate1827(.a(N1215), .O(gate318inter8));
  nand2 gate1828(.a(gate318inter8), .b(gate318inter7), .O(gate318inter9));
  nand2 gate1829(.a(s_135), .b(gate318inter3), .O(gate318inter10));
  nor2  gate1830(.a(gate318inter10), .b(gate318inter9), .O(gate318inter11));
  nor2  gate1831(.a(gate318inter11), .b(gate318inter6), .O(gate318inter12));
  nand2 gate1832(.a(gate318inter12), .b(gate318inter1), .O(N1314));
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );

  xor2  gate2085(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate2086(.a(gate326inter0), .b(s_172), .O(gate326inter1));
  and2  gate2087(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate2088(.a(s_172), .O(gate326inter3));
  inv1  gate2089(.a(s_173), .O(gate326inter4));
  nand2 gate2090(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate2091(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate2092(.a(N733), .O(gate326inter7));
  inv1  gate2093(.a(N1241), .O(gate326inter8));
  nand2 gate2094(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate2095(.a(s_173), .b(gate326inter3), .O(gate326inter10));
  nor2  gate2096(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate2097(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate2098(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );

  xor2  gate1273(.a(N894), .b(N1249), .O(gate329inter0));
  nand2 gate1274(.a(gate329inter0), .b(s_56), .O(gate329inter1));
  and2  gate1275(.a(N894), .b(N1249), .O(gate329inter2));
  inv1  gate1276(.a(s_56), .O(gate329inter3));
  inv1  gate1277(.a(s_57), .O(gate329inter4));
  nand2 gate1278(.a(gate329inter4), .b(gate329inter3), .O(gate329inter5));
  nor2  gate1279(.a(gate329inter5), .b(gate329inter2), .O(gate329inter6));
  inv1  gate1280(.a(N1249), .O(gate329inter7));
  inv1  gate1281(.a(N894), .O(gate329inter8));
  nand2 gate1282(.a(gate329inter8), .b(gate329inter7), .O(gate329inter9));
  nand2 gate1283(.a(s_57), .b(gate329inter3), .O(gate329inter10));
  nor2  gate1284(.a(gate329inter10), .b(gate329inter9), .O(gate329inter11));
  nor2  gate1285(.a(gate329inter11), .b(gate329inter6), .O(gate329inter12));
  nand2 gate1286(.a(gate329inter12), .b(gate329inter1), .O(N1345));
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );

  xor2  gate923(.a(N1216), .b(N1314), .O(gate340inter0));
  nand2 gate924(.a(gate340inter0), .b(s_6), .O(gate340inter1));
  and2  gate925(.a(N1216), .b(N1314), .O(gate340inter2));
  inv1  gate926(.a(s_6), .O(gate340inter3));
  inv1  gate927(.a(s_7), .O(gate340inter4));
  nand2 gate928(.a(gate340inter4), .b(gate340inter3), .O(gate340inter5));
  nor2  gate929(.a(gate340inter5), .b(gate340inter2), .O(gate340inter6));
  inv1  gate930(.a(N1314), .O(gate340inter7));
  inv1  gate931(.a(N1216), .O(gate340inter8));
  nand2 gate932(.a(gate340inter8), .b(gate340inter7), .O(gate340inter9));
  nand2 gate933(.a(s_7), .b(gate340inter3), .O(gate340inter10));
  nor2  gate934(.a(gate340inter10), .b(gate340inter9), .O(gate340inter11));
  nor2  gate935(.a(gate340inter11), .b(gate340inter6), .O(gate340inter12));
  nand2 gate936(.a(gate340inter12), .b(gate340inter1), .O(N1367));
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );

  xor2  gate2057(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate2058(.a(gate342inter0), .b(s_168), .O(gate342inter1));
  and2  gate2059(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate2060(.a(s_168), .O(gate342inter3));
  inv1  gate2061(.a(s_169), .O(gate342inter4));
  nand2 gate2062(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate2063(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate2064(.a(N1316), .O(gate342inter7));
  inv1  gate2065(.a(N1224), .O(gate342inter8));
  nand2 gate2066(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate2067(.a(s_169), .b(gate342inter3), .O(gate342inter10));
  nor2  gate2068(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate2069(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate2070(.a(gate342inter12), .b(gate342inter1), .O(N1373));
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );

  xor2  gate1049(.a(N1229), .b(N1318), .O(gate344inter0));
  nand2 gate1050(.a(gate344inter0), .b(s_24), .O(gate344inter1));
  and2  gate1051(.a(N1229), .b(N1318), .O(gate344inter2));
  inv1  gate1052(.a(s_24), .O(gate344inter3));
  inv1  gate1053(.a(s_25), .O(gate344inter4));
  nand2 gate1054(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate1055(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate1056(.a(N1318), .O(gate344inter7));
  inv1  gate1057(.a(N1229), .O(gate344inter8));
  nand2 gate1058(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate1059(.a(s_25), .b(gate344inter3), .O(gate344inter10));
  nor2  gate1060(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate1061(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate1062(.a(gate344inter12), .b(gate344inter1), .O(N1379));

  xor2  gate1959(.a(N1231), .b(N1322), .O(gate345inter0));
  nand2 gate1960(.a(gate345inter0), .b(s_154), .O(gate345inter1));
  and2  gate1961(.a(N1231), .b(N1322), .O(gate345inter2));
  inv1  gate1962(.a(s_154), .O(gate345inter3));
  inv1  gate1963(.a(s_155), .O(gate345inter4));
  nand2 gate1964(.a(gate345inter4), .b(gate345inter3), .O(gate345inter5));
  nor2  gate1965(.a(gate345inter5), .b(gate345inter2), .O(gate345inter6));
  inv1  gate1966(.a(N1322), .O(gate345inter7));
  inv1  gate1967(.a(N1231), .O(gate345inter8));
  nand2 gate1968(.a(gate345inter8), .b(gate345inter7), .O(gate345inter9));
  nand2 gate1969(.a(s_155), .b(gate345inter3), .O(gate345inter10));
  nor2  gate1970(.a(gate345inter10), .b(gate345inter9), .O(gate345inter11));
  nor2  gate1971(.a(gate345inter11), .b(gate345inter6), .O(gate345inter12));
  nand2 gate1972(.a(gate345inter12), .b(gate345inter1), .O(N1383));
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );

  xor2  gate1231(.a(N1242), .b(N1328), .O(gate351inter0));
  nand2 gate1232(.a(gate351inter0), .b(s_50), .O(gate351inter1));
  and2  gate1233(.a(N1242), .b(N1328), .O(gate351inter2));
  inv1  gate1234(.a(s_50), .O(gate351inter3));
  inv1  gate1235(.a(s_51), .O(gate351inter4));
  nand2 gate1236(.a(gate351inter4), .b(gate351inter3), .O(gate351inter5));
  nor2  gate1237(.a(gate351inter5), .b(gate351inter2), .O(gate351inter6));
  inv1  gate1238(.a(N1328), .O(gate351inter7));
  inv1  gate1239(.a(N1242), .O(gate351inter8));
  nand2 gate1240(.a(gate351inter8), .b(gate351inter7), .O(gate351inter9));
  nand2 gate1241(.a(s_51), .b(gate351inter3), .O(gate351inter10));
  nor2  gate1242(.a(gate351inter10), .b(gate351inter9), .O(gate351inter11));
  nor2  gate1243(.a(gate351inter11), .b(gate351inter6), .O(gate351inter12));
  nand2 gate1244(.a(gate351inter12), .b(gate351inter1), .O(N1393));
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );

  xor2  gate2099(.a(N1396), .b(N640), .O(gate363inter0));
  nand2 gate2100(.a(gate363inter0), .b(s_174), .O(gate363inter1));
  and2  gate2101(.a(N1396), .b(N640), .O(gate363inter2));
  inv1  gate2102(.a(s_174), .O(gate363inter3));
  inv1  gate2103(.a(s_175), .O(gate363inter4));
  nand2 gate2104(.a(gate363inter4), .b(gate363inter3), .O(gate363inter5));
  nor2  gate2105(.a(gate363inter5), .b(gate363inter2), .O(gate363inter6));
  inv1  gate2106(.a(N640), .O(gate363inter7));
  inv1  gate2107(.a(N1396), .O(gate363inter8));
  nand2 gate2108(.a(gate363inter8), .b(gate363inter7), .O(gate363inter9));
  nand2 gate2109(.a(s_175), .b(gate363inter3), .O(gate363inter10));
  nor2  gate2110(.a(gate363inter10), .b(gate363inter9), .O(gate363inter11));
  nor2  gate2111(.a(gate363inter11), .b(gate363inter6), .O(gate363inter12));
  nand2 gate2112(.a(gate363inter12), .b(gate363inter1), .O(N1438));
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );

  xor2  gate979(.a(N1157), .b(N1379), .O(gate380inter0));
  nand2 gate980(.a(gate380inter0), .b(s_14), .O(gate380inter1));
  and2  gate981(.a(N1157), .b(N1379), .O(gate380inter2));
  inv1  gate982(.a(s_14), .O(gate380inter3));
  inv1  gate983(.a(s_15), .O(gate380inter4));
  nand2 gate984(.a(gate380inter4), .b(gate380inter3), .O(gate380inter5));
  nor2  gate985(.a(gate380inter5), .b(gate380inter2), .O(gate380inter6));
  inv1  gate986(.a(N1379), .O(gate380inter7));
  inv1  gate987(.a(N1157), .O(gate380inter8));
  nand2 gate988(.a(gate380inter8), .b(gate380inter7), .O(gate380inter9));
  nand2 gate989(.a(s_15), .b(gate380inter3), .O(gate380inter10));
  nor2  gate990(.a(gate380inter10), .b(gate380inter9), .O(gate380inter11));
  nor2  gate991(.a(gate380inter11), .b(gate380inter6), .O(gate380inter12));
  nand2 gate992(.a(gate380inter12), .b(gate380inter1), .O(N1459));
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate2295(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate2296(.a(gate383inter0), .b(s_202), .O(gate383inter1));
  and2  gate2297(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate2298(.a(s_202), .O(gate383inter3));
  inv1  gate2299(.a(s_203), .O(gate383inter4));
  nand2 gate2300(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate2301(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate2302(.a(N1393), .O(gate383inter7));
  inv1  gate2303(.a(N1161), .O(gate383inter8));
  nand2 gate2304(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate2305(.a(s_203), .b(gate383inter3), .O(gate383inter10));
  nor2  gate2306(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate2307(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate2308(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );

  xor2  gate1833(.a(N1444), .b(N939), .O(gate396inter0));
  nand2 gate1834(.a(gate396inter0), .b(s_136), .O(gate396inter1));
  and2  gate1835(.a(N1444), .b(N939), .O(gate396inter2));
  inv1  gate1836(.a(s_136), .O(gate396inter3));
  inv1  gate1837(.a(s_137), .O(gate396inter4));
  nand2 gate1838(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1839(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1840(.a(N939), .O(gate396inter7));
  inv1  gate1841(.a(N1444), .O(gate396inter8));
  nand2 gate1842(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1843(.a(s_137), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1844(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1845(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1846(.a(gate396inter12), .b(gate396inter1), .O(N1487));

  xor2  gate1917(.a(N1446), .b(N935), .O(gate397inter0));
  nand2 gate1918(.a(gate397inter0), .b(s_148), .O(gate397inter1));
  and2  gate1919(.a(N1446), .b(N935), .O(gate397inter2));
  inv1  gate1920(.a(s_148), .O(gate397inter3));
  inv1  gate1921(.a(s_149), .O(gate397inter4));
  nand2 gate1922(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1923(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1924(.a(N935), .O(gate397inter7));
  inv1  gate1925(.a(N1446), .O(gate397inter8));
  nand2 gate1926(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1927(.a(s_149), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1928(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1929(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1930(.a(gate397inter12), .b(gate397inter1), .O(N1488));
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );

  xor2  gate1119(.a(N1468), .b(N965), .O(gate408inter0));
  nand2 gate1120(.a(gate408inter0), .b(s_34), .O(gate408inter1));
  and2  gate1121(.a(N1468), .b(N965), .O(gate408inter2));
  inv1  gate1122(.a(s_34), .O(gate408inter3));
  inv1  gate1123(.a(s_35), .O(gate408inter4));
  nand2 gate1124(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1125(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1126(.a(N965), .O(gate408inter7));
  inv1  gate1127(.a(N1468), .O(gate408inter8));
  nand2 gate1128(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1129(.a(s_35), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1130(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1131(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1132(.a(gate408inter12), .b(gate408inter1), .O(N1500));
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );

  xor2  gate2183(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate2184(.a(gate410inter0), .b(s_186), .O(gate410inter1));
  and2  gate2185(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate2186(.a(s_186), .O(gate410inter3));
  inv1  gate2187(.a(s_187), .O(gate410inter4));
  nand2 gate2188(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2189(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2190(.a(N994), .O(gate410inter7));
  inv1  gate2191(.a(N1475), .O(gate410inter8));
  nand2 gate2192(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2193(.a(s_187), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2194(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2195(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2196(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );

  xor2  gate2029(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate2030(.a(gate413inter0), .b(s_164), .O(gate413inter1));
  and2  gate2031(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate2032(.a(s_164), .O(gate413inter3));
  inv1  gate2033(.a(s_165), .O(gate413inter4));
  nand2 gate2034(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2035(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2036(.a(N1445), .O(gate413inter7));
  inv1  gate2037(.a(N1488), .O(gate413inter8));
  nand2 gate2038(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2039(.a(s_165), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2040(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2041(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2042(.a(gate413inter12), .b(gate413inter1), .O(N1514));
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );

  xor2  gate2225(.a(N1494), .b(N1455), .O(gate417inter0));
  nand2 gate2226(.a(gate417inter0), .b(s_192), .O(gate417inter1));
  and2  gate2227(.a(N1494), .b(N1455), .O(gate417inter2));
  inv1  gate2228(.a(s_192), .O(gate417inter3));
  inv1  gate2229(.a(s_193), .O(gate417inter4));
  nand2 gate2230(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2231(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2232(.a(N1455), .O(gate417inter7));
  inv1  gate2233(.a(N1494), .O(gate417inter8));
  nand2 gate2234(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2235(.a(s_193), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2236(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2237(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2238(.a(gate417inter12), .b(gate417inter1), .O(N1522));

  xor2  gate1567(.a(N1495), .b(N1457), .O(gate418inter0));
  nand2 gate1568(.a(gate418inter0), .b(s_98), .O(gate418inter1));
  and2  gate1569(.a(N1495), .b(N1457), .O(gate418inter2));
  inv1  gate1570(.a(s_98), .O(gate418inter3));
  inv1  gate1571(.a(s_99), .O(gate418inter4));
  nand2 gate1572(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1573(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1574(.a(N1457), .O(gate418inter7));
  inv1  gate1575(.a(N1495), .O(gate418inter8));
  nand2 gate1576(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1577(.a(s_99), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1578(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1579(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1580(.a(gate418inter12), .b(gate418inter1), .O(N1526));
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );

  xor2  gate1945(.a(N1500), .b(N1469), .O(gate426inter0));
  nand2 gate1946(.a(gate426inter0), .b(s_152), .O(gate426inter1));
  and2  gate1947(.a(N1500), .b(N1469), .O(gate426inter2));
  inv1  gate1948(.a(s_152), .O(gate426inter3));
  inv1  gate1949(.a(s_153), .O(gate426inter4));
  nand2 gate1950(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1951(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1952(.a(N1469), .O(gate426inter7));
  inv1  gate1953(.a(N1500), .O(gate426inter8));
  nand2 gate1954(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1955(.a(s_153), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1956(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1957(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1958(.a(gate426inter12), .b(gate426inter1), .O(N1537));
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );

  xor2  gate1217(.a(N1532), .b(N1481), .O(gate433inter0));
  nand2 gate1218(.a(gate433inter0), .b(s_48), .O(gate433inter1));
  and2  gate1219(.a(N1532), .b(N1481), .O(gate433inter2));
  inv1  gate1220(.a(s_48), .O(gate433inter3));
  inv1  gate1221(.a(s_49), .O(gate433inter4));
  nand2 gate1222(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1223(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1224(.a(N1481), .O(gate433inter7));
  inv1  gate1225(.a(N1532), .O(gate433inter8));
  nand2 gate1226(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1227(.a(s_49), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1228(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1229(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1230(.a(gate433inter12), .b(gate433inter1), .O(N1568));
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );

  xor2  gate2197(.a(N1568), .b(N1567), .O(gate442inter0));
  nand2 gate2198(.a(gate442inter0), .b(s_188), .O(gate442inter1));
  and2  gate2199(.a(N1568), .b(N1567), .O(gate442inter2));
  inv1  gate2200(.a(s_188), .O(gate442inter3));
  inv1  gate2201(.a(s_189), .O(gate442inter4));
  nand2 gate2202(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2203(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2204(.a(N1567), .O(gate442inter7));
  inv1  gate2205(.a(N1568), .O(gate442inter8));
  nand2 gate2206(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2207(.a(s_189), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2208(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2209(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2210(.a(gate442inter12), .b(gate442inter1), .O(N1596));
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );

  xor2  gate1427(.a(N1595), .b(N1478), .O(gate452inter0));
  nand2 gate1428(.a(gate452inter0), .b(s_78), .O(gate452inter1));
  and2  gate1429(.a(N1595), .b(N1478), .O(gate452inter2));
  inv1  gate1430(.a(s_78), .O(gate452inter3));
  inv1  gate1431(.a(s_79), .O(gate452inter4));
  nand2 gate1432(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1433(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1434(.a(N1478), .O(gate452inter7));
  inv1  gate1435(.a(N1595), .O(gate452inter8));
  nand2 gate1436(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1437(.a(s_79), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1438(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1439(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1440(.a(gate452inter12), .b(gate452inter1), .O(N1636));

  xor2  gate1903(.a(N1569), .b(N1576), .O(gate453inter0));
  nand2 gate1904(.a(gate453inter0), .b(s_146), .O(gate453inter1));
  and2  gate1905(.a(N1569), .b(N1576), .O(gate453inter2));
  inv1  gate1906(.a(s_146), .O(gate453inter3));
  inv1  gate1907(.a(s_147), .O(gate453inter4));
  nand2 gate1908(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1909(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1910(.a(N1576), .O(gate453inter7));
  inv1  gate1911(.a(N1569), .O(gate453inter8));
  nand2 gate1912(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1913(.a(s_147), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1914(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1915(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1916(.a(gate453inter12), .b(gate453inter1), .O(N1638));
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );

  xor2  gate2337(.a(N1636), .b(N1594), .O(gate472inter0));
  nand2 gate2338(.a(gate472inter0), .b(s_208), .O(gate472inter1));
  and2  gate2339(.a(N1636), .b(N1594), .O(gate472inter2));
  inv1  gate2340(.a(s_208), .O(gate472inter3));
  inv1  gate2341(.a(s_209), .O(gate472inter4));
  nand2 gate2342(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2343(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2344(.a(N1594), .O(gate472inter7));
  inv1  gate2345(.a(N1636), .O(gate472inter8));
  nand2 gate2346(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2347(.a(s_209), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2348(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2349(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2350(.a(gate472inter12), .b(gate472inter1), .O(N1685));

  xor2  gate1203(.a(N1639), .b(N1510), .O(gate473inter0));
  nand2 gate1204(.a(gate473inter0), .b(s_46), .O(gate473inter1));
  and2  gate1205(.a(N1639), .b(N1510), .O(gate473inter2));
  inv1  gate1206(.a(s_46), .O(gate473inter3));
  inv1  gate1207(.a(s_47), .O(gate473inter4));
  nand2 gate1208(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1209(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1210(.a(N1510), .O(gate473inter7));
  inv1  gate1211(.a(N1639), .O(gate473inter8));
  nand2 gate1212(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1213(.a(s_47), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1214(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1215(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1216(.a(gate473inter12), .b(gate473inter1), .O(N1688));
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );

  xor2  gate1553(.a(N1709), .b(N1600), .O(gate497inter0));
  nand2 gate1554(.a(gate497inter0), .b(s_96), .O(gate497inter1));
  and2  gate1555(.a(N1709), .b(N1600), .O(gate497inter2));
  inv1  gate1556(.a(s_96), .O(gate497inter3));
  inv1  gate1557(.a(s_97), .O(gate497inter4));
  nand2 gate1558(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1559(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1560(.a(N1600), .O(gate497inter7));
  inv1  gate1561(.a(N1709), .O(gate497inter8));
  nand2 gate1562(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1563(.a(s_97), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1564(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1565(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1566(.a(gate497inter12), .b(gate497inter1), .O(N1746));
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );

  xor2  gate951(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate952(.a(gate499inter0), .b(s_10), .O(gate499inter1));
  and2  gate953(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate954(.a(s_10), .O(gate499inter3));
  inv1  gate955(.a(s_11), .O(gate499inter4));
  nand2 gate956(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate957(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate958(.a(N1678), .O(gate499inter7));
  inv1  gate959(.a(N1712), .O(gate499inter8));
  nand2 gate960(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate961(.a(s_11), .b(gate499inter3), .O(gate499inter10));
  nor2  gate962(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate963(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate964(.a(gate499inter12), .b(gate499inter1), .O(N1748));
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );

  xor2  gate1021(.a(N1721), .b(N1537), .O(gate501inter0));
  nand2 gate1022(.a(gate501inter0), .b(s_20), .O(gate501inter1));
  and2  gate1023(.a(N1721), .b(N1537), .O(gate501inter2));
  inv1  gate1024(.a(s_20), .O(gate501inter3));
  inv1  gate1025(.a(s_21), .O(gate501inter4));
  nand2 gate1026(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1027(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1028(.a(N1537), .O(gate501inter7));
  inv1  gate1029(.a(N1721), .O(gate501inter8));
  nand2 gate1030(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1031(.a(s_21), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1032(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1033(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1034(.a(gate501inter12), .b(gate501inter1), .O(N1759));
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate1931(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate1932(.a(gate503inter0), .b(s_150), .O(gate503inter1));
  and2  gate1933(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate1934(.a(s_150), .O(gate503inter3));
  inv1  gate1935(.a(s_151), .O(gate503inter4));
  nand2 gate1936(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1937(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1938(.a(N1697), .O(gate503inter7));
  inv1  gate1939(.a(N1727), .O(gate503inter8));
  nand2 gate1940(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1941(.a(s_151), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1942(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1943(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1944(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );

  xor2  gate1581(.a(N1730), .b(N1701), .O(gate505inter0));
  nand2 gate1582(.a(gate505inter0), .b(s_100), .O(gate505inter1));
  and2  gate1583(.a(N1730), .b(N1701), .O(gate505inter2));
  inv1  gate1584(.a(s_100), .O(gate505inter3));
  inv1  gate1585(.a(s_101), .O(gate505inter4));
  nand2 gate1586(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1587(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1588(.a(N1701), .O(gate505inter7));
  inv1  gate1589(.a(N1730), .O(gate505inter8));
  nand2 gate1590(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1591(.a(s_101), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1592(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1593(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1594(.a(gate505inter12), .b(gate505inter1), .O(N1764));
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1329(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1330(.a(gate513inter0), .b(s_64), .O(gate513inter1));
  and2  gate1331(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1332(.a(s_64), .O(gate513inter3));
  inv1  gate1333(.a(s_65), .O(gate513inter4));
  nand2 gate1334(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1335(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1336(.a(N1731), .O(gate513inter7));
  inv1  gate1337(.a(N1682), .O(gate513inter8));
  nand2 gate1338(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1339(.a(s_65), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1340(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1341(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1342(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );

  xor2  gate1287(.a(N1759), .b(N1720), .O(gate517inter0));
  nand2 gate1288(.a(gate517inter0), .b(s_58), .O(gate517inter1));
  and2  gate1289(.a(N1759), .b(N1720), .O(gate517inter2));
  inv1  gate1290(.a(s_58), .O(gate517inter3));
  inv1  gate1291(.a(s_59), .O(gate517inter4));
  nand2 gate1292(.a(gate517inter4), .b(gate517inter3), .O(gate517inter5));
  nor2  gate1293(.a(gate517inter5), .b(gate517inter2), .O(gate517inter6));
  inv1  gate1294(.a(N1720), .O(gate517inter7));
  inv1  gate1295(.a(N1759), .O(gate517inter8));
  nand2 gate1296(.a(gate517inter8), .b(gate517inter7), .O(gate517inter9));
  nand2 gate1297(.a(s_59), .b(gate517inter3), .O(gate517inter10));
  nor2  gate1298(.a(gate517inter10), .b(gate517inter9), .O(gate517inter11));
  nor2  gate1299(.a(gate517inter11), .b(gate517inter6), .O(gate517inter12));
  nand2 gate1300(.a(gate517inter12), .b(gate517inter1), .O(N1788));

  xor2  gate1665(.a(N1761), .b(N1661), .O(gate518inter0));
  nand2 gate1666(.a(gate518inter0), .b(s_112), .O(gate518inter1));
  and2  gate1667(.a(N1761), .b(N1661), .O(gate518inter2));
  inv1  gate1668(.a(s_112), .O(gate518inter3));
  inv1  gate1669(.a(s_113), .O(gate518inter4));
  nand2 gate1670(.a(gate518inter4), .b(gate518inter3), .O(gate518inter5));
  nor2  gate1671(.a(gate518inter5), .b(gate518inter2), .O(gate518inter6));
  inv1  gate1672(.a(N1661), .O(gate518inter7));
  inv1  gate1673(.a(N1761), .O(gate518inter8));
  nand2 gate1674(.a(gate518inter8), .b(gate518inter7), .O(gate518inter9));
  nand2 gate1675(.a(s_113), .b(gate518inter3), .O(gate518inter10));
  nor2  gate1676(.a(gate518inter10), .b(gate518inter9), .O(gate518inter11));
  nor2  gate1677(.a(gate518inter11), .b(gate518inter6), .O(gate518inter12));
  nand2 gate1678(.a(gate518inter12), .b(gate518inter1), .O(N1791));
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate1469(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate1470(.a(gate522inter0), .b(s_84), .O(gate522inter1));
  and2  gate1471(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate1472(.a(s_84), .O(gate522inter3));
  inv1  gate1473(.a(s_85), .O(gate522inter4));
  nand2 gate1474(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate1475(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate1476(.a(N1740), .O(gate522inter7));
  inv1  gate1477(.a(N1769), .O(gate522inter8));
  nand2 gate1478(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate1479(.a(s_85), .b(gate522inter3), .O(gate522inter10));
  nor2  gate1480(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate1481(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate1482(.a(gate522inter12), .b(gate522inter1), .O(N1798));
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );

  xor2  gate1875(.a(N290), .b(N1742), .O(gate524inter0));
  nand2 gate1876(.a(gate524inter0), .b(s_142), .O(gate524inter1));
  and2  gate1877(.a(N290), .b(N1742), .O(gate524inter2));
  inv1  gate1878(.a(s_142), .O(gate524inter3));
  inv1  gate1879(.a(s_143), .O(gate524inter4));
  nand2 gate1880(.a(gate524inter4), .b(gate524inter3), .O(gate524inter5));
  nor2  gate1881(.a(gate524inter5), .b(gate524inter2), .O(gate524inter6));
  inv1  gate1882(.a(N1742), .O(gate524inter7));
  inv1  gate1883(.a(N290), .O(gate524inter8));
  nand2 gate1884(.a(gate524inter8), .b(gate524inter7), .O(gate524inter9));
  nand2 gate1885(.a(s_143), .b(gate524inter3), .O(gate524inter10));
  nor2  gate1886(.a(gate524inter10), .b(gate524inter9), .O(gate524inter11));
  nor2  gate1887(.a(gate524inter11), .b(gate524inter6), .O(gate524inter12));
  nand2 gate1888(.a(gate524inter12), .b(gate524inter1), .O(N1802));
inv1 gate525( .a(N1748), .O(N1807) );

  xor2  gate1525(.a(N1218), .b(N1748), .O(gate526inter0));
  nand2 gate1526(.a(gate526inter0), .b(s_92), .O(gate526inter1));
  and2  gate1527(.a(N1218), .b(N1748), .O(gate526inter2));
  inv1  gate1528(.a(s_92), .O(gate526inter3));
  inv1  gate1529(.a(s_93), .O(gate526inter4));
  nand2 gate1530(.a(gate526inter4), .b(gate526inter3), .O(gate526inter5));
  nor2  gate1531(.a(gate526inter5), .b(gate526inter2), .O(gate526inter6));
  inv1  gate1532(.a(N1748), .O(gate526inter7));
  inv1  gate1533(.a(N1218), .O(gate526inter8));
  nand2 gate1534(.a(gate526inter8), .b(gate526inter7), .O(gate526inter9));
  nand2 gate1535(.a(s_93), .b(gate526inter3), .O(gate526inter10));
  nor2  gate1536(.a(gate526inter10), .b(gate526inter9), .O(gate526inter11));
  nor2  gate1537(.a(gate526inter11), .b(gate526inter6), .O(gate526inter12));
  nand2 gate1538(.a(gate526inter12), .b(gate526inter1), .O(N1808));

  xor2  gate1035(.a(N1783), .b(N1612), .O(gate527inter0));
  nand2 gate1036(.a(gate527inter0), .b(s_22), .O(gate527inter1));
  and2  gate1037(.a(N1783), .b(N1612), .O(gate527inter2));
  inv1  gate1038(.a(s_22), .O(gate527inter3));
  inv1  gate1039(.a(s_23), .O(gate527inter4));
  nand2 gate1040(.a(gate527inter4), .b(gate527inter3), .O(gate527inter5));
  nor2  gate1041(.a(gate527inter5), .b(gate527inter2), .O(gate527inter6));
  inv1  gate1042(.a(N1612), .O(gate527inter7));
  inv1  gate1043(.a(N1783), .O(gate527inter8));
  nand2 gate1044(.a(gate527inter8), .b(gate527inter7), .O(gate527inter9));
  nand2 gate1045(.a(s_23), .b(gate527inter3), .O(gate527inter10));
  nor2  gate1046(.a(gate527inter10), .b(gate527inter9), .O(gate527inter11));
  nor2  gate1047(.a(gate527inter11), .b(gate527inter6), .O(gate527inter12));
  nand2 gate1048(.a(gate527inter12), .b(gate527inter1), .O(N1809));
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );

  xor2  gate1679(.a(N1764), .b(N1792), .O(gate530inter0));
  nand2 gate1680(.a(gate530inter0), .b(s_114), .O(gate530inter1));
  and2  gate1681(.a(N1764), .b(N1792), .O(gate530inter2));
  inv1  gate1682(.a(s_114), .O(gate530inter3));
  inv1  gate1683(.a(s_115), .O(gate530inter4));
  nand2 gate1684(.a(gate530inter4), .b(gate530inter3), .O(gate530inter5));
  nor2  gate1685(.a(gate530inter5), .b(gate530inter2), .O(gate530inter6));
  inv1  gate1686(.a(N1792), .O(gate530inter7));
  inv1  gate1687(.a(N1764), .O(gate530inter8));
  nand2 gate1688(.a(gate530inter8), .b(gate530inter7), .O(gate530inter9));
  nand2 gate1689(.a(s_115), .b(gate530inter3), .O(gate530inter10));
  nor2  gate1690(.a(gate530inter10), .b(gate530inter9), .O(gate530inter11));
  nor2  gate1691(.a(gate530inter11), .b(gate530inter6), .O(gate530inter12));
  nand2 gate1692(.a(gate530inter12), .b(gate530inter1), .O(N1815));
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );

  xor2  gate2309(.a(N1491), .b(N1774), .O(gate534inter0));
  nand2 gate2310(.a(gate534inter0), .b(s_204), .O(gate534inter1));
  and2  gate2311(.a(N1491), .b(N1774), .O(gate534inter2));
  inv1  gate2312(.a(s_204), .O(gate534inter3));
  inv1  gate2313(.a(s_205), .O(gate534inter4));
  nand2 gate2314(.a(gate534inter4), .b(gate534inter3), .O(gate534inter5));
  nor2  gate2315(.a(gate534inter5), .b(gate534inter2), .O(gate534inter6));
  inv1  gate2316(.a(N1774), .O(gate534inter7));
  inv1  gate2317(.a(N1491), .O(gate534inter8));
  nand2 gate2318(.a(gate534inter8), .b(gate534inter7), .O(gate534inter9));
  nand2 gate2319(.a(s_205), .b(gate534inter3), .O(gate534inter10));
  nor2  gate2320(.a(gate534inter10), .b(gate534inter9), .O(gate534inter11));
  nor2  gate2321(.a(gate534inter11), .b(gate534inter6), .O(gate534inter12));
  nand2 gate2322(.a(gate534inter12), .b(gate534inter1), .O(N1823));
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );

  xor2  gate1497(.a(N1801), .b(N1772), .O(gate539inter0));
  nand2 gate1498(.a(gate539inter0), .b(s_88), .O(gate539inter1));
  and2  gate1499(.a(N1801), .b(N1772), .O(gate539inter2));
  inv1  gate1500(.a(s_88), .O(gate539inter3));
  inv1  gate1501(.a(s_89), .O(gate539inter4));
  nand2 gate1502(.a(gate539inter4), .b(gate539inter3), .O(gate539inter5));
  nor2  gate1503(.a(gate539inter5), .b(gate539inter2), .O(gate539inter6));
  inv1  gate1504(.a(N1772), .O(gate539inter7));
  inv1  gate1505(.a(N1801), .O(gate539inter8));
  nand2 gate1506(.a(gate539inter8), .b(gate539inter7), .O(gate539inter9));
  nand2 gate1507(.a(s_89), .b(gate539inter3), .O(gate539inter10));
  nor2  gate1508(.a(gate539inter10), .b(gate539inter9), .O(gate539inter11));
  nor2  gate1509(.a(gate539inter11), .b(gate539inter6), .O(gate539inter12));
  nand2 gate1510(.a(gate539inter12), .b(gate539inter1), .O(N1830));
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );

  xor2  gate1693(.a(N1822), .b(N1419), .O(gate543inter0));
  nand2 gate1694(.a(gate543inter0), .b(s_116), .O(gate543inter1));
  and2  gate1695(.a(N1822), .b(N1419), .O(gate543inter2));
  inv1  gate1696(.a(s_116), .O(gate543inter3));
  inv1  gate1697(.a(s_117), .O(gate543inter4));
  nand2 gate1698(.a(gate543inter4), .b(gate543inter3), .O(gate543inter5));
  nor2  gate1699(.a(gate543inter5), .b(gate543inter2), .O(gate543inter6));
  inv1  gate1700(.a(N1419), .O(gate543inter7));
  inv1  gate1701(.a(N1822), .O(gate543inter8));
  nand2 gate1702(.a(gate543inter8), .b(gate543inter7), .O(gate543inter9));
  nand2 gate1703(.a(s_117), .b(gate543inter3), .O(gate543inter10));
  nor2  gate1704(.a(gate543inter10), .b(gate543inter9), .O(gate543inter11));
  nor2  gate1705(.a(gate543inter11), .b(gate543inter6), .O(gate543inter12));
  nand2 gate1706(.a(gate543inter12), .b(gate543inter1), .O(N1848));

  xor2  gate1511(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate1512(.a(gate544inter0), .b(s_90), .O(gate544inter1));
  and2  gate1513(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate1514(.a(s_90), .O(gate544inter3));
  inv1  gate1515(.a(s_91), .O(gate544inter4));
  nand2 gate1516(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate1517(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate1518(.a(N1416), .O(gate544inter7));
  inv1  gate1519(.a(N1824), .O(gate544inter8));
  nand2 gate1520(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate1521(.a(s_91), .b(gate544inter3), .O(gate544inter10));
  nor2  gate1522(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate1523(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate1524(.a(gate544inter12), .b(gate544inter1), .O(N1849));
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );

  xor2  gate2141(.a(N1848), .b(N1821), .O(gate557inter0));
  nand2 gate2142(.a(gate557inter0), .b(s_180), .O(gate557inter1));
  and2  gate2143(.a(N1848), .b(N1821), .O(gate557inter2));
  inv1  gate2144(.a(s_180), .O(gate557inter3));
  inv1  gate2145(.a(s_181), .O(gate557inter4));
  nand2 gate2146(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate2147(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate2148(.a(N1821), .O(gate557inter7));
  inv1  gate2149(.a(N1848), .O(gate557inter8));
  nand2 gate2150(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate2151(.a(s_181), .b(gate557inter3), .O(gate557inter10));
  nor2  gate2152(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate2153(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate2154(.a(gate557inter12), .b(gate557inter1), .O(N1878));
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );

  xor2  gate1609(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate1610(.a(gate562inter0), .b(s_104), .O(gate562inter1));
  and2  gate1611(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate1612(.a(s_104), .O(gate562inter3));
  inv1  gate1613(.a(s_105), .O(gate562inter4));
  nand2 gate1614(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate1615(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate1616(.a(N1643), .O(gate562inter7));
  inv1  gate1617(.a(N1856), .O(gate562inter8));
  nand2 gate1618(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate1619(.a(s_105), .b(gate562inter3), .O(gate562inter10));
  nor2  gate1620(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate1621(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate1622(.a(gate562inter12), .b(gate562inter1), .O(N1885));
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate2281(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate2282(.a(gate565inter0), .b(s_200), .O(gate565inter1));
  and2  gate2283(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate2284(.a(s_200), .O(gate565inter3));
  inv1  gate2285(.a(s_201), .O(gate565inter4));
  nand2 gate2286(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate2287(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate2288(.a(N1838), .O(gate565inter7));
  inv1  gate2289(.a(N1785), .O(gate565inter8));
  nand2 gate2290(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate2291(.a(s_201), .b(gate565inter3), .O(gate565inter10));
  nor2  gate2292(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate2293(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate2294(.a(gate565inter12), .b(gate565inter1), .O(N1896));

  xor2  gate1175(.a(N1864), .b(N1640), .O(gate566inter0));
  nand2 gate1176(.a(gate566inter0), .b(s_42), .O(gate566inter1));
  and2  gate1177(.a(N1864), .b(N1640), .O(gate566inter2));
  inv1  gate1178(.a(s_42), .O(gate566inter3));
  inv1  gate1179(.a(s_43), .O(gate566inter4));
  nand2 gate1180(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate1181(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate1182(.a(N1640), .O(gate566inter7));
  inv1  gate1183(.a(N1864), .O(gate566inter8));
  nand2 gate1184(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate1185(.a(s_43), .b(gate566inter3), .O(gate566inter10));
  nor2  gate1186(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate1187(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate1188(.a(gate566inter12), .b(gate566inter1), .O(N1897));
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );

  xor2  gate1539(.a(N1897), .b(N1865), .O(gate582inter0));
  nand2 gate1540(.a(gate582inter0), .b(s_94), .O(gate582inter1));
  and2  gate1541(.a(N1897), .b(N1865), .O(gate582inter2));
  inv1  gate1542(.a(s_94), .O(gate582inter3));
  inv1  gate1543(.a(s_95), .O(gate582inter4));
  nand2 gate1544(.a(gate582inter4), .b(gate582inter3), .O(gate582inter5));
  nor2  gate1545(.a(gate582inter5), .b(gate582inter2), .O(gate582inter6));
  inv1  gate1546(.a(N1865), .O(gate582inter7));
  inv1  gate1547(.a(N1897), .O(gate582inter8));
  nand2 gate1548(.a(gate582inter8), .b(gate582inter7), .O(gate582inter9));
  nand2 gate1549(.a(s_95), .b(gate582inter3), .O(gate582inter10));
  nor2  gate1550(.a(gate582inter10), .b(gate582inter9), .O(gate582inter11));
  nor2  gate1551(.a(gate582inter11), .b(gate582inter6), .O(gate582inter12));
  nand2 gate1552(.a(gate582inter12), .b(gate582inter1), .O(N1933));
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate2113(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate2114(.a(gate596inter0), .b(s_176), .O(gate596inter1));
  and2  gate2115(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate2116(.a(s_176), .O(gate596inter3));
  inv1  gate2117(.a(s_177), .O(gate596inter4));
  nand2 gate2118(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate2119(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate2120(.a(N1930), .O(gate596inter7));
  inv1  gate2121(.a(N917), .O(gate596inter8));
  nand2 gate2122(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate2123(.a(s_177), .b(gate596inter3), .O(gate596inter10));
  nor2  gate2124(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate2125(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate2126(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );

  xor2  gate1301(.a(N1941), .b(N1919), .O(gate600inter0));
  nand2 gate1302(.a(gate600inter0), .b(s_60), .O(gate600inter1));
  and2  gate1303(.a(N1941), .b(N1919), .O(gate600inter2));
  inv1  gate1304(.a(s_60), .O(gate600inter3));
  inv1  gate1305(.a(s_61), .O(gate600inter4));
  nand2 gate1306(.a(gate600inter4), .b(gate600inter3), .O(gate600inter5));
  nor2  gate1307(.a(gate600inter5), .b(gate600inter2), .O(gate600inter6));
  inv1  gate1308(.a(N1919), .O(gate600inter7));
  inv1  gate1309(.a(N1941), .O(gate600inter8));
  nand2 gate1310(.a(gate600inter8), .b(gate600inter7), .O(gate600inter9));
  nand2 gate1311(.a(s_61), .b(gate600inter3), .O(gate600inter10));
  nor2  gate1312(.a(gate600inter10), .b(gate600inter9), .O(gate600inter11));
  nor2  gate1313(.a(gate600inter11), .b(gate600inter6), .O(gate600inter12));
  nand2 gate1314(.a(gate600inter12), .b(gate600inter1), .O(N1979));
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );

  xor2  gate2001(.a(N1350), .b(N1953), .O(gate608inter0));
  nand2 gate2002(.a(gate608inter0), .b(s_160), .O(gate608inter1));
  and2  gate2003(.a(N1350), .b(N1953), .O(gate608inter2));
  inv1  gate2004(.a(s_160), .O(gate608inter3));
  inv1  gate2005(.a(s_161), .O(gate608inter4));
  nand2 gate2006(.a(gate608inter4), .b(gate608inter3), .O(gate608inter5));
  nor2  gate2007(.a(gate608inter5), .b(gate608inter2), .O(gate608inter6));
  inv1  gate2008(.a(N1953), .O(gate608inter7));
  inv1  gate2009(.a(N1350), .O(gate608inter8));
  nand2 gate2010(.a(gate608inter8), .b(gate608inter7), .O(gate608inter9));
  nand2 gate2011(.a(s_161), .b(gate608inter3), .O(gate608inter10));
  nor2  gate2012(.a(gate608inter10), .b(gate608inter9), .O(gate608inter11));
  nor2  gate2013(.a(gate608inter11), .b(gate608inter6), .O(gate608inter12));
  nand2 gate2014(.a(gate608inter12), .b(gate608inter1), .O(N2004));
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate2015(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate2016(.a(gate612inter0), .b(s_162), .O(gate612inter1));
  and2  gate2017(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate2018(.a(s_162), .O(gate612inter3));
  inv1  gate2019(.a(s_163), .O(gate612inter4));
  nand2 gate2020(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate2021(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate2022(.a(N673), .O(gate612inter7));
  inv1  gate2023(.a(N1976), .O(gate612inter8));
  nand2 gate2024(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate2025(.a(s_163), .b(gate612inter3), .O(gate612inter10));
  nor2  gate2026(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate2027(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate2028(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );

  xor2  gate1441(.a(N1923), .b(N1958), .O(gate616inter0));
  nand2 gate1442(.a(gate616inter0), .b(s_80), .O(gate616inter1));
  and2  gate1443(.a(N1923), .b(N1958), .O(gate616inter2));
  inv1  gate1444(.a(s_80), .O(gate616inter3));
  inv1  gate1445(.a(s_81), .O(gate616inter4));
  nand2 gate1446(.a(gate616inter4), .b(gate616inter3), .O(gate616inter5));
  nor2  gate1447(.a(gate616inter5), .b(gate616inter2), .O(gate616inter6));
  inv1  gate1448(.a(N1958), .O(gate616inter7));
  inv1  gate1449(.a(N1923), .O(gate616inter8));
  nand2 gate1450(.a(gate616inter8), .b(gate616inter7), .O(gate616inter9));
  nand2 gate1451(.a(s_81), .b(gate616inter3), .O(gate616inter10));
  nor2  gate1452(.a(gate616inter10), .b(gate616inter9), .O(gate616inter11));
  nor2  gate1453(.a(gate616inter11), .b(gate616inter6), .O(gate616inter12));
  nand2 gate1454(.a(gate616inter12), .b(gate616inter1), .O(N2014));
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );

  xor2  gate2253(.a(N2002), .b(N1440), .O(gate624inter0));
  nand2 gate2254(.a(gate624inter0), .b(s_196), .O(gate624inter1));
  and2  gate2255(.a(N2002), .b(N1440), .O(gate624inter2));
  inv1  gate2256(.a(s_196), .O(gate624inter3));
  inv1  gate2257(.a(s_197), .O(gate624inter4));
  nand2 gate2258(.a(gate624inter4), .b(gate624inter3), .O(gate624inter5));
  nor2  gate2259(.a(gate624inter5), .b(gate624inter2), .O(gate624inter6));
  inv1  gate2260(.a(N1440), .O(gate624inter7));
  inv1  gate2261(.a(N2002), .O(gate624inter8));
  nand2 gate2262(.a(gate624inter8), .b(gate624inter7), .O(gate624inter9));
  nand2 gate2263(.a(s_197), .b(gate624inter3), .O(gate624inter10));
  nor2  gate2264(.a(gate624inter10), .b(gate624inter9), .O(gate624inter11));
  nor2  gate2265(.a(gate624inter11), .b(gate624inter6), .O(gate624inter12));
  nand2 gate2266(.a(gate624inter12), .b(gate624inter1), .O(N2023));
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );

  xor2  gate1847(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate1848(.a(gate627inter0), .b(s_138), .O(gate627inter1));
  and2  gate1849(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate1850(.a(s_138), .O(gate627inter3));
  inv1  gate1851(.a(s_139), .O(gate627inter4));
  nand2 gate1852(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate1853(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate1854(.a(N1975), .O(gate627inter7));
  inv1  gate1855(.a(N2008), .O(gate627inter8));
  nand2 gate1856(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate1857(.a(s_139), .b(gate627inter3), .O(gate627inter10));
  nor2  gate1858(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate1859(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate1860(.a(gate627inter12), .b(gate627inter1), .O(N2026));

  xor2  gate1763(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1764(.a(gate628inter0), .b(s_126), .O(gate628inter1));
  and2  gate1765(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1766(.a(s_126), .O(gate628inter3));
  inv1  gate1767(.a(s_127), .O(gate628inter4));
  nand2 gate1768(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1769(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1770(.a(N1977), .O(gate628inter7));
  inv1  gate1771(.a(N2009), .O(gate628inter8));
  nand2 gate1772(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1773(.a(s_127), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1774(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1775(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1776(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate1399(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate1400(.a(gate633inter0), .b(s_74), .O(gate633inter1));
  and2  gate1401(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate1402(.a(s_74), .O(gate633inter3));
  inv1  gate1403(.a(s_75), .O(gate633inter4));
  nand2 gate1404(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate1405(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate1406(.a(N2020), .O(gate633inter7));
  inv1  gate1407(.a(N2000), .O(gate633inter8));
  nand2 gate1408(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate1409(.a(s_75), .b(gate633inter3), .O(gate633inter10));
  nor2  gate1410(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate1411(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate1412(.a(gate633inter12), .b(gate633inter1), .O(N2038));
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );

  xor2  gate1973(.a(N2025), .b(N2006), .O(gate637inter0));
  nand2 gate1974(.a(gate637inter0), .b(s_156), .O(gate637inter1));
  and2  gate1975(.a(N2025), .b(N2006), .O(gate637inter2));
  inv1  gate1976(.a(s_156), .O(gate637inter3));
  inv1  gate1977(.a(s_157), .O(gate637inter4));
  nand2 gate1978(.a(gate637inter4), .b(gate637inter3), .O(gate637inter5));
  nor2  gate1979(.a(gate637inter5), .b(gate637inter2), .O(gate637inter6));
  inv1  gate1980(.a(N2006), .O(gate637inter7));
  inv1  gate1981(.a(N2025), .O(gate637inter8));
  nand2 gate1982(.a(gate637inter8), .b(gate637inter7), .O(gate637inter9));
  nand2 gate1983(.a(s_157), .b(gate637inter3), .O(gate637inter10));
  nor2  gate1984(.a(gate637inter10), .b(gate637inter9), .O(gate637inter11));
  nor2  gate1985(.a(gate637inter11), .b(gate637inter6), .O(gate637inter12));
  nand2 gate1986(.a(gate637inter12), .b(gate637inter1), .O(N2042));
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );

  xor2  gate1483(.a(N290), .b(N2060), .O(gate649inter0));
  nand2 gate1484(.a(gate649inter0), .b(s_86), .O(gate649inter1));
  and2  gate1485(.a(N290), .b(N2060), .O(gate649inter2));
  inv1  gate1486(.a(s_86), .O(gate649inter3));
  inv1  gate1487(.a(s_87), .O(gate649inter4));
  nand2 gate1488(.a(gate649inter4), .b(gate649inter3), .O(gate649inter5));
  nor2  gate1489(.a(gate649inter5), .b(gate649inter2), .O(gate649inter6));
  inv1  gate1490(.a(N2060), .O(gate649inter7));
  inv1  gate1491(.a(N290), .O(gate649inter8));
  nand2 gate1492(.a(gate649inter8), .b(gate649inter7), .O(gate649inter9));
  nand2 gate1493(.a(s_87), .b(gate649inter3), .O(gate649inter10));
  nor2  gate1494(.a(gate649inter10), .b(gate649inter9), .O(gate649inter11));
  nor2  gate1495(.a(gate649inter11), .b(gate649inter6), .O(gate649inter12));
  nand2 gate1496(.a(gate649inter12), .b(gate649inter1), .O(N2078));
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );

  xor2  gate2211(.a(N915), .b(N2151), .O(gate663inter0));
  nand2 gate2212(.a(gate663inter0), .b(s_190), .O(gate663inter1));
  and2  gate2213(.a(N915), .b(N2151), .O(gate663inter2));
  inv1  gate2214(.a(s_190), .O(gate663inter3));
  inv1  gate2215(.a(s_191), .O(gate663inter4));
  nand2 gate2216(.a(gate663inter4), .b(gate663inter3), .O(gate663inter5));
  nor2  gate2217(.a(gate663inter5), .b(gate663inter2), .O(gate663inter6));
  inv1  gate2218(.a(N2151), .O(gate663inter7));
  inv1  gate2219(.a(N915), .O(gate663inter8));
  nand2 gate2220(.a(gate663inter8), .b(gate663inter7), .O(gate663inter9));
  nand2 gate2221(.a(s_191), .b(gate663inter3), .O(gate663inter10));
  nor2  gate2222(.a(gate663inter10), .b(gate663inter9), .O(gate663inter11));
  nor2  gate2223(.a(gate663inter11), .b(gate663inter6), .O(gate663inter12));
  nand2 gate2224(.a(gate663inter12), .b(gate663inter1), .O(N2214));
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate1455(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate1456(.a(gate671inter0), .b(s_82), .O(gate671inter1));
  and2  gate1457(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate1458(.a(s_82), .O(gate671inter3));
  inv1  gate1459(.a(s_83), .O(gate671inter4));
  nand2 gate1460(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate1461(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate1462(.a(N2205), .O(gate671inter7));
  inv1  gate1463(.a(N913), .O(gate671inter8));
  nand2 gate1464(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate1465(.a(s_83), .b(gate671inter3), .O(gate671inter10));
  nor2  gate1466(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate1467(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate1468(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );

  xor2  gate1007(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate1008(.a(gate678inter0), .b(s_18), .O(gate678inter1));
  and2  gate1009(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate1010(.a(s_18), .O(gate678inter3));
  inv1  gate1011(.a(s_19), .O(gate678inter4));
  nand2 gate1012(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate1013(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate1014(.a(N1252), .O(gate678inter7));
  inv1  gate1015(.a(N2225), .O(gate678inter8));
  nand2 gate1016(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate1017(.a(s_19), .b(gate678inter3), .O(gate678inter10));
  nor2  gate1018(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate1019(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate1020(.a(gate678inter12), .b(gate678inter1), .O(N2233));
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );

  xor2  gate1987(.a(N2230), .b(N2214), .O(gate681inter0));
  nand2 gate1988(.a(gate681inter0), .b(s_158), .O(gate681inter1));
  and2  gate1989(.a(N2230), .b(N2214), .O(gate681inter2));
  inv1  gate1990(.a(s_158), .O(gate681inter3));
  inv1  gate1991(.a(s_159), .O(gate681inter4));
  nand2 gate1992(.a(gate681inter4), .b(gate681inter3), .O(gate681inter5));
  nor2  gate1993(.a(gate681inter5), .b(gate681inter2), .O(gate681inter6));
  inv1  gate1994(.a(N2214), .O(gate681inter7));
  inv1  gate1995(.a(N2230), .O(gate681inter8));
  nand2 gate1996(.a(gate681inter8), .b(gate681inter7), .O(gate681inter9));
  nand2 gate1997(.a(s_159), .b(gate681inter3), .O(gate681inter10));
  nor2  gate1998(.a(gate681inter10), .b(gate681inter9), .O(gate681inter11));
  nor2  gate1999(.a(gate681inter11), .b(gate681inter6), .O(gate681inter12));
  nand2 gate2000(.a(gate681inter12), .b(gate681inter1), .O(N2236));
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );

  xor2  gate1861(.a(N535), .b(N2561), .O(gate752inter0));
  nand2 gate1862(.a(gate752inter0), .b(s_140), .O(gate752inter1));
  and2  gate1863(.a(N535), .b(N2561), .O(gate752inter2));
  inv1  gate1864(.a(s_140), .O(gate752inter3));
  inv1  gate1865(.a(s_141), .O(gate752inter4));
  nand2 gate1866(.a(gate752inter4), .b(gate752inter3), .O(gate752inter5));
  nor2  gate1867(.a(gate752inter5), .b(gate752inter2), .O(gate752inter6));
  inv1  gate1868(.a(N2561), .O(gate752inter7));
  inv1  gate1869(.a(N535), .O(gate752inter8));
  nand2 gate1870(.a(gate752inter8), .b(gate752inter7), .O(gate752inter9));
  nand2 gate1871(.a(s_141), .b(gate752inter3), .O(gate752inter10));
  nor2  gate1872(.a(gate752inter10), .b(gate752inter9), .O(gate752inter11));
  nor2  gate1873(.a(gate752inter11), .b(gate752inter6), .O(gate752inter12));
  nand2 gate1874(.a(gate752inter12), .b(gate752inter1), .O(N2671));
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate1147(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate1148(.a(gate754inter0), .b(s_38), .O(gate754inter1));
  and2  gate1149(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate1150(.a(s_38), .O(gate754inter3));
  inv1  gate1151(.a(s_39), .O(gate754inter4));
  nand2 gate1152(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1153(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1154(.a(N2564), .O(gate754inter7));
  inv1  gate1155(.a(N536), .O(gate754inter8));
  nand2 gate1156(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1157(.a(s_39), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1158(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1159(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1160(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );

  xor2  gate993(.a(N2670), .b(N343), .O(gate765inter0));
  nand2 gate994(.a(gate765inter0), .b(s_16), .O(gate765inter1));
  and2  gate995(.a(N2670), .b(N343), .O(gate765inter2));
  inv1  gate996(.a(s_16), .O(gate765inter3));
  inv1  gate997(.a(s_17), .O(gate765inter4));
  nand2 gate998(.a(gate765inter4), .b(gate765inter3), .O(gate765inter5));
  nor2  gate999(.a(gate765inter5), .b(gate765inter2), .O(gate765inter6));
  inv1  gate1000(.a(N343), .O(gate765inter7));
  inv1  gate1001(.a(N2670), .O(gate765inter8));
  nand2 gate1002(.a(gate765inter8), .b(gate765inter7), .O(gate765inter9));
  nand2 gate1003(.a(s_17), .b(gate765inter3), .O(gate765inter10));
  nor2  gate1004(.a(gate765inter10), .b(gate765inter9), .O(gate765inter11));
  nor2  gate1005(.a(gate765inter11), .b(gate765inter6), .O(gate765inter12));
  nand2 gate1006(.a(gate765inter12), .b(gate765inter1), .O(N2720));
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );

  xor2  gate1189(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate1190(.a(gate768inter0), .b(s_44), .O(gate768inter1));
  and2  gate1191(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate1192(.a(s_44), .O(gate768inter3));
  inv1  gate1193(.a(s_45), .O(gate768inter4));
  nand2 gate1194(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate1195(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate1196(.a(N352), .O(gate768inter7));
  inv1  gate1197(.a(N2676), .O(gate768inter8));
  nand2 gate1198(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate1199(.a(s_45), .b(gate768inter3), .O(gate768inter10));
  nor2  gate1200(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate1201(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate1202(.a(gate768inter12), .b(gate768inter1), .O(N2723));
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );

  xor2  gate2351(.a(N539), .b(N2642), .O(gate771inter0));
  nand2 gate2352(.a(gate771inter0), .b(s_210), .O(gate771inter1));
  and2  gate2353(.a(N539), .b(N2642), .O(gate771inter2));
  inv1  gate2354(.a(s_210), .O(gate771inter3));
  inv1  gate2355(.a(s_211), .O(gate771inter4));
  nand2 gate2356(.a(gate771inter4), .b(gate771inter3), .O(gate771inter5));
  nor2  gate2357(.a(gate771inter5), .b(gate771inter2), .O(gate771inter6));
  inv1  gate2358(.a(N2642), .O(gate771inter7));
  inv1  gate2359(.a(N539), .O(gate771inter8));
  nand2 gate2360(.a(gate771inter8), .b(gate771inter7), .O(gate771inter9));
  nand2 gate2361(.a(s_211), .b(gate771inter3), .O(gate771inter10));
  nor2  gate2362(.a(gate771inter10), .b(gate771inter9), .O(gate771inter11));
  nor2  gate2363(.a(gate771inter11), .b(gate771inter6), .O(gate771inter12));
  nand2 gate2364(.a(gate771inter12), .b(gate771inter1), .O(N2726));
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate1805(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate1806(.a(gate773inter0), .b(s_132), .O(gate773inter1));
  and2  gate1807(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate1808(.a(s_132), .O(gate773inter3));
  inv1  gate1809(.a(s_133), .O(gate773inter4));
  nand2 gate1810(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate1811(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate1812(.a(N2645), .O(gate773inter7));
  inv1  gate1813(.a(N540), .O(gate773inter8));
  nand2 gate1814(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate1815(.a(s_133), .b(gate773inter3), .O(gate773inter10));
  nor2  gate1816(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate1817(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate1818(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );

  xor2  gate2043(.a(N542), .b(N2651), .O(gate777inter0));
  nand2 gate2044(.a(gate777inter0), .b(s_166), .O(gate777inter1));
  and2  gate2045(.a(N542), .b(N2651), .O(gate777inter2));
  inv1  gate2046(.a(s_166), .O(gate777inter3));
  inv1  gate2047(.a(s_167), .O(gate777inter4));
  nand2 gate2048(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate2049(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate2050(.a(N2651), .O(gate777inter7));
  inv1  gate2051(.a(N542), .O(gate777inter8));
  nand2 gate2052(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate2053(.a(s_167), .b(gate777inter3), .O(gate777inter10));
  nor2  gate2054(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate2055(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate2056(.a(gate777inter12), .b(gate777inter1), .O(N2732));
inv1 gate778( .a(N2651), .O(N2733) );

  xor2  gate2155(.a(N2683), .b(N370), .O(gate779inter0));
  nand2 gate2156(.a(gate779inter0), .b(s_182), .O(gate779inter1));
  and2  gate2157(.a(N2683), .b(N370), .O(gate779inter2));
  inv1  gate2158(.a(s_182), .O(gate779inter3));
  inv1  gate2159(.a(s_183), .O(gate779inter4));
  nand2 gate2160(.a(gate779inter4), .b(gate779inter3), .O(gate779inter5));
  nor2  gate2161(.a(gate779inter5), .b(gate779inter2), .O(gate779inter6));
  inv1  gate2162(.a(N370), .O(gate779inter7));
  inv1  gate2163(.a(N2683), .O(gate779inter8));
  nand2 gate2164(.a(gate779inter8), .b(gate779inter7), .O(gate779inter9));
  nand2 gate2165(.a(s_183), .b(gate779inter3), .O(gate779inter10));
  nor2  gate2166(.a(gate779inter10), .b(gate779inter9), .O(gate779inter11));
  nor2  gate2167(.a(gate779inter11), .b(gate779inter6), .O(gate779inter12));
  nand2 gate2168(.a(gate779inter12), .b(gate779inter1), .O(N2734));
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );

  xor2  gate1735(.a(N547), .b(N2664), .O(gate786inter0));
  nand2 gate1736(.a(gate786inter0), .b(s_122), .O(gate786inter1));
  and2  gate1737(.a(N547), .b(N2664), .O(gate786inter2));
  inv1  gate1738(.a(s_122), .O(gate786inter3));
  inv1  gate1739(.a(s_123), .O(gate786inter4));
  nand2 gate1740(.a(gate786inter4), .b(gate786inter3), .O(gate786inter5));
  nor2  gate1741(.a(gate786inter5), .b(gate786inter2), .O(gate786inter6));
  inv1  gate1742(.a(N2664), .O(gate786inter7));
  inv1  gate1743(.a(N547), .O(gate786inter8));
  nand2 gate1744(.a(gate786inter8), .b(gate786inter7), .O(gate786inter9));
  nand2 gate1745(.a(s_123), .b(gate786inter3), .O(gate786inter10));
  nor2  gate1746(.a(gate786inter10), .b(gate786inter9), .O(gate786inter11));
  nor2  gate1747(.a(gate786inter11), .b(gate786inter6), .O(gate786inter12));
  nand2 gate1748(.a(gate786inter12), .b(gate786inter1), .O(N2741));
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );

  xor2  gate1357(.a(N2720), .b(N2669), .O(gate794inter0));
  nand2 gate1358(.a(gate794inter0), .b(s_68), .O(gate794inter1));
  and2  gate1359(.a(N2720), .b(N2669), .O(gate794inter2));
  inv1  gate1360(.a(s_68), .O(gate794inter3));
  inv1  gate1361(.a(s_69), .O(gate794inter4));
  nand2 gate1362(.a(gate794inter4), .b(gate794inter3), .O(gate794inter5));
  nor2  gate1363(.a(gate794inter5), .b(gate794inter2), .O(gate794inter6));
  inv1  gate1364(.a(N2669), .O(gate794inter7));
  inv1  gate1365(.a(N2720), .O(gate794inter8));
  nand2 gate1366(.a(gate794inter8), .b(gate794inter7), .O(gate794inter9));
  nand2 gate1367(.a(s_69), .b(gate794inter3), .O(gate794inter10));
  nor2  gate1368(.a(gate794inter10), .b(gate794inter9), .O(gate794inter11));
  nor2  gate1369(.a(gate794inter11), .b(gate794inter6), .O(gate794inter12));
  nand2 gate1370(.a(gate794inter12), .b(gate794inter1), .O(N2753));
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );

  xor2  gate1889(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate1890(.a(gate799inter0), .b(s_144), .O(gate799inter1));
  and2  gate1891(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate1892(.a(s_144), .O(gate799inter3));
  inv1  gate1893(.a(s_145), .O(gate799inter4));
  nand2 gate1894(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate1895(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate1896(.a(N358), .O(gate799inter7));
  inv1  gate1897(.a(N2727), .O(gate799inter8));
  nand2 gate1898(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate1899(.a(s_145), .b(gate799inter3), .O(gate799inter10));
  nor2  gate1900(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate1901(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate1902(.a(gate799inter12), .b(gate799inter1), .O(N2758));
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );

  xor2  gate1343(.a(N2733), .b(N367), .O(gate802inter0));
  nand2 gate1344(.a(gate802inter0), .b(s_66), .O(gate802inter1));
  and2  gate1345(.a(N2733), .b(N367), .O(gate802inter2));
  inv1  gate1346(.a(s_66), .O(gate802inter3));
  inv1  gate1347(.a(s_67), .O(gate802inter4));
  nand2 gate1348(.a(gate802inter4), .b(gate802inter3), .O(gate802inter5));
  nor2  gate1349(.a(gate802inter5), .b(gate802inter2), .O(gate802inter6));
  inv1  gate1350(.a(N367), .O(gate802inter7));
  inv1  gate1351(.a(N2733), .O(gate802inter8));
  nand2 gate1352(.a(gate802inter8), .b(gate802inter7), .O(gate802inter9));
  nand2 gate1353(.a(s_67), .b(gate802inter3), .O(gate802inter10));
  nor2  gate1354(.a(gate802inter10), .b(gate802inter9), .O(gate802inter11));
  nor2  gate1355(.a(gate802inter11), .b(gate802inter6), .O(gate802inter12));
  nand2 gate1356(.a(gate802inter12), .b(gate802inter1), .O(N2761));
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );

  xor2  gate2169(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate2170(.a(gate806inter0), .b(s_184), .O(gate806inter1));
  and2  gate2171(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate2172(.a(s_184), .O(gate806inter3));
  inv1  gate2173(.a(s_185), .O(gate806inter4));
  nand2 gate2174(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate2175(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate2176(.a(N379), .O(gate806inter7));
  inv1  gate2177(.a(N2740), .O(gate806inter8));
  nand2 gate2178(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate2179(.a(s_185), .b(gate806inter3), .O(gate806inter10));
  nor2  gate2180(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate2181(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate2182(.a(gate806inter12), .b(gate806inter1), .O(N2765));
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );

  xor2  gate909(.a(N2743), .b(N2688), .O(gate808inter0));
  nand2 gate910(.a(gate808inter0), .b(s_4), .O(gate808inter1));
  and2  gate911(.a(N2743), .b(N2688), .O(gate808inter2));
  inv1  gate912(.a(s_4), .O(gate808inter3));
  inv1  gate913(.a(s_5), .O(gate808inter4));
  nand2 gate914(.a(gate808inter4), .b(gate808inter3), .O(gate808inter5));
  nor2  gate915(.a(gate808inter5), .b(gate808inter2), .O(gate808inter6));
  inv1  gate916(.a(N2688), .O(gate808inter7));
  inv1  gate917(.a(N2743), .O(gate808inter8));
  nand2 gate918(.a(gate808inter8), .b(gate808inter7), .O(gate808inter9));
  nand2 gate919(.a(s_5), .b(gate808inter3), .O(gate808inter10));
  nor2  gate920(.a(gate808inter10), .b(gate808inter9), .O(gate808inter11));
  nor2  gate921(.a(gate808inter11), .b(gate808inter6), .O(gate808inter12));
  nand2 gate922(.a(gate808inter12), .b(gate808inter1), .O(N2767));

  xor2  gate1651(.a(N2744), .b(N2690), .O(gate809inter0));
  nand2 gate1652(.a(gate809inter0), .b(s_110), .O(gate809inter1));
  and2  gate1653(.a(N2744), .b(N2690), .O(gate809inter2));
  inv1  gate1654(.a(s_110), .O(gate809inter3));
  inv1  gate1655(.a(s_111), .O(gate809inter4));
  nand2 gate1656(.a(gate809inter4), .b(gate809inter3), .O(gate809inter5));
  nor2  gate1657(.a(gate809inter5), .b(gate809inter2), .O(gate809inter6));
  inv1  gate1658(.a(N2690), .O(gate809inter7));
  inv1  gate1659(.a(N2744), .O(gate809inter8));
  nand2 gate1660(.a(gate809inter8), .b(gate809inter7), .O(gate809inter9));
  nand2 gate1661(.a(s_111), .b(gate809inter3), .O(gate809inter10));
  nor2  gate1662(.a(gate809inter10), .b(gate809inter9), .O(gate809inter11));
  nor2  gate1663(.a(gate809inter11), .b(gate809inter6), .O(gate809inter12));
  nand2 gate1664(.a(gate809inter12), .b(gate809inter1), .O(N2768));
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );

  xor2  gate2239(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate2240(.a(gate815inter0), .b(s_194), .O(gate815inter1));
  and2  gate2241(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate2242(.a(s_194), .O(gate815inter3));
  inv1  gate2243(.a(s_195), .O(gate815inter4));
  nand2 gate2244(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate2245(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate2246(.a(N2730), .O(gate815inter7));
  inv1  gate2247(.a(N2760), .O(gate815inter8));
  nand2 gate2248(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate2249(.a(s_195), .b(gate815inter3), .O(gate815inter10));
  nor2  gate2250(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate2251(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate2252(.a(gate815inter12), .b(gate815inter1), .O(N2782));
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );

  xor2  gate1245(.a(N2764), .b(N2737), .O(gate818inter0));
  nand2 gate1246(.a(gate818inter0), .b(s_52), .O(gate818inter1));
  and2  gate1247(.a(N2764), .b(N2737), .O(gate818inter2));
  inv1  gate1248(.a(s_52), .O(gate818inter3));
  inv1  gate1249(.a(s_53), .O(gate818inter4));
  nand2 gate1250(.a(gate818inter4), .b(gate818inter3), .O(gate818inter5));
  nor2  gate1251(.a(gate818inter5), .b(gate818inter2), .O(gate818inter6));
  inv1  gate1252(.a(N2737), .O(gate818inter7));
  inv1  gate1253(.a(N2764), .O(gate818inter8));
  nand2 gate1254(.a(gate818inter8), .b(gate818inter7), .O(gate818inter9));
  nand2 gate1255(.a(s_53), .b(gate818inter3), .O(gate818inter10));
  nor2  gate1256(.a(gate818inter10), .b(gate818inter9), .O(gate818inter11));
  nor2  gate1257(.a(gate818inter11), .b(gate818inter6), .O(gate818inter12));
  nand2 gate1258(.a(gate818inter12), .b(gate818inter1), .O(N2785));
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );

  xor2  gate2127(.a(N2800), .b(N2384), .O(gate828inter0));
  nand2 gate2128(.a(gate828inter0), .b(s_178), .O(gate828inter1));
  and2  gate2129(.a(N2800), .b(N2384), .O(gate828inter2));
  inv1  gate2130(.a(s_178), .O(gate828inter3));
  inv1  gate2131(.a(s_179), .O(gate828inter4));
  nand2 gate2132(.a(gate828inter4), .b(gate828inter3), .O(gate828inter5));
  nor2  gate2133(.a(gate828inter5), .b(gate828inter2), .O(gate828inter6));
  inv1  gate2134(.a(N2384), .O(gate828inter7));
  inv1  gate2135(.a(N2800), .O(gate828inter8));
  nand2 gate2136(.a(gate828inter8), .b(gate828inter7), .O(gate828inter9));
  nand2 gate2137(.a(s_179), .b(gate828inter3), .O(gate828inter10));
  nor2  gate2138(.a(gate828inter10), .b(gate828inter9), .O(gate828inter11));
  nor2  gate2139(.a(gate828inter11), .b(gate828inter6), .O(gate828inter12));
  nand2 gate2140(.a(gate828inter12), .b(gate828inter1), .O(N2811));
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );

  xor2  gate1707(.a(N2828), .b(N2809), .O(gate838inter0));
  nand2 gate1708(.a(gate838inter0), .b(s_118), .O(gate838inter1));
  and2  gate1709(.a(N2828), .b(N2809), .O(gate838inter2));
  inv1  gate1710(.a(s_118), .O(gate838inter3));
  inv1  gate1711(.a(s_119), .O(gate838inter4));
  nand2 gate1712(.a(gate838inter4), .b(gate838inter3), .O(gate838inter5));
  nor2  gate1713(.a(gate838inter5), .b(gate838inter2), .O(gate838inter6));
  inv1  gate1714(.a(N2809), .O(gate838inter7));
  inv1  gate1715(.a(N2828), .O(gate838inter8));
  nand2 gate1716(.a(gate838inter8), .b(gate838inter7), .O(gate838inter9));
  nand2 gate1717(.a(s_119), .b(gate838inter3), .O(gate838inter10));
  nor2  gate1718(.a(gate838inter10), .b(gate838inter9), .O(gate838inter11));
  nor2  gate1719(.a(gate838inter11), .b(gate838inter6), .O(gate838inter12));
  nand2 gate1720(.a(gate838inter12), .b(gate838inter1), .O(N2846));

  xor2  gate2071(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate2072(.a(gate839inter0), .b(s_170), .O(gate839inter1));
  and2  gate2073(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate2074(.a(s_170), .O(gate839inter3));
  inv1  gate2075(.a(s_171), .O(gate839inter4));
  nand2 gate2076(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate2077(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate2078(.a(N2812), .O(gate839inter7));
  inv1  gate2079(.a(N2076), .O(gate839inter8));
  nand2 gate2080(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate2081(.a(s_171), .b(gate839inter3), .O(gate839inter10));
  nor2  gate2082(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate2083(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate2084(.a(gate839inter12), .b(gate839inter1), .O(N2850));

  xor2  gate1161(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate1162(.a(gate840inter0), .b(s_40), .O(gate840inter1));
  and2  gate1163(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate1164(.a(s_40), .O(gate840inter3));
  inv1  gate1165(.a(s_41), .O(gate840inter4));
  nand2 gate1166(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate1167(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate1168(.a(N2815), .O(gate840inter7));
  inv1  gate1169(.a(N2077), .O(gate840inter8));
  nand2 gate1170(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate1171(.a(s_41), .b(gate840inter3), .O(gate840inter10));
  nor2  gate1172(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate1173(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate1174(.a(gate840inter12), .b(gate840inter1), .O(N2851));
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );

  xor2  gate895(.a(N887), .b(N2846), .O(gate858inter0));
  nand2 gate896(.a(gate858inter0), .b(s_2), .O(gate858inter1));
  and2  gate897(.a(N887), .b(N2846), .O(gate858inter2));
  inv1  gate898(.a(s_2), .O(gate858inter3));
  inv1  gate899(.a(s_3), .O(gate858inter4));
  nand2 gate900(.a(gate858inter4), .b(gate858inter3), .O(gate858inter5));
  nor2  gate901(.a(gate858inter5), .b(gate858inter2), .O(gate858inter6));
  inv1  gate902(.a(N2846), .O(gate858inter7));
  inv1  gate903(.a(N887), .O(gate858inter8));
  nand2 gate904(.a(gate858inter8), .b(gate858inter7), .O(gate858inter9));
  nand2 gate905(.a(s_3), .b(gate858inter3), .O(gate858inter10));
  nor2  gate906(.a(gate858inter10), .b(gate858inter9), .O(gate858inter11));
  nor2  gate907(.a(gate858inter11), .b(gate858inter6), .O(gate858inter12));
  nand2 gate908(.a(gate858inter12), .b(gate858inter1), .O(N2873));
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );

  xor2  gate1777(.a(N2850), .b(N2866), .O(gate861inter0));
  nand2 gate1778(.a(gate861inter0), .b(s_128), .O(gate861inter1));
  and2  gate1779(.a(N2850), .b(N2866), .O(gate861inter2));
  inv1  gate1780(.a(s_128), .O(gate861inter3));
  inv1  gate1781(.a(s_129), .O(gate861inter4));
  nand2 gate1782(.a(gate861inter4), .b(gate861inter3), .O(gate861inter5));
  nor2  gate1783(.a(gate861inter5), .b(gate861inter2), .O(gate861inter6));
  inv1  gate1784(.a(N2866), .O(gate861inter7));
  inv1  gate1785(.a(N2850), .O(gate861inter8));
  nand2 gate1786(.a(gate861inter8), .b(gate861inter7), .O(gate861inter9));
  nand2 gate1787(.a(s_129), .b(gate861inter3), .O(gate861inter10));
  nor2  gate1788(.a(gate861inter10), .b(gate861inter9), .O(gate861inter11));
  nor2  gate1789(.a(gate861inter11), .b(gate861inter6), .O(gate861inter12));
  nand2 gate1790(.a(gate861inter12), .b(gate861inter1), .O(N2876));
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );

  xor2  gate937(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate938(.a(gate865inter0), .b(s_8), .O(gate865inter1));
  and2  gate939(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate940(.a(s_8), .O(gate865inter3));
  inv1  gate941(.a(s_9), .O(gate865inter4));
  nand2 gate942(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate943(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate944(.a(N2870), .O(gate865inter7));
  inv1  gate945(.a(N2854), .O(gate865inter8));
  nand2 gate946(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate947(.a(s_9), .b(gate865inter3), .O(gate865inter10));
  nor2  gate948(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate949(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate950(.a(gate865inter12), .b(gate865inter1), .O(N2880));
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule