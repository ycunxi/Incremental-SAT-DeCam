module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate547(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate548(.a(gate10inter0), .b(s_0), .O(gate10inter1));
  and2  gate549(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate550(.a(s_0), .O(gate10inter3));
  inv1  gate551(.a(s_1), .O(gate10inter4));
  nand2 gate552(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate553(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate554(.a(G3), .O(gate10inter7));
  inv1  gate555(.a(G4), .O(gate10inter8));
  nand2 gate556(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate557(.a(s_1), .b(gate10inter3), .O(gate10inter10));
  nor2  gate558(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate559(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate560(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1765(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1766(.a(gate18inter0), .b(s_174), .O(gate18inter1));
  and2  gate1767(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1768(.a(s_174), .O(gate18inter3));
  inv1  gate1769(.a(s_175), .O(gate18inter4));
  nand2 gate1770(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1771(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1772(.a(G19), .O(gate18inter7));
  inv1  gate1773(.a(G20), .O(gate18inter8));
  nand2 gate1774(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1775(.a(s_175), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1776(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1777(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1778(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1163(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1164(.a(gate20inter0), .b(s_88), .O(gate20inter1));
  and2  gate1165(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1166(.a(s_88), .O(gate20inter3));
  inv1  gate1167(.a(s_89), .O(gate20inter4));
  nand2 gate1168(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1169(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1170(.a(G23), .O(gate20inter7));
  inv1  gate1171(.a(G24), .O(gate20inter8));
  nand2 gate1172(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1173(.a(s_89), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1174(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1175(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1176(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1429(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1430(.a(gate40inter0), .b(s_126), .O(gate40inter1));
  and2  gate1431(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1432(.a(s_126), .O(gate40inter3));
  inv1  gate1433(.a(s_127), .O(gate40inter4));
  nand2 gate1434(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1435(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1436(.a(G28), .O(gate40inter7));
  inv1  gate1437(.a(G32), .O(gate40inter8));
  nand2 gate1438(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1439(.a(s_127), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1440(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1441(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1442(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1863(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1864(.a(gate41inter0), .b(s_188), .O(gate41inter1));
  and2  gate1865(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1866(.a(s_188), .O(gate41inter3));
  inv1  gate1867(.a(s_189), .O(gate41inter4));
  nand2 gate1868(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1869(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1870(.a(G1), .O(gate41inter7));
  inv1  gate1871(.a(G266), .O(gate41inter8));
  nand2 gate1872(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1873(.a(s_189), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1874(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1875(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1876(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1135(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1136(.a(gate42inter0), .b(s_84), .O(gate42inter1));
  and2  gate1137(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1138(.a(s_84), .O(gate42inter3));
  inv1  gate1139(.a(s_85), .O(gate42inter4));
  nand2 gate1140(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1141(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1142(.a(G2), .O(gate42inter7));
  inv1  gate1143(.a(G266), .O(gate42inter8));
  nand2 gate1144(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1145(.a(s_85), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1146(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1147(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1148(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1625(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1626(.a(gate44inter0), .b(s_154), .O(gate44inter1));
  and2  gate1627(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1628(.a(s_154), .O(gate44inter3));
  inv1  gate1629(.a(s_155), .O(gate44inter4));
  nand2 gate1630(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1631(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1632(.a(G4), .O(gate44inter7));
  inv1  gate1633(.a(G269), .O(gate44inter8));
  nand2 gate1634(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1635(.a(s_155), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1636(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1637(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1638(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1471(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1472(.a(gate52inter0), .b(s_132), .O(gate52inter1));
  and2  gate1473(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1474(.a(s_132), .O(gate52inter3));
  inv1  gate1475(.a(s_133), .O(gate52inter4));
  nand2 gate1476(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1477(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1478(.a(G12), .O(gate52inter7));
  inv1  gate1479(.a(G281), .O(gate52inter8));
  nand2 gate1480(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1481(.a(s_133), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1482(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1483(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1484(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate715(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate716(.a(gate55inter0), .b(s_24), .O(gate55inter1));
  and2  gate717(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate718(.a(s_24), .O(gate55inter3));
  inv1  gate719(.a(s_25), .O(gate55inter4));
  nand2 gate720(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate721(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate722(.a(G15), .O(gate55inter7));
  inv1  gate723(.a(G287), .O(gate55inter8));
  nand2 gate724(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate725(.a(s_25), .b(gate55inter3), .O(gate55inter10));
  nor2  gate726(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate727(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate728(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate645(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate646(.a(gate59inter0), .b(s_14), .O(gate59inter1));
  and2  gate647(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate648(.a(s_14), .O(gate59inter3));
  inv1  gate649(.a(s_15), .O(gate59inter4));
  nand2 gate650(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate651(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate652(.a(G19), .O(gate59inter7));
  inv1  gate653(.a(G293), .O(gate59inter8));
  nand2 gate654(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate655(.a(s_15), .b(gate59inter3), .O(gate59inter10));
  nor2  gate656(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate657(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate658(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate617(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate618(.a(gate63inter0), .b(s_10), .O(gate63inter1));
  and2  gate619(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate620(.a(s_10), .O(gate63inter3));
  inv1  gate621(.a(s_11), .O(gate63inter4));
  nand2 gate622(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate623(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate624(.a(G23), .O(gate63inter7));
  inv1  gate625(.a(G299), .O(gate63inter8));
  nand2 gate626(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate627(.a(s_11), .b(gate63inter3), .O(gate63inter10));
  nor2  gate628(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate629(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate630(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1345(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1346(.a(gate64inter0), .b(s_114), .O(gate64inter1));
  and2  gate1347(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1348(.a(s_114), .O(gate64inter3));
  inv1  gate1349(.a(s_115), .O(gate64inter4));
  nand2 gate1350(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1351(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1352(.a(G24), .O(gate64inter7));
  inv1  gate1353(.a(G299), .O(gate64inter8));
  nand2 gate1354(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1355(.a(s_115), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1356(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1357(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1358(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate799(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate800(.a(gate71inter0), .b(s_36), .O(gate71inter1));
  and2  gate801(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate802(.a(s_36), .O(gate71inter3));
  inv1  gate803(.a(s_37), .O(gate71inter4));
  nand2 gate804(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate805(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate806(.a(G31), .O(gate71inter7));
  inv1  gate807(.a(G311), .O(gate71inter8));
  nand2 gate808(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate809(.a(s_37), .b(gate71inter3), .O(gate71inter10));
  nor2  gate810(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate811(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate812(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1541(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1542(.a(gate72inter0), .b(s_142), .O(gate72inter1));
  and2  gate1543(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1544(.a(s_142), .O(gate72inter3));
  inv1  gate1545(.a(s_143), .O(gate72inter4));
  nand2 gate1546(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1547(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1548(.a(G32), .O(gate72inter7));
  inv1  gate1549(.a(G311), .O(gate72inter8));
  nand2 gate1550(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1551(.a(s_143), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1552(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1553(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1554(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate897(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate898(.a(gate75inter0), .b(s_50), .O(gate75inter1));
  and2  gate899(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate900(.a(s_50), .O(gate75inter3));
  inv1  gate901(.a(s_51), .O(gate75inter4));
  nand2 gate902(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate903(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate904(.a(G9), .O(gate75inter7));
  inv1  gate905(.a(G317), .O(gate75inter8));
  nand2 gate906(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate907(.a(s_51), .b(gate75inter3), .O(gate75inter10));
  nor2  gate908(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate909(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate910(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate701(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate702(.a(gate78inter0), .b(s_22), .O(gate78inter1));
  and2  gate703(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate704(.a(s_22), .O(gate78inter3));
  inv1  gate705(.a(s_23), .O(gate78inter4));
  nand2 gate706(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate707(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate708(.a(G6), .O(gate78inter7));
  inv1  gate709(.a(G320), .O(gate78inter8));
  nand2 gate710(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate711(.a(s_23), .b(gate78inter3), .O(gate78inter10));
  nor2  gate712(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate713(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate714(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate813(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate814(.a(gate87inter0), .b(s_38), .O(gate87inter1));
  and2  gate815(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate816(.a(s_38), .O(gate87inter3));
  inv1  gate817(.a(s_39), .O(gate87inter4));
  nand2 gate818(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate819(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate820(.a(G12), .O(gate87inter7));
  inv1  gate821(.a(G335), .O(gate87inter8));
  nand2 gate822(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate823(.a(s_39), .b(gate87inter3), .O(gate87inter10));
  nor2  gate824(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate825(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate826(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1709(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1710(.a(gate89inter0), .b(s_166), .O(gate89inter1));
  and2  gate1711(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1712(.a(s_166), .O(gate89inter3));
  inv1  gate1713(.a(s_167), .O(gate89inter4));
  nand2 gate1714(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1715(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1716(.a(G17), .O(gate89inter7));
  inv1  gate1717(.a(G338), .O(gate89inter8));
  nand2 gate1718(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1719(.a(s_167), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1720(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1721(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1722(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1835(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1836(.a(gate98inter0), .b(s_184), .O(gate98inter1));
  and2  gate1837(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1838(.a(s_184), .O(gate98inter3));
  inv1  gate1839(.a(s_185), .O(gate98inter4));
  nand2 gate1840(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1841(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1842(.a(G23), .O(gate98inter7));
  inv1  gate1843(.a(G350), .O(gate98inter8));
  nand2 gate1844(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1845(.a(s_185), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1846(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1847(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1848(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate995(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate996(.a(gate100inter0), .b(s_64), .O(gate100inter1));
  and2  gate997(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate998(.a(s_64), .O(gate100inter3));
  inv1  gate999(.a(s_65), .O(gate100inter4));
  nand2 gate1000(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1001(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1002(.a(G31), .O(gate100inter7));
  inv1  gate1003(.a(G353), .O(gate100inter8));
  nand2 gate1004(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1005(.a(s_65), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1006(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1007(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1008(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1653(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1654(.a(gate101inter0), .b(s_158), .O(gate101inter1));
  and2  gate1655(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1656(.a(s_158), .O(gate101inter3));
  inv1  gate1657(.a(s_159), .O(gate101inter4));
  nand2 gate1658(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1659(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1660(.a(G20), .O(gate101inter7));
  inv1  gate1661(.a(G356), .O(gate101inter8));
  nand2 gate1662(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1663(.a(s_159), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1664(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1665(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1666(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1177(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1178(.a(gate104inter0), .b(s_90), .O(gate104inter1));
  and2  gate1179(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1180(.a(s_90), .O(gate104inter3));
  inv1  gate1181(.a(s_91), .O(gate104inter4));
  nand2 gate1182(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1183(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1184(.a(G32), .O(gate104inter7));
  inv1  gate1185(.a(G359), .O(gate104inter8));
  nand2 gate1186(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1187(.a(s_91), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1188(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1189(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1190(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate673(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate674(.a(gate106inter0), .b(s_18), .O(gate106inter1));
  and2  gate675(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate676(.a(s_18), .O(gate106inter3));
  inv1  gate677(.a(s_19), .O(gate106inter4));
  nand2 gate678(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate679(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate680(.a(G364), .O(gate106inter7));
  inv1  gate681(.a(G365), .O(gate106inter8));
  nand2 gate682(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate683(.a(s_19), .b(gate106inter3), .O(gate106inter10));
  nor2  gate684(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate685(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate686(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate925(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate926(.a(gate108inter0), .b(s_54), .O(gate108inter1));
  and2  gate927(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate928(.a(s_54), .O(gate108inter3));
  inv1  gate929(.a(s_55), .O(gate108inter4));
  nand2 gate930(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate931(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate932(.a(G368), .O(gate108inter7));
  inv1  gate933(.a(G369), .O(gate108inter8));
  nand2 gate934(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate935(.a(s_55), .b(gate108inter3), .O(gate108inter10));
  nor2  gate936(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate937(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate938(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate743(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate744(.a(gate114inter0), .b(s_28), .O(gate114inter1));
  and2  gate745(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate746(.a(s_28), .O(gate114inter3));
  inv1  gate747(.a(s_29), .O(gate114inter4));
  nand2 gate748(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate749(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate750(.a(G380), .O(gate114inter7));
  inv1  gate751(.a(G381), .O(gate114inter8));
  nand2 gate752(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate753(.a(s_29), .b(gate114inter3), .O(gate114inter10));
  nor2  gate754(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate755(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate756(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1583(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1584(.a(gate117inter0), .b(s_148), .O(gate117inter1));
  and2  gate1585(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1586(.a(s_148), .O(gate117inter3));
  inv1  gate1587(.a(s_149), .O(gate117inter4));
  nand2 gate1588(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1589(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1590(.a(G386), .O(gate117inter7));
  inv1  gate1591(.a(G387), .O(gate117inter8));
  nand2 gate1592(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1593(.a(s_149), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1594(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1595(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1596(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate1275(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1276(.a(gate118inter0), .b(s_104), .O(gate118inter1));
  and2  gate1277(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1278(.a(s_104), .O(gate118inter3));
  inv1  gate1279(.a(s_105), .O(gate118inter4));
  nand2 gate1280(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1281(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1282(.a(G388), .O(gate118inter7));
  inv1  gate1283(.a(G389), .O(gate118inter8));
  nand2 gate1284(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1285(.a(s_105), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1286(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1287(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1288(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1751(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1752(.a(gate119inter0), .b(s_172), .O(gate119inter1));
  and2  gate1753(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1754(.a(s_172), .O(gate119inter3));
  inv1  gate1755(.a(s_173), .O(gate119inter4));
  nand2 gate1756(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1757(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1758(.a(G390), .O(gate119inter7));
  inv1  gate1759(.a(G391), .O(gate119inter8));
  nand2 gate1760(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1761(.a(s_173), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1762(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1763(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1764(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate827(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate828(.a(gate120inter0), .b(s_40), .O(gate120inter1));
  and2  gate829(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate830(.a(s_40), .O(gate120inter3));
  inv1  gate831(.a(s_41), .O(gate120inter4));
  nand2 gate832(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate833(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate834(.a(G392), .O(gate120inter7));
  inv1  gate835(.a(G393), .O(gate120inter8));
  nand2 gate836(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate837(.a(s_41), .b(gate120inter3), .O(gate120inter10));
  nor2  gate838(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate839(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate840(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1695(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1696(.a(gate137inter0), .b(s_164), .O(gate137inter1));
  and2  gate1697(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1698(.a(s_164), .O(gate137inter3));
  inv1  gate1699(.a(s_165), .O(gate137inter4));
  nand2 gate1700(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1701(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1702(.a(G426), .O(gate137inter7));
  inv1  gate1703(.a(G429), .O(gate137inter8));
  nand2 gate1704(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1705(.a(s_165), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1706(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1707(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1708(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1331(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1332(.a(gate138inter0), .b(s_112), .O(gate138inter1));
  and2  gate1333(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1334(.a(s_112), .O(gate138inter3));
  inv1  gate1335(.a(s_113), .O(gate138inter4));
  nand2 gate1336(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1337(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1338(.a(G432), .O(gate138inter7));
  inv1  gate1339(.a(G435), .O(gate138inter8));
  nand2 gate1340(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1341(.a(s_113), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1342(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1343(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1344(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate561(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate562(.a(gate145inter0), .b(s_2), .O(gate145inter1));
  and2  gate563(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate564(.a(s_2), .O(gate145inter3));
  inv1  gate565(.a(s_3), .O(gate145inter4));
  nand2 gate566(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate567(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate568(.a(G474), .O(gate145inter7));
  inv1  gate569(.a(G477), .O(gate145inter8));
  nand2 gate570(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate571(.a(s_3), .b(gate145inter3), .O(gate145inter10));
  nor2  gate572(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate573(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate574(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1723(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1724(.a(gate148inter0), .b(s_168), .O(gate148inter1));
  and2  gate1725(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1726(.a(s_168), .O(gate148inter3));
  inv1  gate1727(.a(s_169), .O(gate148inter4));
  nand2 gate1728(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1729(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1730(.a(G492), .O(gate148inter7));
  inv1  gate1731(.a(G495), .O(gate148inter8));
  nand2 gate1732(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1733(.a(s_169), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1734(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1735(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1736(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1499(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1500(.a(gate150inter0), .b(s_136), .O(gate150inter1));
  and2  gate1501(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1502(.a(s_136), .O(gate150inter3));
  inv1  gate1503(.a(s_137), .O(gate150inter4));
  nand2 gate1504(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1505(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1506(.a(G504), .O(gate150inter7));
  inv1  gate1507(.a(G507), .O(gate150inter8));
  nand2 gate1508(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1509(.a(s_137), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1510(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1511(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1512(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1247(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1248(.a(gate151inter0), .b(s_100), .O(gate151inter1));
  and2  gate1249(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1250(.a(s_100), .O(gate151inter3));
  inv1  gate1251(.a(s_101), .O(gate151inter4));
  nand2 gate1252(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1253(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1254(.a(G510), .O(gate151inter7));
  inv1  gate1255(.a(G513), .O(gate151inter8));
  nand2 gate1256(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1257(.a(s_101), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1258(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1259(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1260(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1289(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1290(.a(gate163inter0), .b(s_106), .O(gate163inter1));
  and2  gate1291(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1292(.a(s_106), .O(gate163inter3));
  inv1  gate1293(.a(s_107), .O(gate163inter4));
  nand2 gate1294(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1295(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1296(.a(G456), .O(gate163inter7));
  inv1  gate1297(.a(G537), .O(gate163inter8));
  nand2 gate1298(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1299(.a(s_107), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1300(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1301(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1302(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1233(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1234(.a(gate169inter0), .b(s_98), .O(gate169inter1));
  and2  gate1235(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1236(.a(s_98), .O(gate169inter3));
  inv1  gate1237(.a(s_99), .O(gate169inter4));
  nand2 gate1238(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1239(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1240(.a(G474), .O(gate169inter7));
  inv1  gate1241(.a(G546), .O(gate169inter8));
  nand2 gate1242(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1243(.a(s_99), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1244(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1245(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1246(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1877(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1878(.a(gate171inter0), .b(s_190), .O(gate171inter1));
  and2  gate1879(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1880(.a(s_190), .O(gate171inter3));
  inv1  gate1881(.a(s_191), .O(gate171inter4));
  nand2 gate1882(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1883(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1884(.a(G480), .O(gate171inter7));
  inv1  gate1885(.a(G549), .O(gate171inter8));
  nand2 gate1886(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1887(.a(s_191), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1888(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1889(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1890(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1611(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1612(.a(gate174inter0), .b(s_152), .O(gate174inter1));
  and2  gate1613(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1614(.a(s_152), .O(gate174inter3));
  inv1  gate1615(.a(s_153), .O(gate174inter4));
  nand2 gate1616(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1617(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1618(.a(G489), .O(gate174inter7));
  inv1  gate1619(.a(G552), .O(gate174inter8));
  nand2 gate1620(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1621(.a(s_153), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1622(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1623(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1624(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1597(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1598(.a(gate178inter0), .b(s_150), .O(gate178inter1));
  and2  gate1599(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1600(.a(s_150), .O(gate178inter3));
  inv1  gate1601(.a(s_151), .O(gate178inter4));
  nand2 gate1602(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1603(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1604(.a(G501), .O(gate178inter7));
  inv1  gate1605(.a(G558), .O(gate178inter8));
  nand2 gate1606(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1607(.a(s_151), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1608(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1609(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1610(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate757(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate758(.a(gate180inter0), .b(s_30), .O(gate180inter1));
  and2  gate759(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate760(.a(s_30), .O(gate180inter3));
  inv1  gate761(.a(s_31), .O(gate180inter4));
  nand2 gate762(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate763(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate764(.a(G507), .O(gate180inter7));
  inv1  gate765(.a(G561), .O(gate180inter8));
  nand2 gate766(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate767(.a(s_31), .b(gate180inter3), .O(gate180inter10));
  nor2  gate768(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate769(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate770(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1359(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1360(.a(gate187inter0), .b(s_116), .O(gate187inter1));
  and2  gate1361(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1362(.a(s_116), .O(gate187inter3));
  inv1  gate1363(.a(s_117), .O(gate187inter4));
  nand2 gate1364(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1365(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1366(.a(G574), .O(gate187inter7));
  inv1  gate1367(.a(G575), .O(gate187inter8));
  nand2 gate1368(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1369(.a(s_117), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1370(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1371(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1372(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate855(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate856(.a(gate188inter0), .b(s_44), .O(gate188inter1));
  and2  gate857(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate858(.a(s_44), .O(gate188inter3));
  inv1  gate859(.a(s_45), .O(gate188inter4));
  nand2 gate860(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate861(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate862(.a(G576), .O(gate188inter7));
  inv1  gate863(.a(G577), .O(gate188inter8));
  nand2 gate864(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate865(.a(s_45), .b(gate188inter3), .O(gate188inter10));
  nor2  gate866(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate867(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate868(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1555(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1556(.a(gate190inter0), .b(s_144), .O(gate190inter1));
  and2  gate1557(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1558(.a(s_144), .O(gate190inter3));
  inv1  gate1559(.a(s_145), .O(gate190inter4));
  nand2 gate1560(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1561(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1562(.a(G580), .O(gate190inter7));
  inv1  gate1563(.a(G581), .O(gate190inter8));
  nand2 gate1564(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1565(.a(s_145), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1566(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1567(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1568(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate659(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate660(.a(gate194inter0), .b(s_16), .O(gate194inter1));
  and2  gate661(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate662(.a(s_16), .O(gate194inter3));
  inv1  gate663(.a(s_17), .O(gate194inter4));
  nand2 gate664(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate665(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate666(.a(G588), .O(gate194inter7));
  inv1  gate667(.a(G589), .O(gate194inter8));
  nand2 gate668(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate669(.a(s_17), .b(gate194inter3), .O(gate194inter10));
  nor2  gate670(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate671(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate672(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate883(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate884(.a(gate195inter0), .b(s_48), .O(gate195inter1));
  and2  gate885(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate886(.a(s_48), .O(gate195inter3));
  inv1  gate887(.a(s_49), .O(gate195inter4));
  nand2 gate888(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate889(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate890(.a(G590), .O(gate195inter7));
  inv1  gate891(.a(G591), .O(gate195inter8));
  nand2 gate892(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate893(.a(s_49), .b(gate195inter3), .O(gate195inter10));
  nor2  gate894(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate895(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate896(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1387(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1388(.a(gate196inter0), .b(s_120), .O(gate196inter1));
  and2  gate1389(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1390(.a(s_120), .O(gate196inter3));
  inv1  gate1391(.a(s_121), .O(gate196inter4));
  nand2 gate1392(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1393(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1394(.a(G592), .O(gate196inter7));
  inv1  gate1395(.a(G593), .O(gate196inter8));
  nand2 gate1396(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1397(.a(s_121), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1398(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1399(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1400(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1919(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1920(.a(gate204inter0), .b(s_196), .O(gate204inter1));
  and2  gate1921(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1922(.a(s_196), .O(gate204inter3));
  inv1  gate1923(.a(s_197), .O(gate204inter4));
  nand2 gate1924(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1925(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1926(.a(G607), .O(gate204inter7));
  inv1  gate1927(.a(G617), .O(gate204inter8));
  nand2 gate1928(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1929(.a(s_197), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1930(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1931(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1932(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate953(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate954(.a(gate208inter0), .b(s_58), .O(gate208inter1));
  and2  gate955(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate956(.a(s_58), .O(gate208inter3));
  inv1  gate957(.a(s_59), .O(gate208inter4));
  nand2 gate958(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate959(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate960(.a(G627), .O(gate208inter7));
  inv1  gate961(.a(G637), .O(gate208inter8));
  nand2 gate962(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate963(.a(s_59), .b(gate208inter3), .O(gate208inter10));
  nor2  gate964(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate965(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate966(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate967(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate968(.a(gate218inter0), .b(s_60), .O(gate218inter1));
  and2  gate969(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate970(.a(s_60), .O(gate218inter3));
  inv1  gate971(.a(s_61), .O(gate218inter4));
  nand2 gate972(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate973(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate974(.a(G627), .O(gate218inter7));
  inv1  gate975(.a(G678), .O(gate218inter8));
  nand2 gate976(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate977(.a(s_61), .b(gate218inter3), .O(gate218inter10));
  nor2  gate978(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate979(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate980(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1891(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1892(.a(gate225inter0), .b(s_192), .O(gate225inter1));
  and2  gate1893(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1894(.a(s_192), .O(gate225inter3));
  inv1  gate1895(.a(s_193), .O(gate225inter4));
  nand2 gate1896(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1897(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1898(.a(G690), .O(gate225inter7));
  inv1  gate1899(.a(G691), .O(gate225inter8));
  nand2 gate1900(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1901(.a(s_193), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1902(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1903(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1904(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate729(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate730(.a(gate226inter0), .b(s_26), .O(gate226inter1));
  and2  gate731(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate732(.a(s_26), .O(gate226inter3));
  inv1  gate733(.a(s_27), .O(gate226inter4));
  nand2 gate734(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate735(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate736(.a(G692), .O(gate226inter7));
  inv1  gate737(.a(G693), .O(gate226inter8));
  nand2 gate738(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate739(.a(s_27), .b(gate226inter3), .O(gate226inter10));
  nor2  gate740(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate741(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate742(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1527(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1528(.a(gate228inter0), .b(s_140), .O(gate228inter1));
  and2  gate1529(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1530(.a(s_140), .O(gate228inter3));
  inv1  gate1531(.a(s_141), .O(gate228inter4));
  nand2 gate1532(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1533(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1534(.a(G696), .O(gate228inter7));
  inv1  gate1535(.a(G697), .O(gate228inter8));
  nand2 gate1536(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1537(.a(s_141), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1538(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1539(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1540(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate869(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate870(.a(gate237inter0), .b(s_46), .O(gate237inter1));
  and2  gate871(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate872(.a(s_46), .O(gate237inter3));
  inv1  gate873(.a(s_47), .O(gate237inter4));
  nand2 gate874(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate875(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate876(.a(G254), .O(gate237inter7));
  inv1  gate877(.a(G706), .O(gate237inter8));
  nand2 gate878(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate879(.a(s_47), .b(gate237inter3), .O(gate237inter10));
  nor2  gate880(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate881(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate882(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1415(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1416(.a(gate238inter0), .b(s_124), .O(gate238inter1));
  and2  gate1417(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1418(.a(s_124), .O(gate238inter3));
  inv1  gate1419(.a(s_125), .O(gate238inter4));
  nand2 gate1420(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1421(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1422(.a(G257), .O(gate238inter7));
  inv1  gate1423(.a(G709), .O(gate238inter8));
  nand2 gate1424(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1425(.a(s_125), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1426(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1427(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1428(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate911(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate912(.a(gate243inter0), .b(s_52), .O(gate243inter1));
  and2  gate913(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate914(.a(s_52), .O(gate243inter3));
  inv1  gate915(.a(s_53), .O(gate243inter4));
  nand2 gate916(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate917(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate918(.a(G245), .O(gate243inter7));
  inv1  gate919(.a(G733), .O(gate243inter8));
  nand2 gate920(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate921(.a(s_53), .b(gate243inter3), .O(gate243inter10));
  nor2  gate922(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate923(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate924(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1401(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1402(.a(gate249inter0), .b(s_122), .O(gate249inter1));
  and2  gate1403(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1404(.a(s_122), .O(gate249inter3));
  inv1  gate1405(.a(s_123), .O(gate249inter4));
  nand2 gate1406(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1407(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1408(.a(G254), .O(gate249inter7));
  inv1  gate1409(.a(G742), .O(gate249inter8));
  nand2 gate1410(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1411(.a(s_123), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1412(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1413(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1414(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1667(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1668(.a(gate250inter0), .b(s_160), .O(gate250inter1));
  and2  gate1669(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1670(.a(s_160), .O(gate250inter3));
  inv1  gate1671(.a(s_161), .O(gate250inter4));
  nand2 gate1672(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1673(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1674(.a(G706), .O(gate250inter7));
  inv1  gate1675(.a(G742), .O(gate250inter8));
  nand2 gate1676(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1677(.a(s_161), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1678(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1679(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1680(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1219(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1220(.a(gate252inter0), .b(s_96), .O(gate252inter1));
  and2  gate1221(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1222(.a(s_96), .O(gate252inter3));
  inv1  gate1223(.a(s_97), .O(gate252inter4));
  nand2 gate1224(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1225(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1226(.a(G709), .O(gate252inter7));
  inv1  gate1227(.a(G745), .O(gate252inter8));
  nand2 gate1228(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1229(.a(s_97), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1230(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1231(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1232(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1303(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1304(.a(gate257inter0), .b(s_108), .O(gate257inter1));
  and2  gate1305(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1306(.a(s_108), .O(gate257inter3));
  inv1  gate1307(.a(s_109), .O(gate257inter4));
  nand2 gate1308(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1309(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1310(.a(G754), .O(gate257inter7));
  inv1  gate1311(.a(G755), .O(gate257inter8));
  nand2 gate1312(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1313(.a(s_109), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1314(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1315(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1316(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1485(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1486(.a(gate260inter0), .b(s_134), .O(gate260inter1));
  and2  gate1487(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1488(.a(s_134), .O(gate260inter3));
  inv1  gate1489(.a(s_135), .O(gate260inter4));
  nand2 gate1490(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1491(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1492(.a(G760), .O(gate260inter7));
  inv1  gate1493(.a(G761), .O(gate260inter8));
  nand2 gate1494(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1495(.a(s_135), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1496(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1497(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1498(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1821(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1822(.a(gate261inter0), .b(s_182), .O(gate261inter1));
  and2  gate1823(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1824(.a(s_182), .O(gate261inter3));
  inv1  gate1825(.a(s_183), .O(gate261inter4));
  nand2 gate1826(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1827(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1828(.a(G762), .O(gate261inter7));
  inv1  gate1829(.a(G763), .O(gate261inter8));
  nand2 gate1830(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1831(.a(s_183), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1832(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1833(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1834(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate589(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate590(.a(gate266inter0), .b(s_6), .O(gate266inter1));
  and2  gate591(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate592(.a(s_6), .O(gate266inter3));
  inv1  gate593(.a(s_7), .O(gate266inter4));
  nand2 gate594(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate595(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate596(.a(G645), .O(gate266inter7));
  inv1  gate597(.a(G773), .O(gate266inter8));
  nand2 gate598(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate599(.a(s_7), .b(gate266inter3), .O(gate266inter10));
  nor2  gate600(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate601(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate602(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate841(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate842(.a(gate267inter0), .b(s_42), .O(gate267inter1));
  and2  gate843(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate844(.a(s_42), .O(gate267inter3));
  inv1  gate845(.a(s_43), .O(gate267inter4));
  nand2 gate846(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate847(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate848(.a(G648), .O(gate267inter7));
  inv1  gate849(.a(G776), .O(gate267inter8));
  nand2 gate850(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate851(.a(s_43), .b(gate267inter3), .O(gate267inter10));
  nor2  gate852(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate853(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate854(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1205(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1206(.a(gate268inter0), .b(s_94), .O(gate268inter1));
  and2  gate1207(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1208(.a(s_94), .O(gate268inter3));
  inv1  gate1209(.a(s_95), .O(gate268inter4));
  nand2 gate1210(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1211(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1212(.a(G651), .O(gate268inter7));
  inv1  gate1213(.a(G779), .O(gate268inter8));
  nand2 gate1214(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1215(.a(s_95), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1216(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1217(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1218(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1569(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1570(.a(gate270inter0), .b(s_146), .O(gate270inter1));
  and2  gate1571(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1572(.a(s_146), .O(gate270inter3));
  inv1  gate1573(.a(s_147), .O(gate270inter4));
  nand2 gate1574(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1575(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1576(.a(G657), .O(gate270inter7));
  inv1  gate1577(.a(G785), .O(gate270inter8));
  nand2 gate1578(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1579(.a(s_147), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1580(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1581(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1582(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate603(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate604(.a(gate278inter0), .b(s_8), .O(gate278inter1));
  and2  gate605(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate606(.a(s_8), .O(gate278inter3));
  inv1  gate607(.a(s_9), .O(gate278inter4));
  nand2 gate608(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate609(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate610(.a(G776), .O(gate278inter7));
  inv1  gate611(.a(G800), .O(gate278inter8));
  nand2 gate612(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate613(.a(s_9), .b(gate278inter3), .O(gate278inter10));
  nor2  gate614(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate615(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate616(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1051(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1052(.a(gate281inter0), .b(s_72), .O(gate281inter1));
  and2  gate1053(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1054(.a(s_72), .O(gate281inter3));
  inv1  gate1055(.a(s_73), .O(gate281inter4));
  nand2 gate1056(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1057(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1058(.a(G654), .O(gate281inter7));
  inv1  gate1059(.a(G806), .O(gate281inter8));
  nand2 gate1060(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1061(.a(s_73), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1062(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1063(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1064(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate785(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate786(.a(gate282inter0), .b(s_34), .O(gate282inter1));
  and2  gate787(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate788(.a(s_34), .O(gate282inter3));
  inv1  gate789(.a(s_35), .O(gate282inter4));
  nand2 gate790(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate791(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate792(.a(G782), .O(gate282inter7));
  inv1  gate793(.a(G806), .O(gate282inter8));
  nand2 gate794(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate795(.a(s_35), .b(gate282inter3), .O(gate282inter10));
  nor2  gate796(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate797(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate798(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1191(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1192(.a(gate283inter0), .b(s_92), .O(gate283inter1));
  and2  gate1193(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1194(.a(s_92), .O(gate283inter3));
  inv1  gate1195(.a(s_93), .O(gate283inter4));
  nand2 gate1196(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1197(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1198(.a(G657), .O(gate283inter7));
  inv1  gate1199(.a(G809), .O(gate283inter8));
  nand2 gate1200(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1201(.a(s_93), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1202(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1203(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1204(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1443(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1444(.a(gate289inter0), .b(s_128), .O(gate289inter1));
  and2  gate1445(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1446(.a(s_128), .O(gate289inter3));
  inv1  gate1447(.a(s_129), .O(gate289inter4));
  nand2 gate1448(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1449(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1450(.a(G818), .O(gate289inter7));
  inv1  gate1451(.a(G819), .O(gate289inter8));
  nand2 gate1452(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1453(.a(s_129), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1454(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1455(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1456(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1065(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1066(.a(gate391inter0), .b(s_74), .O(gate391inter1));
  and2  gate1067(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1068(.a(s_74), .O(gate391inter3));
  inv1  gate1069(.a(s_75), .O(gate391inter4));
  nand2 gate1070(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1071(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1072(.a(G5), .O(gate391inter7));
  inv1  gate1073(.a(G1048), .O(gate391inter8));
  nand2 gate1074(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1075(.a(s_75), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1076(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1077(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1078(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1093(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1094(.a(gate395inter0), .b(s_78), .O(gate395inter1));
  and2  gate1095(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1096(.a(s_78), .O(gate395inter3));
  inv1  gate1097(.a(s_79), .O(gate395inter4));
  nand2 gate1098(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1099(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1100(.a(G9), .O(gate395inter7));
  inv1  gate1101(.a(G1060), .O(gate395inter8));
  nand2 gate1102(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1103(.a(s_79), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1104(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1105(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1106(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1947(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1948(.a(gate402inter0), .b(s_200), .O(gate402inter1));
  and2  gate1949(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1950(.a(s_200), .O(gate402inter3));
  inv1  gate1951(.a(s_201), .O(gate402inter4));
  nand2 gate1952(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1953(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1954(.a(G16), .O(gate402inter7));
  inv1  gate1955(.a(G1081), .O(gate402inter8));
  nand2 gate1956(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1957(.a(s_201), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1958(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1959(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1960(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1639(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1640(.a(gate410inter0), .b(s_156), .O(gate410inter1));
  and2  gate1641(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1642(.a(s_156), .O(gate410inter3));
  inv1  gate1643(.a(s_157), .O(gate410inter4));
  nand2 gate1644(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1645(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1646(.a(G24), .O(gate410inter7));
  inv1  gate1647(.a(G1105), .O(gate410inter8));
  nand2 gate1648(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1649(.a(s_157), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1650(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1651(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1652(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1009(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1010(.a(gate411inter0), .b(s_66), .O(gate411inter1));
  and2  gate1011(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1012(.a(s_66), .O(gate411inter3));
  inv1  gate1013(.a(s_67), .O(gate411inter4));
  nand2 gate1014(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1015(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1016(.a(G25), .O(gate411inter7));
  inv1  gate1017(.a(G1108), .O(gate411inter8));
  nand2 gate1018(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1019(.a(s_67), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1020(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1021(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1022(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1681(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1682(.a(gate413inter0), .b(s_162), .O(gate413inter1));
  and2  gate1683(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1684(.a(s_162), .O(gate413inter3));
  inv1  gate1685(.a(s_163), .O(gate413inter4));
  nand2 gate1686(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1687(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1688(.a(G27), .O(gate413inter7));
  inv1  gate1689(.a(G1114), .O(gate413inter8));
  nand2 gate1690(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1691(.a(s_163), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1692(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1693(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1694(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1037(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1038(.a(gate416inter0), .b(s_70), .O(gate416inter1));
  and2  gate1039(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1040(.a(s_70), .O(gate416inter3));
  inv1  gate1041(.a(s_71), .O(gate416inter4));
  nand2 gate1042(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1043(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1044(.a(G30), .O(gate416inter7));
  inv1  gate1045(.a(G1123), .O(gate416inter8));
  nand2 gate1046(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1047(.a(s_71), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1048(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1049(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1050(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1513(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1514(.a(gate421inter0), .b(s_138), .O(gate421inter1));
  and2  gate1515(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1516(.a(s_138), .O(gate421inter3));
  inv1  gate1517(.a(s_139), .O(gate421inter4));
  nand2 gate1518(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1519(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1520(.a(G2), .O(gate421inter7));
  inv1  gate1521(.a(G1135), .O(gate421inter8));
  nand2 gate1522(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1523(.a(s_139), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1524(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1525(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1526(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1457(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1458(.a(gate435inter0), .b(s_130), .O(gate435inter1));
  and2  gate1459(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1460(.a(s_130), .O(gate435inter3));
  inv1  gate1461(.a(s_131), .O(gate435inter4));
  nand2 gate1462(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1463(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1464(.a(G9), .O(gate435inter7));
  inv1  gate1465(.a(G1156), .O(gate435inter8));
  nand2 gate1466(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1467(.a(s_131), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1468(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1469(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1470(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1905(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1906(.a(gate437inter0), .b(s_194), .O(gate437inter1));
  and2  gate1907(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1908(.a(s_194), .O(gate437inter3));
  inv1  gate1909(.a(s_195), .O(gate437inter4));
  nand2 gate1910(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1911(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1912(.a(G10), .O(gate437inter7));
  inv1  gate1913(.a(G1159), .O(gate437inter8));
  nand2 gate1914(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1915(.a(s_195), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1916(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1917(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1918(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate575(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate576(.a(gate440inter0), .b(s_4), .O(gate440inter1));
  and2  gate577(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate578(.a(s_4), .O(gate440inter3));
  inv1  gate579(.a(s_5), .O(gate440inter4));
  nand2 gate580(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate581(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate582(.a(G1066), .O(gate440inter7));
  inv1  gate583(.a(G1162), .O(gate440inter8));
  nand2 gate584(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate585(.a(s_5), .b(gate440inter3), .O(gate440inter10));
  nor2  gate586(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate587(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate588(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate939(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate940(.a(gate442inter0), .b(s_56), .O(gate442inter1));
  and2  gate941(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate942(.a(s_56), .O(gate442inter3));
  inv1  gate943(.a(s_57), .O(gate442inter4));
  nand2 gate944(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate945(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate946(.a(G1069), .O(gate442inter7));
  inv1  gate947(.a(G1165), .O(gate442inter8));
  nand2 gate948(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate949(.a(s_57), .b(gate442inter3), .O(gate442inter10));
  nor2  gate950(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate951(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate952(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1779(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1780(.a(gate444inter0), .b(s_176), .O(gate444inter1));
  and2  gate1781(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1782(.a(s_176), .O(gate444inter3));
  inv1  gate1783(.a(s_177), .O(gate444inter4));
  nand2 gate1784(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1785(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1786(.a(G1072), .O(gate444inter7));
  inv1  gate1787(.a(G1168), .O(gate444inter8));
  nand2 gate1788(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1789(.a(s_177), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1790(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1791(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1792(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1849(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1850(.a(gate446inter0), .b(s_186), .O(gate446inter1));
  and2  gate1851(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1852(.a(s_186), .O(gate446inter3));
  inv1  gate1853(.a(s_187), .O(gate446inter4));
  nand2 gate1854(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1855(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1856(.a(G1075), .O(gate446inter7));
  inv1  gate1857(.a(G1171), .O(gate446inter8));
  nand2 gate1858(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1859(.a(s_187), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1860(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1861(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1862(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1807(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1808(.a(gate448inter0), .b(s_180), .O(gate448inter1));
  and2  gate1809(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1810(.a(s_180), .O(gate448inter3));
  inv1  gate1811(.a(s_181), .O(gate448inter4));
  nand2 gate1812(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1813(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1814(.a(G1078), .O(gate448inter7));
  inv1  gate1815(.a(G1174), .O(gate448inter8));
  nand2 gate1816(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1817(.a(s_181), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1818(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1819(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1820(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate771(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate772(.a(gate449inter0), .b(s_32), .O(gate449inter1));
  and2  gate773(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate774(.a(s_32), .O(gate449inter3));
  inv1  gate775(.a(s_33), .O(gate449inter4));
  nand2 gate776(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate777(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate778(.a(G16), .O(gate449inter7));
  inv1  gate779(.a(G1177), .O(gate449inter8));
  nand2 gate780(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate781(.a(s_33), .b(gate449inter3), .O(gate449inter10));
  nor2  gate782(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate783(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate784(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1079(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1080(.a(gate452inter0), .b(s_76), .O(gate452inter1));
  and2  gate1081(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1082(.a(s_76), .O(gate452inter3));
  inv1  gate1083(.a(s_77), .O(gate452inter4));
  nand2 gate1084(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1085(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1086(.a(G1084), .O(gate452inter7));
  inv1  gate1087(.a(G1180), .O(gate452inter8));
  nand2 gate1088(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1089(.a(s_77), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1090(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1091(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1092(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1107(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1108(.a(gate462inter0), .b(s_80), .O(gate462inter1));
  and2  gate1109(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1110(.a(s_80), .O(gate462inter3));
  inv1  gate1111(.a(s_81), .O(gate462inter4));
  nand2 gate1112(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1113(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1114(.a(G1099), .O(gate462inter7));
  inv1  gate1115(.a(G1195), .O(gate462inter8));
  nand2 gate1116(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1117(.a(s_81), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1118(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1119(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1120(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate687(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate688(.a(gate465inter0), .b(s_20), .O(gate465inter1));
  and2  gate689(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate690(.a(s_20), .O(gate465inter3));
  inv1  gate691(.a(s_21), .O(gate465inter4));
  nand2 gate692(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate693(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate694(.a(G24), .O(gate465inter7));
  inv1  gate695(.a(G1201), .O(gate465inter8));
  nand2 gate696(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate697(.a(s_21), .b(gate465inter3), .O(gate465inter10));
  nor2  gate698(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate699(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate700(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate981(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate982(.a(gate472inter0), .b(s_62), .O(gate472inter1));
  and2  gate983(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate984(.a(s_62), .O(gate472inter3));
  inv1  gate985(.a(s_63), .O(gate472inter4));
  nand2 gate986(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate987(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate988(.a(G1114), .O(gate472inter7));
  inv1  gate989(.a(G1210), .O(gate472inter8));
  nand2 gate990(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate991(.a(s_63), .b(gate472inter3), .O(gate472inter10));
  nor2  gate992(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate993(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate994(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1149(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1150(.a(gate473inter0), .b(s_86), .O(gate473inter1));
  and2  gate1151(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1152(.a(s_86), .O(gate473inter3));
  inv1  gate1153(.a(s_87), .O(gate473inter4));
  nand2 gate1154(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1155(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1156(.a(G28), .O(gate473inter7));
  inv1  gate1157(.a(G1213), .O(gate473inter8));
  nand2 gate1158(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1159(.a(s_87), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1160(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1161(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1162(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1933(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1934(.a(gate475inter0), .b(s_198), .O(gate475inter1));
  and2  gate1935(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1936(.a(s_198), .O(gate475inter3));
  inv1  gate1937(.a(s_199), .O(gate475inter4));
  nand2 gate1938(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1939(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1940(.a(G29), .O(gate475inter7));
  inv1  gate1941(.a(G1216), .O(gate475inter8));
  nand2 gate1942(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1943(.a(s_199), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1944(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1945(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1946(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1023(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1024(.a(gate477inter0), .b(s_68), .O(gate477inter1));
  and2  gate1025(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1026(.a(s_68), .O(gate477inter3));
  inv1  gate1027(.a(s_69), .O(gate477inter4));
  nand2 gate1028(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1029(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1030(.a(G30), .O(gate477inter7));
  inv1  gate1031(.a(G1219), .O(gate477inter8));
  nand2 gate1032(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1033(.a(s_69), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1034(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1035(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1036(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1317(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1318(.a(gate478inter0), .b(s_110), .O(gate478inter1));
  and2  gate1319(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1320(.a(s_110), .O(gate478inter3));
  inv1  gate1321(.a(s_111), .O(gate478inter4));
  nand2 gate1322(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1323(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1324(.a(G1123), .O(gate478inter7));
  inv1  gate1325(.a(G1219), .O(gate478inter8));
  nand2 gate1326(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1327(.a(s_111), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1328(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1329(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1330(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1261(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1262(.a(gate481inter0), .b(s_102), .O(gate481inter1));
  and2  gate1263(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1264(.a(s_102), .O(gate481inter3));
  inv1  gate1265(.a(s_103), .O(gate481inter4));
  nand2 gate1266(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1267(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1268(.a(G32), .O(gate481inter7));
  inv1  gate1269(.a(G1225), .O(gate481inter8));
  nand2 gate1270(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1271(.a(s_103), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1272(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1273(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1274(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1373(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1374(.a(gate482inter0), .b(s_118), .O(gate482inter1));
  and2  gate1375(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1376(.a(s_118), .O(gate482inter3));
  inv1  gate1377(.a(s_119), .O(gate482inter4));
  nand2 gate1378(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1379(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1380(.a(G1129), .O(gate482inter7));
  inv1  gate1381(.a(G1225), .O(gate482inter8));
  nand2 gate1382(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1383(.a(s_119), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1384(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1385(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1386(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate631(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate632(.a(gate483inter0), .b(s_12), .O(gate483inter1));
  and2  gate633(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate634(.a(s_12), .O(gate483inter3));
  inv1  gate635(.a(s_13), .O(gate483inter4));
  nand2 gate636(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate637(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate638(.a(G1228), .O(gate483inter7));
  inv1  gate639(.a(G1229), .O(gate483inter8));
  nand2 gate640(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate641(.a(s_13), .b(gate483inter3), .O(gate483inter10));
  nor2  gate642(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate643(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate644(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1793(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1794(.a(gate492inter0), .b(s_178), .O(gate492inter1));
  and2  gate1795(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1796(.a(s_178), .O(gate492inter3));
  inv1  gate1797(.a(s_179), .O(gate492inter4));
  nand2 gate1798(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1799(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1800(.a(G1246), .O(gate492inter7));
  inv1  gate1801(.a(G1247), .O(gate492inter8));
  nand2 gate1802(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1803(.a(s_179), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1804(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1805(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1806(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1737(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1738(.a(gate493inter0), .b(s_170), .O(gate493inter1));
  and2  gate1739(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1740(.a(s_170), .O(gate493inter3));
  inv1  gate1741(.a(s_171), .O(gate493inter4));
  nand2 gate1742(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1743(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1744(.a(G1248), .O(gate493inter7));
  inv1  gate1745(.a(G1249), .O(gate493inter8));
  nand2 gate1746(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1747(.a(s_171), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1748(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1749(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1750(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1121(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1122(.a(gate501inter0), .b(s_82), .O(gate501inter1));
  and2  gate1123(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1124(.a(s_82), .O(gate501inter3));
  inv1  gate1125(.a(s_83), .O(gate501inter4));
  nand2 gate1126(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1127(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1128(.a(G1264), .O(gate501inter7));
  inv1  gate1129(.a(G1265), .O(gate501inter8));
  nand2 gate1130(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1131(.a(s_83), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1132(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1133(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1134(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule