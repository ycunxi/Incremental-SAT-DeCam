module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
input s_382,s_383;//RE__ALLOW(00,01,10,11);
input s_384,s_385;//RE__ALLOW(00,01,10,11);
input s_386,s_387;//RE__ALLOW(00,01,10,11);
input s_388,s_389;//RE__ALLOW(00,01,10,11);
input s_390,s_391;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate729(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate730(.a(gate9inter0), .b(s_26), .O(gate9inter1));
  and2  gate731(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate732(.a(s_26), .O(gate9inter3));
  inv1  gate733(.a(s_27), .O(gate9inter4));
  nand2 gate734(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate735(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate736(.a(G1), .O(gate9inter7));
  inv1  gate737(.a(G2), .O(gate9inter8));
  nand2 gate738(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate739(.a(s_27), .b(gate9inter3), .O(gate9inter10));
  nor2  gate740(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate741(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate742(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1051(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1052(.a(gate16inter0), .b(s_72), .O(gate16inter1));
  and2  gate1053(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1054(.a(s_72), .O(gate16inter3));
  inv1  gate1055(.a(s_73), .O(gate16inter4));
  nand2 gate1056(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1057(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1058(.a(G15), .O(gate16inter7));
  inv1  gate1059(.a(G16), .O(gate16inter8));
  nand2 gate1060(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1061(.a(s_73), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1062(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1063(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1064(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2479(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2480(.a(gate18inter0), .b(s_276), .O(gate18inter1));
  and2  gate2481(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2482(.a(s_276), .O(gate18inter3));
  inv1  gate2483(.a(s_277), .O(gate18inter4));
  nand2 gate2484(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2485(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2486(.a(G19), .O(gate18inter7));
  inv1  gate2487(.a(G20), .O(gate18inter8));
  nand2 gate2488(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2489(.a(s_277), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2490(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2491(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2492(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1415(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1416(.a(gate19inter0), .b(s_124), .O(gate19inter1));
  and2  gate1417(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1418(.a(s_124), .O(gate19inter3));
  inv1  gate1419(.a(s_125), .O(gate19inter4));
  nand2 gate1420(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1421(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1422(.a(G21), .O(gate19inter7));
  inv1  gate1423(.a(G22), .O(gate19inter8));
  nand2 gate1424(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1425(.a(s_125), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1426(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1427(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1428(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate3235(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate3236(.a(gate21inter0), .b(s_384), .O(gate21inter1));
  and2  gate3237(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate3238(.a(s_384), .O(gate21inter3));
  inv1  gate3239(.a(s_385), .O(gate21inter4));
  nand2 gate3240(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate3241(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate3242(.a(G25), .O(gate21inter7));
  inv1  gate3243(.a(G26), .O(gate21inter8));
  nand2 gate3244(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate3245(.a(s_385), .b(gate21inter3), .O(gate21inter10));
  nor2  gate3246(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate3247(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate3248(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate589(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate590(.a(gate22inter0), .b(s_6), .O(gate22inter1));
  and2  gate591(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate592(.a(s_6), .O(gate22inter3));
  inv1  gate593(.a(s_7), .O(gate22inter4));
  nand2 gate594(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate595(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate596(.a(G27), .O(gate22inter7));
  inv1  gate597(.a(G28), .O(gate22inter8));
  nand2 gate598(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate599(.a(s_7), .b(gate22inter3), .O(gate22inter10));
  nor2  gate600(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate601(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate602(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1023(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1024(.a(gate23inter0), .b(s_68), .O(gate23inter1));
  and2  gate1025(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1026(.a(s_68), .O(gate23inter3));
  inv1  gate1027(.a(s_69), .O(gate23inter4));
  nand2 gate1028(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1029(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1030(.a(G29), .O(gate23inter7));
  inv1  gate1031(.a(G30), .O(gate23inter8));
  nand2 gate1032(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1033(.a(s_69), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1034(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1035(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1036(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1975(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1976(.a(gate27inter0), .b(s_204), .O(gate27inter1));
  and2  gate1977(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1978(.a(s_204), .O(gate27inter3));
  inv1  gate1979(.a(s_205), .O(gate27inter4));
  nand2 gate1980(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1981(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1982(.a(G2), .O(gate27inter7));
  inv1  gate1983(.a(G6), .O(gate27inter8));
  nand2 gate1984(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1985(.a(s_205), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1986(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1987(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1988(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2689(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2690(.a(gate29inter0), .b(s_306), .O(gate29inter1));
  and2  gate2691(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2692(.a(s_306), .O(gate29inter3));
  inv1  gate2693(.a(s_307), .O(gate29inter4));
  nand2 gate2694(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2695(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2696(.a(G3), .O(gate29inter7));
  inv1  gate2697(.a(G7), .O(gate29inter8));
  nand2 gate2698(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2699(.a(s_307), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2700(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2701(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2702(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate3053(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate3054(.a(gate30inter0), .b(s_358), .O(gate30inter1));
  and2  gate3055(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate3056(.a(s_358), .O(gate30inter3));
  inv1  gate3057(.a(s_359), .O(gate30inter4));
  nand2 gate3058(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate3059(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate3060(.a(G11), .O(gate30inter7));
  inv1  gate3061(.a(G15), .O(gate30inter8));
  nand2 gate3062(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate3063(.a(s_359), .b(gate30inter3), .O(gate30inter10));
  nor2  gate3064(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate3065(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate3066(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate3095(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate3096(.a(gate31inter0), .b(s_364), .O(gate31inter1));
  and2  gate3097(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate3098(.a(s_364), .O(gate31inter3));
  inv1  gate3099(.a(s_365), .O(gate31inter4));
  nand2 gate3100(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate3101(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate3102(.a(G4), .O(gate31inter7));
  inv1  gate3103(.a(G8), .O(gate31inter8));
  nand2 gate3104(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate3105(.a(s_365), .b(gate31inter3), .O(gate31inter10));
  nor2  gate3106(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate3107(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate3108(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1793(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1794(.a(gate33inter0), .b(s_178), .O(gate33inter1));
  and2  gate1795(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1796(.a(s_178), .O(gate33inter3));
  inv1  gate1797(.a(s_179), .O(gate33inter4));
  nand2 gate1798(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1799(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1800(.a(G17), .O(gate33inter7));
  inv1  gate1801(.a(G21), .O(gate33inter8));
  nand2 gate1802(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1803(.a(s_179), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1804(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1805(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1806(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2535(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2536(.a(gate34inter0), .b(s_284), .O(gate34inter1));
  and2  gate2537(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2538(.a(s_284), .O(gate34inter3));
  inv1  gate2539(.a(s_285), .O(gate34inter4));
  nand2 gate2540(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2541(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2542(.a(G25), .O(gate34inter7));
  inv1  gate2543(.a(G29), .O(gate34inter8));
  nand2 gate2544(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2545(.a(s_285), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2546(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2547(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2548(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate2815(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2816(.a(gate35inter0), .b(s_324), .O(gate35inter1));
  and2  gate2817(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2818(.a(s_324), .O(gate35inter3));
  inv1  gate2819(.a(s_325), .O(gate35inter4));
  nand2 gate2820(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2821(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2822(.a(G18), .O(gate35inter7));
  inv1  gate2823(.a(G22), .O(gate35inter8));
  nand2 gate2824(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2825(.a(s_325), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2826(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2827(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2828(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate3109(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate3110(.a(gate37inter0), .b(s_366), .O(gate37inter1));
  and2  gate3111(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate3112(.a(s_366), .O(gate37inter3));
  inv1  gate3113(.a(s_367), .O(gate37inter4));
  nand2 gate3114(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate3115(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate3116(.a(G19), .O(gate37inter7));
  inv1  gate3117(.a(G23), .O(gate37inter8));
  nand2 gate3118(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate3119(.a(s_367), .b(gate37inter3), .O(gate37inter10));
  nor2  gate3120(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate3121(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate3122(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2227(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2228(.a(gate38inter0), .b(s_240), .O(gate38inter1));
  and2  gate2229(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2230(.a(s_240), .O(gate38inter3));
  inv1  gate2231(.a(s_241), .O(gate38inter4));
  nand2 gate2232(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2233(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2234(.a(G27), .O(gate38inter7));
  inv1  gate2235(.a(G31), .O(gate38inter8));
  nand2 gate2236(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2237(.a(s_241), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2238(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2239(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2240(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate855(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate856(.a(gate40inter0), .b(s_44), .O(gate40inter1));
  and2  gate857(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate858(.a(s_44), .O(gate40inter3));
  inv1  gate859(.a(s_45), .O(gate40inter4));
  nand2 gate860(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate861(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate862(.a(G28), .O(gate40inter7));
  inv1  gate863(.a(G32), .O(gate40inter8));
  nand2 gate864(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate865(.a(s_45), .b(gate40inter3), .O(gate40inter10));
  nor2  gate866(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate867(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate868(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1821(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1822(.a(gate47inter0), .b(s_182), .O(gate47inter1));
  and2  gate1823(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1824(.a(s_182), .O(gate47inter3));
  inv1  gate1825(.a(s_183), .O(gate47inter4));
  nand2 gate1826(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1827(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1828(.a(G7), .O(gate47inter7));
  inv1  gate1829(.a(G275), .O(gate47inter8));
  nand2 gate1830(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1831(.a(s_183), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1832(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1833(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1834(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1163(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1164(.a(gate49inter0), .b(s_88), .O(gate49inter1));
  and2  gate1165(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1166(.a(s_88), .O(gate49inter3));
  inv1  gate1167(.a(s_89), .O(gate49inter4));
  nand2 gate1168(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1169(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1170(.a(G9), .O(gate49inter7));
  inv1  gate1171(.a(G278), .O(gate49inter8));
  nand2 gate1172(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1173(.a(s_89), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1174(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1175(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1176(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1919(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1920(.a(gate50inter0), .b(s_196), .O(gate50inter1));
  and2  gate1921(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1922(.a(s_196), .O(gate50inter3));
  inv1  gate1923(.a(s_197), .O(gate50inter4));
  nand2 gate1924(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1925(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1926(.a(G10), .O(gate50inter7));
  inv1  gate1927(.a(G278), .O(gate50inter8));
  nand2 gate1928(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1929(.a(s_197), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1930(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1931(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1932(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2969(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2970(.a(gate51inter0), .b(s_346), .O(gate51inter1));
  and2  gate2971(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2972(.a(s_346), .O(gate51inter3));
  inv1  gate2973(.a(s_347), .O(gate51inter4));
  nand2 gate2974(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2975(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2976(.a(G11), .O(gate51inter7));
  inv1  gate2977(.a(G281), .O(gate51inter8));
  nand2 gate2978(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2979(.a(s_347), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2980(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2981(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2982(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate3151(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate3152(.a(gate53inter0), .b(s_372), .O(gate53inter1));
  and2  gate3153(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate3154(.a(s_372), .O(gate53inter3));
  inv1  gate3155(.a(s_373), .O(gate53inter4));
  nand2 gate3156(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate3157(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate3158(.a(G13), .O(gate53inter7));
  inv1  gate3159(.a(G284), .O(gate53inter8));
  nand2 gate3160(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate3161(.a(s_373), .b(gate53inter3), .O(gate53inter10));
  nor2  gate3162(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate3163(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate3164(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1135(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1136(.a(gate57inter0), .b(s_84), .O(gate57inter1));
  and2  gate1137(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1138(.a(s_84), .O(gate57inter3));
  inv1  gate1139(.a(s_85), .O(gate57inter4));
  nand2 gate1140(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1141(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1142(.a(G17), .O(gate57inter7));
  inv1  gate1143(.a(G290), .O(gate57inter8));
  nand2 gate1144(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1145(.a(s_85), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1146(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1147(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1148(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1401(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1402(.a(gate58inter0), .b(s_122), .O(gate58inter1));
  and2  gate1403(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1404(.a(s_122), .O(gate58inter3));
  inv1  gate1405(.a(s_123), .O(gate58inter4));
  nand2 gate1406(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1407(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1408(.a(G18), .O(gate58inter7));
  inv1  gate1409(.a(G290), .O(gate58inter8));
  nand2 gate1410(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1411(.a(s_123), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1412(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1413(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1414(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate3277(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate3278(.a(gate59inter0), .b(s_390), .O(gate59inter1));
  and2  gate3279(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate3280(.a(s_390), .O(gate59inter3));
  inv1  gate3281(.a(s_391), .O(gate59inter4));
  nand2 gate3282(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate3283(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate3284(.a(G19), .O(gate59inter7));
  inv1  gate3285(.a(G293), .O(gate59inter8));
  nand2 gate3286(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate3287(.a(s_391), .b(gate59inter3), .O(gate59inter10));
  nor2  gate3288(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate3289(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate3290(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate3025(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate3026(.a(gate62inter0), .b(s_354), .O(gate62inter1));
  and2  gate3027(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate3028(.a(s_354), .O(gate62inter3));
  inv1  gate3029(.a(s_355), .O(gate62inter4));
  nand2 gate3030(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate3031(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate3032(.a(G22), .O(gate62inter7));
  inv1  gate3033(.a(G296), .O(gate62inter8));
  nand2 gate3034(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate3035(.a(s_355), .b(gate62inter3), .O(gate62inter10));
  nor2  gate3036(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate3037(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate3038(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1989(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1990(.a(gate63inter0), .b(s_206), .O(gate63inter1));
  and2  gate1991(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1992(.a(s_206), .O(gate63inter3));
  inv1  gate1993(.a(s_207), .O(gate63inter4));
  nand2 gate1994(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1995(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1996(.a(G23), .O(gate63inter7));
  inv1  gate1997(.a(G299), .O(gate63inter8));
  nand2 gate1998(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1999(.a(s_207), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2000(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2001(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2002(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate883(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate884(.a(gate66inter0), .b(s_48), .O(gate66inter1));
  and2  gate885(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate886(.a(s_48), .O(gate66inter3));
  inv1  gate887(.a(s_49), .O(gate66inter4));
  nand2 gate888(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate889(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate890(.a(G26), .O(gate66inter7));
  inv1  gate891(.a(G302), .O(gate66inter8));
  nand2 gate892(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate893(.a(s_49), .b(gate66inter3), .O(gate66inter10));
  nor2  gate894(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate895(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate896(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate561(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate562(.a(gate67inter0), .b(s_2), .O(gate67inter1));
  and2  gate563(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate564(.a(s_2), .O(gate67inter3));
  inv1  gate565(.a(s_3), .O(gate67inter4));
  nand2 gate566(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate567(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate568(.a(G27), .O(gate67inter7));
  inv1  gate569(.a(G305), .O(gate67inter8));
  nand2 gate570(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate571(.a(s_3), .b(gate67inter3), .O(gate67inter10));
  nor2  gate572(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate573(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate574(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate3263(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate3264(.a(gate68inter0), .b(s_388), .O(gate68inter1));
  and2  gate3265(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate3266(.a(s_388), .O(gate68inter3));
  inv1  gate3267(.a(s_389), .O(gate68inter4));
  nand2 gate3268(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate3269(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate3270(.a(G28), .O(gate68inter7));
  inv1  gate3271(.a(G305), .O(gate68inter8));
  nand2 gate3272(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate3273(.a(s_389), .b(gate68inter3), .O(gate68inter10));
  nor2  gate3274(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate3275(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate3276(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2787(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2788(.a(gate70inter0), .b(s_320), .O(gate70inter1));
  and2  gate2789(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2790(.a(s_320), .O(gate70inter3));
  inv1  gate2791(.a(s_321), .O(gate70inter4));
  nand2 gate2792(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2793(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2794(.a(G30), .O(gate70inter7));
  inv1  gate2795(.a(G308), .O(gate70inter8));
  nand2 gate2796(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2797(.a(s_321), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2798(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2799(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2800(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate575(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate576(.a(gate73inter0), .b(s_4), .O(gate73inter1));
  and2  gate577(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate578(.a(s_4), .O(gate73inter3));
  inv1  gate579(.a(s_5), .O(gate73inter4));
  nand2 gate580(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate581(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate582(.a(G1), .O(gate73inter7));
  inv1  gate583(.a(G314), .O(gate73inter8));
  nand2 gate584(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate585(.a(s_5), .b(gate73inter3), .O(gate73inter10));
  nor2  gate586(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate587(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate588(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate3067(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate3068(.a(gate74inter0), .b(s_360), .O(gate74inter1));
  and2  gate3069(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate3070(.a(s_360), .O(gate74inter3));
  inv1  gate3071(.a(s_361), .O(gate74inter4));
  nand2 gate3072(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate3073(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate3074(.a(G5), .O(gate74inter7));
  inv1  gate3075(.a(G314), .O(gate74inter8));
  nand2 gate3076(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate3077(.a(s_361), .b(gate74inter3), .O(gate74inter10));
  nor2  gate3078(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate3079(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate3080(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate2143(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2144(.a(gate75inter0), .b(s_228), .O(gate75inter1));
  and2  gate2145(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2146(.a(s_228), .O(gate75inter3));
  inv1  gate2147(.a(s_229), .O(gate75inter4));
  nand2 gate2148(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2149(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2150(.a(G9), .O(gate75inter7));
  inv1  gate2151(.a(G317), .O(gate75inter8));
  nand2 gate2152(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2153(.a(s_229), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2154(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2155(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2156(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2353(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2354(.a(gate80inter0), .b(s_258), .O(gate80inter1));
  and2  gate2355(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2356(.a(s_258), .O(gate80inter3));
  inv1  gate2357(.a(s_259), .O(gate80inter4));
  nand2 gate2358(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2359(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2360(.a(G14), .O(gate80inter7));
  inv1  gate2361(.a(G323), .O(gate80inter8));
  nand2 gate2362(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2363(.a(s_259), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2364(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2365(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2366(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1751(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1752(.a(gate81inter0), .b(s_172), .O(gate81inter1));
  and2  gate1753(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1754(.a(s_172), .O(gate81inter3));
  inv1  gate1755(.a(s_173), .O(gate81inter4));
  nand2 gate1756(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1757(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1758(.a(G3), .O(gate81inter7));
  inv1  gate1759(.a(G326), .O(gate81inter8));
  nand2 gate1760(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1761(.a(s_173), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1762(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1763(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1764(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1555(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1556(.a(gate82inter0), .b(s_144), .O(gate82inter1));
  and2  gate1557(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1558(.a(s_144), .O(gate82inter3));
  inv1  gate1559(.a(s_145), .O(gate82inter4));
  nand2 gate1560(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1561(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1562(.a(G7), .O(gate82inter7));
  inv1  gate1563(.a(G326), .O(gate82inter8));
  nand2 gate1564(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1565(.a(s_145), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1566(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1567(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1568(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate813(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate814(.a(gate85inter0), .b(s_38), .O(gate85inter1));
  and2  gate815(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate816(.a(s_38), .O(gate85inter3));
  inv1  gate817(.a(s_39), .O(gate85inter4));
  nand2 gate818(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate819(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate820(.a(G4), .O(gate85inter7));
  inv1  gate821(.a(G332), .O(gate85inter8));
  nand2 gate822(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate823(.a(s_39), .b(gate85inter3), .O(gate85inter10));
  nor2  gate824(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate825(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate826(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate743(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate744(.a(gate87inter0), .b(s_28), .O(gate87inter1));
  and2  gate745(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate746(.a(s_28), .O(gate87inter3));
  inv1  gate747(.a(s_29), .O(gate87inter4));
  nand2 gate748(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate749(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate750(.a(G12), .O(gate87inter7));
  inv1  gate751(.a(G335), .O(gate87inter8));
  nand2 gate752(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate753(.a(s_29), .b(gate87inter3), .O(gate87inter10));
  nor2  gate754(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate755(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate756(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate953(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate954(.a(gate91inter0), .b(s_58), .O(gate91inter1));
  and2  gate955(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate956(.a(s_58), .O(gate91inter3));
  inv1  gate957(.a(s_59), .O(gate91inter4));
  nand2 gate958(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate959(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate960(.a(G25), .O(gate91inter7));
  inv1  gate961(.a(G341), .O(gate91inter8));
  nand2 gate962(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate963(.a(s_59), .b(gate91inter3), .O(gate91inter10));
  nor2  gate964(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate965(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate966(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1443(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1444(.a(gate93inter0), .b(s_128), .O(gate93inter1));
  and2  gate1445(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1446(.a(s_128), .O(gate93inter3));
  inv1  gate1447(.a(s_129), .O(gate93inter4));
  nand2 gate1448(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1449(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1450(.a(G18), .O(gate93inter7));
  inv1  gate1451(.a(G344), .O(gate93inter8));
  nand2 gate1452(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1453(.a(s_129), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1454(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1455(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1456(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1009(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1010(.a(gate94inter0), .b(s_66), .O(gate94inter1));
  and2  gate1011(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1012(.a(s_66), .O(gate94inter3));
  inv1  gate1013(.a(s_67), .O(gate94inter4));
  nand2 gate1014(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1015(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1016(.a(G22), .O(gate94inter7));
  inv1  gate1017(.a(G344), .O(gate94inter8));
  nand2 gate1018(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1019(.a(s_67), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1020(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1021(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1022(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate939(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate940(.a(gate95inter0), .b(s_56), .O(gate95inter1));
  and2  gate941(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate942(.a(s_56), .O(gate95inter3));
  inv1  gate943(.a(s_57), .O(gate95inter4));
  nand2 gate944(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate945(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate946(.a(G26), .O(gate95inter7));
  inv1  gate947(.a(G347), .O(gate95inter8));
  nand2 gate948(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate949(.a(s_57), .b(gate95inter3), .O(gate95inter10));
  nor2  gate950(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate951(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate952(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2003(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2004(.a(gate96inter0), .b(s_208), .O(gate96inter1));
  and2  gate2005(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2006(.a(s_208), .O(gate96inter3));
  inv1  gate2007(.a(s_209), .O(gate96inter4));
  nand2 gate2008(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2009(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2010(.a(G30), .O(gate96inter7));
  inv1  gate2011(.a(G347), .O(gate96inter8));
  nand2 gate2012(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2013(.a(s_209), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2014(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2015(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2016(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2297(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2298(.a(gate97inter0), .b(s_250), .O(gate97inter1));
  and2  gate2299(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2300(.a(s_250), .O(gate97inter3));
  inv1  gate2301(.a(s_251), .O(gate97inter4));
  nand2 gate2302(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2303(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2304(.a(G19), .O(gate97inter7));
  inv1  gate2305(.a(G350), .O(gate97inter8));
  nand2 gate2306(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2307(.a(s_251), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2308(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2309(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2310(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1471(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1472(.a(gate99inter0), .b(s_132), .O(gate99inter1));
  and2  gate1473(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1474(.a(s_132), .O(gate99inter3));
  inv1  gate1475(.a(s_133), .O(gate99inter4));
  nand2 gate1476(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1477(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1478(.a(G27), .O(gate99inter7));
  inv1  gate1479(.a(G353), .O(gate99inter8));
  nand2 gate1480(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1481(.a(s_133), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1482(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1483(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1484(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate3207(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate3208(.a(gate100inter0), .b(s_380), .O(gate100inter1));
  and2  gate3209(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate3210(.a(s_380), .O(gate100inter3));
  inv1  gate3211(.a(s_381), .O(gate100inter4));
  nand2 gate3212(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate3213(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate3214(.a(G31), .O(gate100inter7));
  inv1  gate3215(.a(G353), .O(gate100inter8));
  nand2 gate3216(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate3217(.a(s_381), .b(gate100inter3), .O(gate100inter10));
  nor2  gate3218(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate3219(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate3220(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate3123(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate3124(.a(gate101inter0), .b(s_368), .O(gate101inter1));
  and2  gate3125(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate3126(.a(s_368), .O(gate101inter3));
  inv1  gate3127(.a(s_369), .O(gate101inter4));
  nand2 gate3128(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate3129(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate3130(.a(G20), .O(gate101inter7));
  inv1  gate3131(.a(G356), .O(gate101inter8));
  nand2 gate3132(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate3133(.a(s_369), .b(gate101inter3), .O(gate101inter10));
  nor2  gate3134(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate3135(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate3136(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate841(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate842(.a(gate103inter0), .b(s_42), .O(gate103inter1));
  and2  gate843(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate844(.a(s_42), .O(gate103inter3));
  inv1  gate845(.a(s_43), .O(gate103inter4));
  nand2 gate846(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate847(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate848(.a(G28), .O(gate103inter7));
  inv1  gate849(.a(G359), .O(gate103inter8));
  nand2 gate850(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate851(.a(s_43), .b(gate103inter3), .O(gate103inter10));
  nor2  gate852(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate853(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate854(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2213(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2214(.a(gate104inter0), .b(s_238), .O(gate104inter1));
  and2  gate2215(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2216(.a(s_238), .O(gate104inter3));
  inv1  gate2217(.a(s_239), .O(gate104inter4));
  nand2 gate2218(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2219(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2220(.a(G32), .O(gate104inter7));
  inv1  gate2221(.a(G359), .O(gate104inter8));
  nand2 gate2222(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2223(.a(s_239), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2224(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2225(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2226(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1891(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1892(.a(gate105inter0), .b(s_192), .O(gate105inter1));
  and2  gate1893(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1894(.a(s_192), .O(gate105inter3));
  inv1  gate1895(.a(s_193), .O(gate105inter4));
  nand2 gate1896(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1897(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1898(.a(G362), .O(gate105inter7));
  inv1  gate1899(.a(G363), .O(gate105inter8));
  nand2 gate1900(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1901(.a(s_193), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1902(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1903(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1904(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate673(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate674(.a(gate107inter0), .b(s_18), .O(gate107inter1));
  and2  gate675(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate676(.a(s_18), .O(gate107inter3));
  inv1  gate677(.a(s_19), .O(gate107inter4));
  nand2 gate678(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate679(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate680(.a(G366), .O(gate107inter7));
  inv1  gate681(.a(G367), .O(gate107inter8));
  nand2 gate682(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate683(.a(s_19), .b(gate107inter3), .O(gate107inter10));
  nor2  gate684(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate685(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate686(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate2241(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2242(.a(gate109inter0), .b(s_242), .O(gate109inter1));
  and2  gate2243(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2244(.a(s_242), .O(gate109inter3));
  inv1  gate2245(.a(s_243), .O(gate109inter4));
  nand2 gate2246(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2247(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2248(.a(G370), .O(gate109inter7));
  inv1  gate2249(.a(G371), .O(gate109inter8));
  nand2 gate2250(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2251(.a(s_243), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2252(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2253(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2254(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1065(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1066(.a(gate111inter0), .b(s_74), .O(gate111inter1));
  and2  gate1067(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1068(.a(s_74), .O(gate111inter3));
  inv1  gate1069(.a(s_75), .O(gate111inter4));
  nand2 gate1070(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1071(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1072(.a(G374), .O(gate111inter7));
  inv1  gate1073(.a(G375), .O(gate111inter8));
  nand2 gate1074(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1075(.a(s_75), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1076(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1077(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1078(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2073(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2074(.a(gate112inter0), .b(s_218), .O(gate112inter1));
  and2  gate2075(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2076(.a(s_218), .O(gate112inter3));
  inv1  gate2077(.a(s_219), .O(gate112inter4));
  nand2 gate2078(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2079(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2080(.a(G376), .O(gate112inter7));
  inv1  gate2081(.a(G377), .O(gate112inter8));
  nand2 gate2082(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2083(.a(s_219), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2084(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2085(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2086(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2031(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2032(.a(gate114inter0), .b(s_212), .O(gate114inter1));
  and2  gate2033(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2034(.a(s_212), .O(gate114inter3));
  inv1  gate2035(.a(s_213), .O(gate114inter4));
  nand2 gate2036(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2037(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2038(.a(G380), .O(gate114inter7));
  inv1  gate2039(.a(G381), .O(gate114inter8));
  nand2 gate2040(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2041(.a(s_213), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2042(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2043(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2044(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2437(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2438(.a(gate116inter0), .b(s_270), .O(gate116inter1));
  and2  gate2439(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2440(.a(s_270), .O(gate116inter3));
  inv1  gate2441(.a(s_271), .O(gate116inter4));
  nand2 gate2442(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2443(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2444(.a(G384), .O(gate116inter7));
  inv1  gate2445(.a(G385), .O(gate116inter8));
  nand2 gate2446(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2447(.a(s_271), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2448(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2449(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2450(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1639(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1640(.a(gate121inter0), .b(s_156), .O(gate121inter1));
  and2  gate1641(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1642(.a(s_156), .O(gate121inter3));
  inv1  gate1643(.a(s_157), .O(gate121inter4));
  nand2 gate1644(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1645(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1646(.a(G394), .O(gate121inter7));
  inv1  gate1647(.a(G395), .O(gate121inter8));
  nand2 gate1648(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1649(.a(s_157), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1650(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1651(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1652(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2871(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2872(.a(gate126inter0), .b(s_332), .O(gate126inter1));
  and2  gate2873(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2874(.a(s_332), .O(gate126inter3));
  inv1  gate2875(.a(s_333), .O(gate126inter4));
  nand2 gate2876(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2877(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2878(.a(G404), .O(gate126inter7));
  inv1  gate2879(.a(G405), .O(gate126inter8));
  nand2 gate2880(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2881(.a(s_333), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2882(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2883(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2884(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1723(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1724(.a(gate130inter0), .b(s_168), .O(gate130inter1));
  and2  gate1725(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1726(.a(s_168), .O(gate130inter3));
  inv1  gate1727(.a(s_169), .O(gate130inter4));
  nand2 gate1728(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1729(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1730(.a(G412), .O(gate130inter7));
  inv1  gate1731(.a(G413), .O(gate130inter8));
  nand2 gate1732(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1733(.a(s_169), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1734(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1735(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1736(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate785(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate786(.a(gate133inter0), .b(s_34), .O(gate133inter1));
  and2  gate787(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate788(.a(s_34), .O(gate133inter3));
  inv1  gate789(.a(s_35), .O(gate133inter4));
  nand2 gate790(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate791(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate792(.a(G418), .O(gate133inter7));
  inv1  gate793(.a(G419), .O(gate133inter8));
  nand2 gate794(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate795(.a(s_35), .b(gate133inter3), .O(gate133inter10));
  nor2  gate796(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate797(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate798(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate701(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate702(.a(gate135inter0), .b(s_22), .O(gate135inter1));
  and2  gate703(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate704(.a(s_22), .O(gate135inter3));
  inv1  gate705(.a(s_23), .O(gate135inter4));
  nand2 gate706(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate707(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate708(.a(G422), .O(gate135inter7));
  inv1  gate709(.a(G423), .O(gate135inter8));
  nand2 gate710(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate711(.a(s_23), .b(gate135inter3), .O(gate135inter10));
  nor2  gate712(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate713(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate714(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate2395(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2396(.a(gate136inter0), .b(s_264), .O(gate136inter1));
  and2  gate2397(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2398(.a(s_264), .O(gate136inter3));
  inv1  gate2399(.a(s_265), .O(gate136inter4));
  nand2 gate2400(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2401(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2402(.a(G424), .O(gate136inter7));
  inv1  gate2403(.a(G425), .O(gate136inter8));
  nand2 gate2404(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2405(.a(s_265), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2406(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2407(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2408(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate3249(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate3250(.a(gate141inter0), .b(s_386), .O(gate141inter1));
  and2  gate3251(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate3252(.a(s_386), .O(gate141inter3));
  inv1  gate3253(.a(s_387), .O(gate141inter4));
  nand2 gate3254(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate3255(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate3256(.a(G450), .O(gate141inter7));
  inv1  gate3257(.a(G453), .O(gate141inter8));
  nand2 gate3258(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate3259(.a(s_387), .b(gate141inter3), .O(gate141inter10));
  nor2  gate3260(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate3261(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate3262(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1877(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1878(.a(gate146inter0), .b(s_190), .O(gate146inter1));
  and2  gate1879(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1880(.a(s_190), .O(gate146inter3));
  inv1  gate1881(.a(s_191), .O(gate146inter4));
  nand2 gate1882(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1883(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1884(.a(G480), .O(gate146inter7));
  inv1  gate1885(.a(G483), .O(gate146inter8));
  nand2 gate1886(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1887(.a(s_191), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1888(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1889(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1890(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2339(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2340(.a(gate150inter0), .b(s_256), .O(gate150inter1));
  and2  gate2341(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2342(.a(s_256), .O(gate150inter3));
  inv1  gate2343(.a(s_257), .O(gate150inter4));
  nand2 gate2344(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2345(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2346(.a(G504), .O(gate150inter7));
  inv1  gate2347(.a(G507), .O(gate150inter8));
  nand2 gate2348(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2349(.a(s_257), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2350(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2351(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2352(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1499(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1500(.a(gate151inter0), .b(s_136), .O(gate151inter1));
  and2  gate1501(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1502(.a(s_136), .O(gate151inter3));
  inv1  gate1503(.a(s_137), .O(gate151inter4));
  nand2 gate1504(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1505(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1506(.a(G510), .O(gate151inter7));
  inv1  gate1507(.a(G513), .O(gate151inter8));
  nand2 gate1508(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1509(.a(s_137), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1510(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1511(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1512(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2283(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2284(.a(gate155inter0), .b(s_248), .O(gate155inter1));
  and2  gate2285(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2286(.a(s_248), .O(gate155inter3));
  inv1  gate2287(.a(s_249), .O(gate155inter4));
  nand2 gate2288(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2289(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2290(.a(G432), .O(gate155inter7));
  inv1  gate2291(.a(G525), .O(gate155inter8));
  nand2 gate2292(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2293(.a(s_249), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2294(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2295(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2296(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2325(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2326(.a(gate156inter0), .b(s_254), .O(gate156inter1));
  and2  gate2327(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2328(.a(s_254), .O(gate156inter3));
  inv1  gate2329(.a(s_255), .O(gate156inter4));
  nand2 gate2330(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2331(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2332(.a(G435), .O(gate156inter7));
  inv1  gate2333(.a(G525), .O(gate156inter8));
  nand2 gate2334(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2335(.a(s_255), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2336(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2337(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2338(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2549(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2550(.a(gate157inter0), .b(s_286), .O(gate157inter1));
  and2  gate2551(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2552(.a(s_286), .O(gate157inter3));
  inv1  gate2553(.a(s_287), .O(gate157inter4));
  nand2 gate2554(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2555(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2556(.a(G438), .O(gate157inter7));
  inv1  gate2557(.a(G528), .O(gate157inter8));
  nand2 gate2558(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2559(.a(s_287), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2560(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2561(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2562(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2521(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2522(.a(gate159inter0), .b(s_282), .O(gate159inter1));
  and2  gate2523(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2524(.a(s_282), .O(gate159inter3));
  inv1  gate2525(.a(s_283), .O(gate159inter4));
  nand2 gate2526(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2527(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2528(.a(G444), .O(gate159inter7));
  inv1  gate2529(.a(G531), .O(gate159inter8));
  nand2 gate2530(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2531(.a(s_283), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2532(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2533(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2534(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate659(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate660(.a(gate161inter0), .b(s_16), .O(gate161inter1));
  and2  gate661(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate662(.a(s_16), .O(gate161inter3));
  inv1  gate663(.a(s_17), .O(gate161inter4));
  nand2 gate664(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate665(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate666(.a(G450), .O(gate161inter7));
  inv1  gate667(.a(G534), .O(gate161inter8));
  nand2 gate668(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate669(.a(s_17), .b(gate161inter3), .O(gate161inter10));
  nor2  gate670(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate671(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate672(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1709(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1710(.a(gate163inter0), .b(s_166), .O(gate163inter1));
  and2  gate1711(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1712(.a(s_166), .O(gate163inter3));
  inv1  gate1713(.a(s_167), .O(gate163inter4));
  nand2 gate1714(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1715(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1716(.a(G456), .O(gate163inter7));
  inv1  gate1717(.a(G537), .O(gate163inter8));
  nand2 gate1718(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1719(.a(s_167), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1720(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1721(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1722(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2745(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2746(.a(gate164inter0), .b(s_314), .O(gate164inter1));
  and2  gate2747(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2748(.a(s_314), .O(gate164inter3));
  inv1  gate2749(.a(s_315), .O(gate164inter4));
  nand2 gate2750(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2751(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2752(.a(G459), .O(gate164inter7));
  inv1  gate2753(.a(G537), .O(gate164inter8));
  nand2 gate2754(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2755(.a(s_315), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2756(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2757(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2758(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1079(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1080(.a(gate173inter0), .b(s_76), .O(gate173inter1));
  and2  gate1081(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1082(.a(s_76), .O(gate173inter3));
  inv1  gate1083(.a(s_77), .O(gate173inter4));
  nand2 gate1084(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1085(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1086(.a(G486), .O(gate173inter7));
  inv1  gate1087(.a(G552), .O(gate173inter8));
  nand2 gate1088(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1089(.a(s_77), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1090(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1091(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1092(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1653(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1654(.a(gate174inter0), .b(s_158), .O(gate174inter1));
  and2  gate1655(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1656(.a(s_158), .O(gate174inter3));
  inv1  gate1657(.a(s_159), .O(gate174inter4));
  nand2 gate1658(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1659(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1660(.a(G489), .O(gate174inter7));
  inv1  gate1661(.a(G552), .O(gate174inter8));
  nand2 gate1662(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1663(.a(s_159), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1664(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1665(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1666(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2885(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2886(.a(gate175inter0), .b(s_334), .O(gate175inter1));
  and2  gate2887(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2888(.a(s_334), .O(gate175inter3));
  inv1  gate2889(.a(s_335), .O(gate175inter4));
  nand2 gate2890(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2891(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2892(.a(G492), .O(gate175inter7));
  inv1  gate2893(.a(G555), .O(gate175inter8));
  nand2 gate2894(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2895(.a(s_335), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2896(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2897(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2898(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1513(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1514(.a(gate180inter0), .b(s_138), .O(gate180inter1));
  and2  gate1515(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1516(.a(s_138), .O(gate180inter3));
  inv1  gate1517(.a(s_139), .O(gate180inter4));
  nand2 gate1518(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1519(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1520(.a(G507), .O(gate180inter7));
  inv1  gate1521(.a(G561), .O(gate180inter8));
  nand2 gate1522(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1523(.a(s_139), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1524(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1525(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1526(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate2577(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2578(.a(gate181inter0), .b(s_290), .O(gate181inter1));
  and2  gate2579(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2580(.a(s_290), .O(gate181inter3));
  inv1  gate2581(.a(s_291), .O(gate181inter4));
  nand2 gate2582(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2583(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2584(.a(G510), .O(gate181inter7));
  inv1  gate2585(.a(G564), .O(gate181inter8));
  nand2 gate2586(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2587(.a(s_291), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2588(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2589(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2590(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1233(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1234(.a(gate183inter0), .b(s_98), .O(gate183inter1));
  and2  gate1235(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1236(.a(s_98), .O(gate183inter3));
  inv1  gate1237(.a(s_99), .O(gate183inter4));
  nand2 gate1238(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1239(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1240(.a(G516), .O(gate183inter7));
  inv1  gate1241(.a(G567), .O(gate183inter8));
  nand2 gate1242(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1243(.a(s_99), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1244(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1245(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1246(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1205(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1206(.a(gate184inter0), .b(s_94), .O(gate184inter1));
  and2  gate1207(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1208(.a(s_94), .O(gate184inter3));
  inv1  gate1209(.a(s_95), .O(gate184inter4));
  nand2 gate1210(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1211(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1212(.a(G519), .O(gate184inter7));
  inv1  gate1213(.a(G567), .O(gate184inter8));
  nand2 gate1214(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1215(.a(s_95), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1216(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1217(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1218(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1611(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1612(.a(gate188inter0), .b(s_152), .O(gate188inter1));
  and2  gate1613(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1614(.a(s_152), .O(gate188inter3));
  inv1  gate1615(.a(s_153), .O(gate188inter4));
  nand2 gate1616(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1617(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1618(.a(G576), .O(gate188inter7));
  inv1  gate1619(.a(G577), .O(gate188inter8));
  nand2 gate1620(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1621(.a(s_153), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1622(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1623(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1624(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1583(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1584(.a(gate193inter0), .b(s_148), .O(gate193inter1));
  and2  gate1585(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1586(.a(s_148), .O(gate193inter3));
  inv1  gate1587(.a(s_149), .O(gate193inter4));
  nand2 gate1588(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1589(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1590(.a(G586), .O(gate193inter7));
  inv1  gate1591(.a(G587), .O(gate193inter8));
  nand2 gate1592(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1593(.a(s_149), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1594(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1595(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1596(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1317(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1318(.a(gate194inter0), .b(s_110), .O(gate194inter1));
  and2  gate1319(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1320(.a(s_110), .O(gate194inter3));
  inv1  gate1321(.a(s_111), .O(gate194inter4));
  nand2 gate1322(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1323(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1324(.a(G588), .O(gate194inter7));
  inv1  gate1325(.a(G589), .O(gate194inter8));
  nand2 gate1326(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1327(.a(s_111), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1328(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1329(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1330(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2381(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2382(.a(gate195inter0), .b(s_262), .O(gate195inter1));
  and2  gate2383(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2384(.a(s_262), .O(gate195inter3));
  inv1  gate2385(.a(s_263), .O(gate195inter4));
  nand2 gate2386(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2387(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2388(.a(G590), .O(gate195inter7));
  inv1  gate2389(.a(G591), .O(gate195inter8));
  nand2 gate2390(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2391(.a(s_263), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2392(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2393(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2394(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2451(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2452(.a(gate198inter0), .b(s_272), .O(gate198inter1));
  and2  gate2453(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2454(.a(s_272), .O(gate198inter3));
  inv1  gate2455(.a(s_273), .O(gate198inter4));
  nand2 gate2456(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2457(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2458(.a(G596), .O(gate198inter7));
  inv1  gate2459(.a(G597), .O(gate198inter8));
  nand2 gate2460(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2461(.a(s_273), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2462(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2463(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2464(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2017(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2018(.a(gate200inter0), .b(s_210), .O(gate200inter1));
  and2  gate2019(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2020(.a(s_210), .O(gate200inter3));
  inv1  gate2021(.a(s_211), .O(gate200inter4));
  nand2 gate2022(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2023(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2024(.a(G600), .O(gate200inter7));
  inv1  gate2025(.a(G601), .O(gate200inter8));
  nand2 gate2026(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2027(.a(s_211), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2028(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2029(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2030(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1275(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1276(.a(gate204inter0), .b(s_104), .O(gate204inter1));
  and2  gate1277(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1278(.a(s_104), .O(gate204inter3));
  inv1  gate1279(.a(s_105), .O(gate204inter4));
  nand2 gate1280(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1281(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1282(.a(G607), .O(gate204inter7));
  inv1  gate1283(.a(G617), .O(gate204inter8));
  nand2 gate1284(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1285(.a(s_105), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1286(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1287(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1288(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1373(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1374(.a(gate206inter0), .b(s_118), .O(gate206inter1));
  and2  gate1375(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1376(.a(s_118), .O(gate206inter3));
  inv1  gate1377(.a(s_119), .O(gate206inter4));
  nand2 gate1378(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1379(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1380(.a(G632), .O(gate206inter7));
  inv1  gate1381(.a(G637), .O(gate206inter8));
  nand2 gate1382(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1383(.a(s_119), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1384(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1385(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1386(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1429(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1430(.a(gate210inter0), .b(s_126), .O(gate210inter1));
  and2  gate1431(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1432(.a(s_126), .O(gate210inter3));
  inv1  gate1433(.a(s_127), .O(gate210inter4));
  nand2 gate1434(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1435(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1436(.a(G607), .O(gate210inter7));
  inv1  gate1437(.a(G666), .O(gate210inter8));
  nand2 gate1438(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1439(.a(s_127), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1440(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1441(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1442(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1457(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1458(.a(gate213inter0), .b(s_130), .O(gate213inter1));
  and2  gate1459(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1460(.a(s_130), .O(gate213inter3));
  inv1  gate1461(.a(s_131), .O(gate213inter4));
  nand2 gate1462(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1463(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1464(.a(G602), .O(gate213inter7));
  inv1  gate1465(.a(G672), .O(gate213inter8));
  nand2 gate1466(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1467(.a(s_131), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1468(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1469(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1470(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate995(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate996(.a(gate214inter0), .b(s_64), .O(gate214inter1));
  and2  gate997(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate998(.a(s_64), .O(gate214inter3));
  inv1  gate999(.a(s_65), .O(gate214inter4));
  nand2 gate1000(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1001(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1002(.a(G612), .O(gate214inter7));
  inv1  gate1003(.a(G672), .O(gate214inter8));
  nand2 gate1004(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1005(.a(s_65), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1006(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1007(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1008(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate3193(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate3194(.a(gate217inter0), .b(s_378), .O(gate217inter1));
  and2  gate3195(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate3196(.a(s_378), .O(gate217inter3));
  inv1  gate3197(.a(s_379), .O(gate217inter4));
  nand2 gate3198(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate3199(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate3200(.a(G622), .O(gate217inter7));
  inv1  gate3201(.a(G678), .O(gate217inter8));
  nand2 gate3202(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate3203(.a(s_379), .b(gate217inter3), .O(gate217inter10));
  nor2  gate3204(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate3205(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate3206(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2199(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2200(.a(gate222inter0), .b(s_236), .O(gate222inter1));
  and2  gate2201(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2202(.a(s_236), .O(gate222inter3));
  inv1  gate2203(.a(s_237), .O(gate222inter4));
  nand2 gate2204(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2205(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2206(.a(G632), .O(gate222inter7));
  inv1  gate2207(.a(G684), .O(gate222inter8));
  nand2 gate2208(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2209(.a(s_237), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2210(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2211(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2212(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2941(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2942(.a(gate224inter0), .b(s_342), .O(gate224inter1));
  and2  gate2943(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2944(.a(s_342), .O(gate224inter3));
  inv1  gate2945(.a(s_343), .O(gate224inter4));
  nand2 gate2946(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2947(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2948(.a(G637), .O(gate224inter7));
  inv1  gate2949(.a(G687), .O(gate224inter8));
  nand2 gate2950(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2951(.a(s_343), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2952(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2953(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2954(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate3179(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate3180(.a(gate225inter0), .b(s_376), .O(gate225inter1));
  and2  gate3181(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate3182(.a(s_376), .O(gate225inter3));
  inv1  gate3183(.a(s_377), .O(gate225inter4));
  nand2 gate3184(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate3185(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate3186(.a(G690), .O(gate225inter7));
  inv1  gate3187(.a(G691), .O(gate225inter8));
  nand2 gate3188(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate3189(.a(s_377), .b(gate225inter3), .O(gate225inter10));
  nor2  gate3190(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate3191(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate3192(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1289(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1290(.a(gate226inter0), .b(s_106), .O(gate226inter1));
  and2  gate1291(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1292(.a(s_106), .O(gate226inter3));
  inv1  gate1293(.a(s_107), .O(gate226inter4));
  nand2 gate1294(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1295(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1296(.a(G692), .O(gate226inter7));
  inv1  gate1297(.a(G693), .O(gate226inter8));
  nand2 gate1298(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1299(.a(s_107), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1300(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1301(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1302(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate2311(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2312(.a(gate227inter0), .b(s_252), .O(gate227inter1));
  and2  gate2313(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2314(.a(s_252), .O(gate227inter3));
  inv1  gate2315(.a(s_253), .O(gate227inter4));
  nand2 gate2316(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2317(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2318(.a(G694), .O(gate227inter7));
  inv1  gate2319(.a(G695), .O(gate227inter8));
  nand2 gate2320(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2321(.a(s_253), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2322(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2323(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2324(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate2927(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2928(.a(gate228inter0), .b(s_340), .O(gate228inter1));
  and2  gate2929(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2930(.a(s_340), .O(gate228inter3));
  inv1  gate2931(.a(s_341), .O(gate228inter4));
  nand2 gate2932(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2933(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2934(.a(G696), .O(gate228inter7));
  inv1  gate2935(.a(G697), .O(gate228inter8));
  nand2 gate2936(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2937(.a(s_341), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2938(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2939(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2940(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2045(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2046(.a(gate230inter0), .b(s_214), .O(gate230inter1));
  and2  gate2047(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2048(.a(s_214), .O(gate230inter3));
  inv1  gate2049(.a(s_215), .O(gate230inter4));
  nand2 gate2050(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2051(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2052(.a(G700), .O(gate230inter7));
  inv1  gate2053(.a(G701), .O(gate230inter8));
  nand2 gate2054(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2055(.a(s_215), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2056(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2057(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2058(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate771(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate772(.a(gate232inter0), .b(s_32), .O(gate232inter1));
  and2  gate773(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate774(.a(s_32), .O(gate232inter3));
  inv1  gate775(.a(s_33), .O(gate232inter4));
  nand2 gate776(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate777(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate778(.a(G704), .O(gate232inter7));
  inv1  gate779(.a(G705), .O(gate232inter8));
  nand2 gate780(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate781(.a(s_33), .b(gate232inter3), .O(gate232inter10));
  nor2  gate782(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate783(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate784(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate3011(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate3012(.a(gate233inter0), .b(s_352), .O(gate233inter1));
  and2  gate3013(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate3014(.a(s_352), .O(gate233inter3));
  inv1  gate3015(.a(s_353), .O(gate233inter4));
  nand2 gate3016(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate3017(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate3018(.a(G242), .O(gate233inter7));
  inv1  gate3019(.a(G718), .O(gate233inter8));
  nand2 gate3020(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate3021(.a(s_353), .b(gate233inter3), .O(gate233inter10));
  nor2  gate3022(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate3023(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate3024(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1149(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1150(.a(gate234inter0), .b(s_86), .O(gate234inter1));
  and2  gate1151(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1152(.a(s_86), .O(gate234inter3));
  inv1  gate1153(.a(s_87), .O(gate234inter4));
  nand2 gate1154(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1155(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1156(.a(G245), .O(gate234inter7));
  inv1  gate1157(.a(G721), .O(gate234inter8));
  nand2 gate1158(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1159(.a(s_87), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1160(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1161(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1162(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1107(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1108(.a(gate235inter0), .b(s_80), .O(gate235inter1));
  and2  gate1109(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1110(.a(s_80), .O(gate235inter3));
  inv1  gate1111(.a(s_81), .O(gate235inter4));
  nand2 gate1112(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1113(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1114(.a(G248), .O(gate235inter7));
  inv1  gate1115(.a(G724), .O(gate235inter8));
  nand2 gate1116(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1117(.a(s_81), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1118(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1119(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1120(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2115(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2116(.a(gate238inter0), .b(s_224), .O(gate238inter1));
  and2  gate2117(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2118(.a(s_224), .O(gate238inter3));
  inv1  gate2119(.a(s_225), .O(gate238inter4));
  nand2 gate2120(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2121(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2122(.a(G257), .O(gate238inter7));
  inv1  gate2123(.a(G709), .O(gate238inter8));
  nand2 gate2124(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2125(.a(s_225), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2126(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2127(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2128(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2829(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2830(.a(gate239inter0), .b(s_326), .O(gate239inter1));
  and2  gate2831(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2832(.a(s_326), .O(gate239inter3));
  inv1  gate2833(.a(s_327), .O(gate239inter4));
  nand2 gate2834(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2835(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2836(.a(G260), .O(gate239inter7));
  inv1  gate2837(.a(G712), .O(gate239inter8));
  nand2 gate2838(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2839(.a(s_327), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2840(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2841(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2842(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1037(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1038(.a(gate242inter0), .b(s_70), .O(gate242inter1));
  and2  gate1039(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1040(.a(s_70), .O(gate242inter3));
  inv1  gate1041(.a(s_71), .O(gate242inter4));
  nand2 gate1042(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1043(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1044(.a(G718), .O(gate242inter7));
  inv1  gate1045(.a(G730), .O(gate242inter8));
  nand2 gate1046(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1047(.a(s_71), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1048(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1049(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1050(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate631(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate632(.a(gate244inter0), .b(s_12), .O(gate244inter1));
  and2  gate633(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate634(.a(s_12), .O(gate244inter3));
  inv1  gate635(.a(s_13), .O(gate244inter4));
  nand2 gate636(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate637(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate638(.a(G721), .O(gate244inter7));
  inv1  gate639(.a(G733), .O(gate244inter8));
  nand2 gate640(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate641(.a(s_13), .b(gate244inter3), .O(gate244inter10));
  nor2  gate642(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate643(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate644(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1569(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1570(.a(gate246inter0), .b(s_146), .O(gate246inter1));
  and2  gate1571(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1572(.a(s_146), .O(gate246inter3));
  inv1  gate1573(.a(s_147), .O(gate246inter4));
  nand2 gate1574(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1575(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1576(.a(G724), .O(gate246inter7));
  inv1  gate1577(.a(G736), .O(gate246inter8));
  nand2 gate1578(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1579(.a(s_147), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1580(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1581(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1582(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1961(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1962(.a(gate247inter0), .b(s_202), .O(gate247inter1));
  and2  gate1963(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1964(.a(s_202), .O(gate247inter3));
  inv1  gate1965(.a(s_203), .O(gate247inter4));
  nand2 gate1966(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1967(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1968(.a(G251), .O(gate247inter7));
  inv1  gate1969(.a(G739), .O(gate247inter8));
  nand2 gate1970(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1971(.a(s_203), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1972(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1973(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1974(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2367(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2368(.a(gate249inter0), .b(s_260), .O(gate249inter1));
  and2  gate2369(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2370(.a(s_260), .O(gate249inter3));
  inv1  gate2371(.a(s_261), .O(gate249inter4));
  nand2 gate2372(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2373(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2374(.a(G254), .O(gate249inter7));
  inv1  gate2375(.a(G742), .O(gate249inter8));
  nand2 gate2376(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2377(.a(s_261), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2378(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2379(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2380(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate897(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate898(.a(gate250inter0), .b(s_50), .O(gate250inter1));
  and2  gate899(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate900(.a(s_50), .O(gate250inter3));
  inv1  gate901(.a(s_51), .O(gate250inter4));
  nand2 gate902(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate903(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate904(.a(G706), .O(gate250inter7));
  inv1  gate905(.a(G742), .O(gate250inter8));
  nand2 gate906(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate907(.a(s_51), .b(gate250inter3), .O(gate250inter10));
  nor2  gate908(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate909(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate910(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2857(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2858(.a(gate251inter0), .b(s_330), .O(gate251inter1));
  and2  gate2859(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2860(.a(s_330), .O(gate251inter3));
  inv1  gate2861(.a(s_331), .O(gate251inter4));
  nand2 gate2862(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2863(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2864(.a(G257), .O(gate251inter7));
  inv1  gate2865(.a(G745), .O(gate251inter8));
  nand2 gate2866(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2867(.a(s_331), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2868(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2869(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2870(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2465(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2466(.a(gate254inter0), .b(s_274), .O(gate254inter1));
  and2  gate2467(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2468(.a(s_274), .O(gate254inter3));
  inv1  gate2469(.a(s_275), .O(gate254inter4));
  nand2 gate2470(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2471(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2472(.a(G712), .O(gate254inter7));
  inv1  gate2473(.a(G748), .O(gate254inter8));
  nand2 gate2474(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2475(.a(s_275), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2476(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2477(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2478(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1667(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1668(.a(gate255inter0), .b(s_160), .O(gate255inter1));
  and2  gate1669(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1670(.a(s_160), .O(gate255inter3));
  inv1  gate1671(.a(s_161), .O(gate255inter4));
  nand2 gate1672(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1673(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1674(.a(G263), .O(gate255inter7));
  inv1  gate1675(.a(G751), .O(gate255inter8));
  nand2 gate1676(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1677(.a(s_161), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1678(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1679(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1680(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2913(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2914(.a(gate261inter0), .b(s_338), .O(gate261inter1));
  and2  gate2915(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2916(.a(s_338), .O(gate261inter3));
  inv1  gate2917(.a(s_339), .O(gate261inter4));
  nand2 gate2918(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2919(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2920(.a(G762), .O(gate261inter7));
  inv1  gate2921(.a(G763), .O(gate261inter8));
  nand2 gate2922(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2923(.a(s_339), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2924(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2925(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2926(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate603(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate604(.a(gate262inter0), .b(s_8), .O(gate262inter1));
  and2  gate605(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate606(.a(s_8), .O(gate262inter3));
  inv1  gate607(.a(s_9), .O(gate262inter4));
  nand2 gate608(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate609(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate610(.a(G764), .O(gate262inter7));
  inv1  gate611(.a(G765), .O(gate262inter8));
  nand2 gate612(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate613(.a(s_9), .b(gate262inter3), .O(gate262inter10));
  nor2  gate614(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate615(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate616(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate967(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate968(.a(gate263inter0), .b(s_60), .O(gate263inter1));
  and2  gate969(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate970(.a(s_60), .O(gate263inter3));
  inv1  gate971(.a(s_61), .O(gate263inter4));
  nand2 gate972(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate973(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate974(.a(G766), .O(gate263inter7));
  inv1  gate975(.a(G767), .O(gate263inter8));
  nand2 gate976(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate977(.a(s_61), .b(gate263inter3), .O(gate263inter10));
  nor2  gate978(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate979(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate980(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate3165(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate3166(.a(gate268inter0), .b(s_374), .O(gate268inter1));
  and2  gate3167(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate3168(.a(s_374), .O(gate268inter3));
  inv1  gate3169(.a(s_375), .O(gate268inter4));
  nand2 gate3170(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate3171(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate3172(.a(G651), .O(gate268inter7));
  inv1  gate3173(.a(G779), .O(gate268inter8));
  nand2 gate3174(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate3175(.a(s_375), .b(gate268inter3), .O(gate268inter10));
  nor2  gate3176(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate3177(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate3178(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2101(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2102(.a(gate271inter0), .b(s_222), .O(gate271inter1));
  and2  gate2103(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2104(.a(s_222), .O(gate271inter3));
  inv1  gate2105(.a(s_223), .O(gate271inter4));
  nand2 gate2106(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2107(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2108(.a(G660), .O(gate271inter7));
  inv1  gate2109(.a(G788), .O(gate271inter8));
  nand2 gate2110(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2111(.a(s_223), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2112(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2113(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2114(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1331(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1332(.a(gate274inter0), .b(s_112), .O(gate274inter1));
  and2  gate1333(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1334(.a(s_112), .O(gate274inter3));
  inv1  gate1335(.a(s_113), .O(gate274inter4));
  nand2 gate1336(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1337(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1338(.a(G770), .O(gate274inter7));
  inv1  gate1339(.a(G794), .O(gate274inter8));
  nand2 gate1340(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1341(.a(s_113), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1342(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1343(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1344(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1247(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1248(.a(gate279inter0), .b(s_100), .O(gate279inter1));
  and2  gate1249(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1250(.a(s_100), .O(gate279inter3));
  inv1  gate1251(.a(s_101), .O(gate279inter4));
  nand2 gate1252(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1253(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1254(.a(G651), .O(gate279inter7));
  inv1  gate1255(.a(G803), .O(gate279inter8));
  nand2 gate1256(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1257(.a(s_101), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1258(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1259(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1260(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate645(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate646(.a(gate280inter0), .b(s_14), .O(gate280inter1));
  and2  gate647(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate648(.a(s_14), .O(gate280inter3));
  inv1  gate649(.a(s_15), .O(gate280inter4));
  nand2 gate650(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate651(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate652(.a(G779), .O(gate280inter7));
  inv1  gate653(.a(G803), .O(gate280inter8));
  nand2 gate654(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate655(.a(s_15), .b(gate280inter3), .O(gate280inter10));
  nor2  gate656(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate657(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate658(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1527(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1528(.a(gate284inter0), .b(s_140), .O(gate284inter1));
  and2  gate1529(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1530(.a(s_140), .O(gate284inter3));
  inv1  gate1531(.a(s_141), .O(gate284inter4));
  nand2 gate1532(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1533(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1534(.a(G785), .O(gate284inter7));
  inv1  gate1535(.a(G809), .O(gate284inter8));
  nand2 gate1536(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1537(.a(s_141), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1538(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1539(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1540(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2423(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2424(.a(gate285inter0), .b(s_268), .O(gate285inter1));
  and2  gate2425(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2426(.a(s_268), .O(gate285inter3));
  inv1  gate2427(.a(s_269), .O(gate285inter4));
  nand2 gate2428(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2429(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2430(.a(G660), .O(gate285inter7));
  inv1  gate2431(.a(G812), .O(gate285inter8));
  nand2 gate2432(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2433(.a(s_269), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2434(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2435(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2436(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2129(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2130(.a(gate286inter0), .b(s_226), .O(gate286inter1));
  and2  gate2131(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2132(.a(s_226), .O(gate286inter3));
  inv1  gate2133(.a(s_227), .O(gate286inter4));
  nand2 gate2134(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2135(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2136(.a(G788), .O(gate286inter7));
  inv1  gate2137(.a(G812), .O(gate286inter8));
  nand2 gate2138(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2139(.a(s_227), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2140(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2141(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2142(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2591(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2592(.a(gate287inter0), .b(s_292), .O(gate287inter1));
  and2  gate2593(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2594(.a(s_292), .O(gate287inter3));
  inv1  gate2595(.a(s_293), .O(gate287inter4));
  nand2 gate2596(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2597(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2598(.a(G663), .O(gate287inter7));
  inv1  gate2599(.a(G815), .O(gate287inter8));
  nand2 gate2600(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2601(.a(s_293), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2602(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2603(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2604(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2619(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2620(.a(gate289inter0), .b(s_296), .O(gate289inter1));
  and2  gate2621(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2622(.a(s_296), .O(gate289inter3));
  inv1  gate2623(.a(s_297), .O(gate289inter4));
  nand2 gate2624(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2625(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2626(.a(G818), .O(gate289inter7));
  inv1  gate2627(.a(G819), .O(gate289inter8));
  nand2 gate2628(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2629(.a(s_297), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2630(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2631(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2632(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1933(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1934(.a(gate290inter0), .b(s_198), .O(gate290inter1));
  and2  gate1935(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1936(.a(s_198), .O(gate290inter3));
  inv1  gate1937(.a(s_199), .O(gate290inter4));
  nand2 gate1938(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1939(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1940(.a(G820), .O(gate290inter7));
  inv1  gate1941(.a(G821), .O(gate290inter8));
  nand2 gate1942(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1943(.a(s_199), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1944(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1945(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1946(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1863(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1864(.a(gate291inter0), .b(s_188), .O(gate291inter1));
  and2  gate1865(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1866(.a(s_188), .O(gate291inter3));
  inv1  gate1867(.a(s_189), .O(gate291inter4));
  nand2 gate1868(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1869(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1870(.a(G822), .O(gate291inter7));
  inv1  gate1871(.a(G823), .O(gate291inter8));
  nand2 gate1872(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1873(.a(s_189), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1874(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1875(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1876(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1303(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1304(.a(gate293inter0), .b(s_108), .O(gate293inter1));
  and2  gate1305(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1306(.a(s_108), .O(gate293inter3));
  inv1  gate1307(.a(s_109), .O(gate293inter4));
  nand2 gate1308(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1309(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1310(.a(G828), .O(gate293inter7));
  inv1  gate1311(.a(G829), .O(gate293inter8));
  nand2 gate1312(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1313(.a(s_109), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1314(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1315(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1316(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2899(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2900(.a(gate294inter0), .b(s_336), .O(gate294inter1));
  and2  gate2901(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2902(.a(s_336), .O(gate294inter3));
  inv1  gate2903(.a(s_337), .O(gate294inter4));
  nand2 gate2904(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2905(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2906(.a(G832), .O(gate294inter7));
  inv1  gate2907(.a(G833), .O(gate294inter8));
  nand2 gate2908(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2909(.a(s_337), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2910(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2911(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2912(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1597(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1598(.a(gate389inter0), .b(s_150), .O(gate389inter1));
  and2  gate1599(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1600(.a(s_150), .O(gate389inter3));
  inv1  gate1601(.a(s_151), .O(gate389inter4));
  nand2 gate1602(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1603(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1604(.a(G3), .O(gate389inter7));
  inv1  gate1605(.a(G1042), .O(gate389inter8));
  nand2 gate1606(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1607(.a(s_151), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1608(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1609(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1610(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1849(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1850(.a(gate392inter0), .b(s_186), .O(gate392inter1));
  and2  gate1851(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1852(.a(s_186), .O(gate392inter3));
  inv1  gate1853(.a(s_187), .O(gate392inter4));
  nand2 gate1854(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1855(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1856(.a(G6), .O(gate392inter7));
  inv1  gate1857(.a(G1051), .O(gate392inter8));
  nand2 gate1858(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1859(.a(s_187), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1860(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1861(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1862(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1261(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1262(.a(gate393inter0), .b(s_102), .O(gate393inter1));
  and2  gate1263(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1264(.a(s_102), .O(gate393inter3));
  inv1  gate1265(.a(s_103), .O(gate393inter4));
  nand2 gate1266(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1267(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1268(.a(G7), .O(gate393inter7));
  inv1  gate1269(.a(G1054), .O(gate393inter8));
  nand2 gate1270(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1271(.a(s_103), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1272(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1273(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1274(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2507(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2508(.a(gate398inter0), .b(s_280), .O(gate398inter1));
  and2  gate2509(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2510(.a(s_280), .O(gate398inter3));
  inv1  gate2511(.a(s_281), .O(gate398inter4));
  nand2 gate2512(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2513(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2514(.a(G12), .O(gate398inter7));
  inv1  gate2515(.a(G1069), .O(gate398inter8));
  nand2 gate2516(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2517(.a(s_281), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2518(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2519(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2520(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2409(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2410(.a(gate402inter0), .b(s_266), .O(gate402inter1));
  and2  gate2411(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2412(.a(s_266), .O(gate402inter3));
  inv1  gate2413(.a(s_267), .O(gate402inter4));
  nand2 gate2414(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2415(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2416(.a(G16), .O(gate402inter7));
  inv1  gate2417(.a(G1081), .O(gate402inter8));
  nand2 gate2418(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2419(.a(s_267), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2420(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2421(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2422(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1359(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1360(.a(gate403inter0), .b(s_116), .O(gate403inter1));
  and2  gate1361(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1362(.a(s_116), .O(gate403inter3));
  inv1  gate1363(.a(s_117), .O(gate403inter4));
  nand2 gate1364(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1365(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1366(.a(G17), .O(gate403inter7));
  inv1  gate1367(.a(G1084), .O(gate403inter8));
  nand2 gate1368(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1369(.a(s_117), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1370(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1371(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1372(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2605(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2606(.a(gate410inter0), .b(s_294), .O(gate410inter1));
  and2  gate2607(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2608(.a(s_294), .O(gate410inter3));
  inv1  gate2609(.a(s_295), .O(gate410inter4));
  nand2 gate2610(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2611(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2612(.a(G24), .O(gate410inter7));
  inv1  gate2613(.a(G1105), .O(gate410inter8));
  nand2 gate2614(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2615(.a(s_295), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2616(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2617(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2618(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2773(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2774(.a(gate412inter0), .b(s_318), .O(gate412inter1));
  and2  gate2775(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2776(.a(s_318), .O(gate412inter3));
  inv1  gate2777(.a(s_319), .O(gate412inter4));
  nand2 gate2778(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2779(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2780(.a(G26), .O(gate412inter7));
  inv1  gate2781(.a(G1111), .O(gate412inter8));
  nand2 gate2782(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2783(.a(s_319), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2784(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2785(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2786(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1625(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1626(.a(gate413inter0), .b(s_154), .O(gate413inter1));
  and2  gate1627(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1628(.a(s_154), .O(gate413inter3));
  inv1  gate1629(.a(s_155), .O(gate413inter4));
  nand2 gate1630(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1631(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1632(.a(G27), .O(gate413inter7));
  inv1  gate1633(.a(G1114), .O(gate413inter8));
  nand2 gate1634(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1635(.a(s_155), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1636(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1637(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1638(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate617(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate618(.a(gate414inter0), .b(s_10), .O(gate414inter1));
  and2  gate619(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate620(.a(s_10), .O(gate414inter3));
  inv1  gate621(.a(s_11), .O(gate414inter4));
  nand2 gate622(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate623(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate624(.a(G28), .O(gate414inter7));
  inv1  gate625(.a(G1117), .O(gate414inter8));
  nand2 gate626(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate627(.a(s_11), .b(gate414inter3), .O(gate414inter10));
  nor2  gate628(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate629(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate630(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate687(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate688(.a(gate416inter0), .b(s_20), .O(gate416inter1));
  and2  gate689(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate690(.a(s_20), .O(gate416inter3));
  inv1  gate691(.a(s_21), .O(gate416inter4));
  nand2 gate692(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate693(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate694(.a(G30), .O(gate416inter7));
  inv1  gate695(.a(G1123), .O(gate416inter8));
  nand2 gate696(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate697(.a(s_21), .b(gate416inter3), .O(gate416inter10));
  nor2  gate698(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate699(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate700(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2157(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2158(.a(gate417inter0), .b(s_230), .O(gate417inter1));
  and2  gate2159(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2160(.a(s_230), .O(gate417inter3));
  inv1  gate2161(.a(s_231), .O(gate417inter4));
  nand2 gate2162(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2163(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2164(.a(G31), .O(gate417inter7));
  inv1  gate2165(.a(G1126), .O(gate417inter8));
  nand2 gate2166(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2167(.a(s_231), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2168(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2169(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2170(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate925(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate926(.a(gate419inter0), .b(s_54), .O(gate419inter1));
  and2  gate927(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate928(.a(s_54), .O(gate419inter3));
  inv1  gate929(.a(s_55), .O(gate419inter4));
  nand2 gate930(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate931(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate932(.a(G1), .O(gate419inter7));
  inv1  gate933(.a(G1132), .O(gate419inter8));
  nand2 gate934(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate935(.a(s_55), .b(gate419inter3), .O(gate419inter10));
  nor2  gate936(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate937(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate938(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2255(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2256(.a(gate420inter0), .b(s_244), .O(gate420inter1));
  and2  gate2257(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2258(.a(s_244), .O(gate420inter3));
  inv1  gate2259(.a(s_245), .O(gate420inter4));
  nand2 gate2260(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2261(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2262(.a(G1036), .O(gate420inter7));
  inv1  gate2263(.a(G1132), .O(gate420inter8));
  nand2 gate2264(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2265(.a(s_245), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2266(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2267(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2268(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate827(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate828(.a(gate421inter0), .b(s_40), .O(gate421inter1));
  and2  gate829(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate830(.a(s_40), .O(gate421inter3));
  inv1  gate831(.a(s_41), .O(gate421inter4));
  nand2 gate832(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate833(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate834(.a(G2), .O(gate421inter7));
  inv1  gate835(.a(G1135), .O(gate421inter8));
  nand2 gate836(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate837(.a(s_41), .b(gate421inter3), .O(gate421inter10));
  nor2  gate838(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate839(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate840(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2717(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2718(.a(gate423inter0), .b(s_310), .O(gate423inter1));
  and2  gate2719(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2720(.a(s_310), .O(gate423inter3));
  inv1  gate2721(.a(s_311), .O(gate423inter4));
  nand2 gate2722(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2723(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2724(.a(G3), .O(gate423inter7));
  inv1  gate2725(.a(G1138), .O(gate423inter8));
  nand2 gate2726(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2727(.a(s_311), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2728(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2729(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2730(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2269(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2270(.a(gate424inter0), .b(s_246), .O(gate424inter1));
  and2  gate2271(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2272(.a(s_246), .O(gate424inter3));
  inv1  gate2273(.a(s_247), .O(gate424inter4));
  nand2 gate2274(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2275(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2276(.a(G1042), .O(gate424inter7));
  inv1  gate2277(.a(G1138), .O(gate424inter8));
  nand2 gate2278(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2279(.a(s_247), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2280(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2281(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2282(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate3039(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate3040(.a(gate426inter0), .b(s_356), .O(gate426inter1));
  and2  gate3041(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate3042(.a(s_356), .O(gate426inter3));
  inv1  gate3043(.a(s_357), .O(gate426inter4));
  nand2 gate3044(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate3045(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate3046(.a(G1045), .O(gate426inter7));
  inv1  gate3047(.a(G1141), .O(gate426inter8));
  nand2 gate3048(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate3049(.a(s_357), .b(gate426inter3), .O(gate426inter10));
  nor2  gate3050(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate3051(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate3052(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1737(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1738(.a(gate427inter0), .b(s_170), .O(gate427inter1));
  and2  gate1739(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1740(.a(s_170), .O(gate427inter3));
  inv1  gate1741(.a(s_171), .O(gate427inter4));
  nand2 gate1742(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1743(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1744(.a(G5), .O(gate427inter7));
  inv1  gate1745(.a(G1144), .O(gate427inter8));
  nand2 gate1746(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1747(.a(s_171), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1748(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1749(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1750(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1681(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1682(.a(gate428inter0), .b(s_162), .O(gate428inter1));
  and2  gate1683(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1684(.a(s_162), .O(gate428inter3));
  inv1  gate1685(.a(s_163), .O(gate428inter4));
  nand2 gate1686(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1687(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1688(.a(G1048), .O(gate428inter7));
  inv1  gate1689(.a(G1144), .O(gate428inter8));
  nand2 gate1690(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1691(.a(s_163), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1692(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1693(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1694(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate3081(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate3082(.a(gate432inter0), .b(s_362), .O(gate432inter1));
  and2  gate3083(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate3084(.a(s_362), .O(gate432inter3));
  inv1  gate3085(.a(s_363), .O(gate432inter4));
  nand2 gate3086(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate3087(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate3088(.a(G1054), .O(gate432inter7));
  inv1  gate3089(.a(G1150), .O(gate432inter8));
  nand2 gate3090(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate3091(.a(s_363), .b(gate432inter3), .O(gate432inter10));
  nor2  gate3092(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate3093(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate3094(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1177(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1178(.a(gate435inter0), .b(s_90), .O(gate435inter1));
  and2  gate1179(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1180(.a(s_90), .O(gate435inter3));
  inv1  gate1181(.a(s_91), .O(gate435inter4));
  nand2 gate1182(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1183(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1184(.a(G9), .O(gate435inter7));
  inv1  gate1185(.a(G1156), .O(gate435inter8));
  nand2 gate1186(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1187(.a(s_91), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1188(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1189(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1190(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2493(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2494(.a(gate438inter0), .b(s_278), .O(gate438inter1));
  and2  gate2495(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2496(.a(s_278), .O(gate438inter3));
  inv1  gate2497(.a(s_279), .O(gate438inter4));
  nand2 gate2498(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2499(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2500(.a(G1063), .O(gate438inter7));
  inv1  gate2501(.a(G1159), .O(gate438inter8));
  nand2 gate2502(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2503(.a(s_279), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2504(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2505(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2506(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate3221(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate3222(.a(gate440inter0), .b(s_382), .O(gate440inter1));
  and2  gate3223(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate3224(.a(s_382), .O(gate440inter3));
  inv1  gate3225(.a(s_383), .O(gate440inter4));
  nand2 gate3226(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate3227(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate3228(.a(G1066), .O(gate440inter7));
  inv1  gate3229(.a(G1162), .O(gate440inter8));
  nand2 gate3230(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate3231(.a(s_383), .b(gate440inter3), .O(gate440inter10));
  nor2  gate3232(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate3233(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate3234(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate799(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate800(.a(gate442inter0), .b(s_36), .O(gate442inter1));
  and2  gate801(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate802(.a(s_36), .O(gate442inter3));
  inv1  gate803(.a(s_37), .O(gate442inter4));
  nand2 gate804(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate805(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate806(.a(G1069), .O(gate442inter7));
  inv1  gate807(.a(G1165), .O(gate442inter8));
  nand2 gate808(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate809(.a(s_37), .b(gate442inter3), .O(gate442inter10));
  nor2  gate810(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate811(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate812(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1779(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1780(.a(gate444inter0), .b(s_176), .O(gate444inter1));
  and2  gate1781(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1782(.a(s_176), .O(gate444inter3));
  inv1  gate1783(.a(s_177), .O(gate444inter4));
  nand2 gate1784(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1785(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1786(.a(G1072), .O(gate444inter7));
  inv1  gate1787(.a(G1168), .O(gate444inter8));
  nand2 gate1788(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1789(.a(s_177), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1790(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1791(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1792(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate2171(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2172(.a(gate445inter0), .b(s_232), .O(gate445inter1));
  and2  gate2173(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2174(.a(s_232), .O(gate445inter3));
  inv1  gate2175(.a(s_233), .O(gate445inter4));
  nand2 gate2176(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2177(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2178(.a(G14), .O(gate445inter7));
  inv1  gate2179(.a(G1171), .O(gate445inter8));
  nand2 gate2180(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2181(.a(s_233), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2182(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2183(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2184(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2759(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2760(.a(gate448inter0), .b(s_316), .O(gate448inter1));
  and2  gate2761(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2762(.a(s_316), .O(gate448inter3));
  inv1  gate2763(.a(s_317), .O(gate448inter4));
  nand2 gate2764(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2765(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2766(.a(G1078), .O(gate448inter7));
  inv1  gate2767(.a(G1174), .O(gate448inter8));
  nand2 gate2768(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2769(.a(s_317), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2770(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2771(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2772(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2633(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2634(.a(gate449inter0), .b(s_298), .O(gate449inter1));
  and2  gate2635(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2636(.a(s_298), .O(gate449inter3));
  inv1  gate2637(.a(s_299), .O(gate449inter4));
  nand2 gate2638(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2639(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2640(.a(G16), .O(gate449inter7));
  inv1  gate2641(.a(G1177), .O(gate449inter8));
  nand2 gate2642(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2643(.a(s_299), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2644(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2645(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2646(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1191(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1192(.a(gate452inter0), .b(s_92), .O(gate452inter1));
  and2  gate1193(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1194(.a(s_92), .O(gate452inter3));
  inv1  gate1195(.a(s_93), .O(gate452inter4));
  nand2 gate1196(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1197(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1198(.a(G1084), .O(gate452inter7));
  inv1  gate1199(.a(G1180), .O(gate452inter8));
  nand2 gate1200(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1201(.a(s_93), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1202(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1203(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1204(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate981(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate982(.a(gate454inter0), .b(s_62), .O(gate454inter1));
  and2  gate983(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate984(.a(s_62), .O(gate454inter3));
  inv1  gate985(.a(s_63), .O(gate454inter4));
  nand2 gate986(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate987(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate988(.a(G1087), .O(gate454inter7));
  inv1  gate989(.a(G1183), .O(gate454inter8));
  nand2 gate990(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate991(.a(s_63), .b(gate454inter3), .O(gate454inter10));
  nor2  gate992(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate993(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate994(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1387(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1388(.a(gate456inter0), .b(s_120), .O(gate456inter1));
  and2  gate1389(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1390(.a(s_120), .O(gate456inter3));
  inv1  gate1391(.a(s_121), .O(gate456inter4));
  nand2 gate1392(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1393(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1394(.a(G1090), .O(gate456inter7));
  inv1  gate1395(.a(G1186), .O(gate456inter8));
  nand2 gate1396(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1397(.a(s_121), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1398(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1399(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1400(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2703(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2704(.a(gate458inter0), .b(s_308), .O(gate458inter1));
  and2  gate2705(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2706(.a(s_308), .O(gate458inter3));
  inv1  gate2707(.a(s_309), .O(gate458inter4));
  nand2 gate2708(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2709(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2710(.a(G1093), .O(gate458inter7));
  inv1  gate2711(.a(G1189), .O(gate458inter8));
  nand2 gate2712(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2713(.a(s_309), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2714(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2715(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2716(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate3137(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate3138(.a(gate459inter0), .b(s_370), .O(gate459inter1));
  and2  gate3139(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate3140(.a(s_370), .O(gate459inter3));
  inv1  gate3141(.a(s_371), .O(gate459inter4));
  nand2 gate3142(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate3143(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate3144(.a(G21), .O(gate459inter7));
  inv1  gate3145(.a(G1192), .O(gate459inter8));
  nand2 gate3146(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate3147(.a(s_371), .b(gate459inter3), .O(gate459inter10));
  nor2  gate3148(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate3149(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate3150(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2843(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2844(.a(gate461inter0), .b(s_328), .O(gate461inter1));
  and2  gate2845(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2846(.a(s_328), .O(gate461inter3));
  inv1  gate2847(.a(s_329), .O(gate461inter4));
  nand2 gate2848(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2849(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2850(.a(G22), .O(gate461inter7));
  inv1  gate2851(.a(G1195), .O(gate461inter8));
  nand2 gate2852(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2853(.a(s_329), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2854(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2855(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2856(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2731(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2732(.a(gate462inter0), .b(s_312), .O(gate462inter1));
  and2  gate2733(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2734(.a(s_312), .O(gate462inter3));
  inv1  gate2735(.a(s_313), .O(gate462inter4));
  nand2 gate2736(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2737(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2738(.a(G1099), .O(gate462inter7));
  inv1  gate2739(.a(G1195), .O(gate462inter8));
  nand2 gate2740(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2741(.a(s_313), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2742(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2743(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2744(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2185(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2186(.a(gate463inter0), .b(s_234), .O(gate463inter1));
  and2  gate2187(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2188(.a(s_234), .O(gate463inter3));
  inv1  gate2189(.a(s_235), .O(gate463inter4));
  nand2 gate2190(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2191(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2192(.a(G23), .O(gate463inter7));
  inv1  gate2193(.a(G1198), .O(gate463inter8));
  nand2 gate2194(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2195(.a(s_235), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2196(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2197(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2198(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2955(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2956(.a(gate465inter0), .b(s_344), .O(gate465inter1));
  and2  gate2957(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2958(.a(s_344), .O(gate465inter3));
  inv1  gate2959(.a(s_345), .O(gate465inter4));
  nand2 gate2960(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2961(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2962(.a(G24), .O(gate465inter7));
  inv1  gate2963(.a(G1201), .O(gate465inter8));
  nand2 gate2964(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2965(.a(s_345), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2966(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2967(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2968(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1695(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1696(.a(gate466inter0), .b(s_164), .O(gate466inter1));
  and2  gate1697(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1698(.a(s_164), .O(gate466inter3));
  inv1  gate1699(.a(s_165), .O(gate466inter4));
  nand2 gate1700(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1701(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1702(.a(G1105), .O(gate466inter7));
  inv1  gate1703(.a(G1201), .O(gate466inter8));
  nand2 gate1704(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1705(.a(s_165), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1706(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1707(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1708(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2675(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2676(.a(gate470inter0), .b(s_304), .O(gate470inter1));
  and2  gate2677(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2678(.a(s_304), .O(gate470inter3));
  inv1  gate2679(.a(s_305), .O(gate470inter4));
  nand2 gate2680(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2681(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2682(.a(G1111), .O(gate470inter7));
  inv1  gate2683(.a(G1207), .O(gate470inter8));
  nand2 gate2684(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2685(.a(s_305), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2686(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2687(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2688(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2059(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2060(.a(gate471inter0), .b(s_216), .O(gate471inter1));
  and2  gate2061(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2062(.a(s_216), .O(gate471inter3));
  inv1  gate2063(.a(s_217), .O(gate471inter4));
  nand2 gate2064(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2065(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2066(.a(G27), .O(gate471inter7));
  inv1  gate2067(.a(G1210), .O(gate471inter8));
  nand2 gate2068(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2069(.a(s_217), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2070(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2071(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2072(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2647(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2648(.a(gate474inter0), .b(s_300), .O(gate474inter1));
  and2  gate2649(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2650(.a(s_300), .O(gate474inter3));
  inv1  gate2651(.a(s_301), .O(gate474inter4));
  nand2 gate2652(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2653(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2654(.a(G1117), .O(gate474inter7));
  inv1  gate2655(.a(G1213), .O(gate474inter8));
  nand2 gate2656(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2657(.a(s_301), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2658(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2659(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2660(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2997(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2998(.a(gate476inter0), .b(s_350), .O(gate476inter1));
  and2  gate2999(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate3000(.a(s_350), .O(gate476inter3));
  inv1  gate3001(.a(s_351), .O(gate476inter4));
  nand2 gate3002(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate3003(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate3004(.a(G1120), .O(gate476inter7));
  inv1  gate3005(.a(G1216), .O(gate476inter8));
  nand2 gate3006(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate3007(.a(s_351), .b(gate476inter3), .O(gate476inter10));
  nor2  gate3008(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate3009(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate3010(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1807(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1808(.a(gate478inter0), .b(s_180), .O(gate478inter1));
  and2  gate1809(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1810(.a(s_180), .O(gate478inter3));
  inv1  gate1811(.a(s_181), .O(gate478inter4));
  nand2 gate1812(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1813(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1814(.a(G1123), .O(gate478inter7));
  inv1  gate1815(.a(G1219), .O(gate478inter8));
  nand2 gate1816(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1817(.a(s_181), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1818(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1819(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1820(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate2983(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2984(.a(gate481inter0), .b(s_348), .O(gate481inter1));
  and2  gate2985(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2986(.a(s_348), .O(gate481inter3));
  inv1  gate2987(.a(s_349), .O(gate481inter4));
  nand2 gate2988(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2989(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2990(.a(G32), .O(gate481inter7));
  inv1  gate2991(.a(G1225), .O(gate481inter8));
  nand2 gate2992(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2993(.a(s_349), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2994(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2995(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2996(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1093(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1094(.a(gate482inter0), .b(s_78), .O(gate482inter1));
  and2  gate1095(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1096(.a(s_78), .O(gate482inter3));
  inv1  gate1097(.a(s_79), .O(gate482inter4));
  nand2 gate1098(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1099(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1100(.a(G1129), .O(gate482inter7));
  inv1  gate1101(.a(G1225), .O(gate482inter8));
  nand2 gate1102(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1103(.a(s_79), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1104(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1105(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1106(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1121(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1122(.a(gate484inter0), .b(s_82), .O(gate484inter1));
  and2  gate1123(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1124(.a(s_82), .O(gate484inter3));
  inv1  gate1125(.a(s_83), .O(gate484inter4));
  nand2 gate1126(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1127(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1128(.a(G1230), .O(gate484inter7));
  inv1  gate1129(.a(G1231), .O(gate484inter8));
  nand2 gate1130(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1131(.a(s_83), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1132(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1133(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1134(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2661(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2662(.a(gate485inter0), .b(s_302), .O(gate485inter1));
  and2  gate2663(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2664(.a(s_302), .O(gate485inter3));
  inv1  gate2665(.a(s_303), .O(gate485inter4));
  nand2 gate2666(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2667(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2668(.a(G1232), .O(gate485inter7));
  inv1  gate2669(.a(G1233), .O(gate485inter8));
  nand2 gate2670(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2671(.a(s_303), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2672(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2673(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2674(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate911(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate912(.a(gate489inter0), .b(s_52), .O(gate489inter1));
  and2  gate913(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate914(.a(s_52), .O(gate489inter3));
  inv1  gate915(.a(s_53), .O(gate489inter4));
  nand2 gate916(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate917(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate918(.a(G1240), .O(gate489inter7));
  inv1  gate919(.a(G1241), .O(gate489inter8));
  nand2 gate920(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate921(.a(s_53), .b(gate489inter3), .O(gate489inter10));
  nor2  gate922(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate923(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate924(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate869(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate870(.a(gate491inter0), .b(s_46), .O(gate491inter1));
  and2  gate871(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate872(.a(s_46), .O(gate491inter3));
  inv1  gate873(.a(s_47), .O(gate491inter4));
  nand2 gate874(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate875(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate876(.a(G1244), .O(gate491inter7));
  inv1  gate877(.a(G1245), .O(gate491inter8));
  nand2 gate878(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate879(.a(s_47), .b(gate491inter3), .O(gate491inter10));
  nor2  gate880(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate881(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate882(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2087(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2088(.a(gate493inter0), .b(s_220), .O(gate493inter1));
  and2  gate2089(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2090(.a(s_220), .O(gate493inter3));
  inv1  gate2091(.a(s_221), .O(gate493inter4));
  nand2 gate2092(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2093(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2094(.a(G1248), .O(gate493inter7));
  inv1  gate2095(.a(G1249), .O(gate493inter8));
  nand2 gate2096(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2097(.a(s_221), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2098(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2099(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2100(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1485(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1486(.a(gate494inter0), .b(s_134), .O(gate494inter1));
  and2  gate1487(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1488(.a(s_134), .O(gate494inter3));
  inv1  gate1489(.a(s_135), .O(gate494inter4));
  nand2 gate1490(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1491(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1492(.a(G1250), .O(gate494inter7));
  inv1  gate1493(.a(G1251), .O(gate494inter8));
  nand2 gate1494(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1495(.a(s_135), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1496(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1497(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1498(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1905(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1906(.a(gate495inter0), .b(s_194), .O(gate495inter1));
  and2  gate1907(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1908(.a(s_194), .O(gate495inter3));
  inv1  gate1909(.a(s_195), .O(gate495inter4));
  nand2 gate1910(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1911(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1912(.a(G1252), .O(gate495inter7));
  inv1  gate1913(.a(G1253), .O(gate495inter8));
  nand2 gate1914(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1915(.a(s_195), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1916(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1917(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1918(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate757(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate758(.a(gate497inter0), .b(s_30), .O(gate497inter1));
  and2  gate759(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate760(.a(s_30), .O(gate497inter3));
  inv1  gate761(.a(s_31), .O(gate497inter4));
  nand2 gate762(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate763(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate764(.a(G1256), .O(gate497inter7));
  inv1  gate765(.a(G1257), .O(gate497inter8));
  nand2 gate766(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate767(.a(s_31), .b(gate497inter3), .O(gate497inter10));
  nor2  gate768(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate769(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate770(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1765(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1766(.a(gate500inter0), .b(s_174), .O(gate500inter1));
  and2  gate1767(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1768(.a(s_174), .O(gate500inter3));
  inv1  gate1769(.a(s_175), .O(gate500inter4));
  nand2 gate1770(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1771(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1772(.a(G1262), .O(gate500inter7));
  inv1  gate1773(.a(G1263), .O(gate500inter8));
  nand2 gate1774(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1775(.a(s_175), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1776(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1777(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1778(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2563(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2564(.a(gate501inter0), .b(s_288), .O(gate501inter1));
  and2  gate2565(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2566(.a(s_288), .O(gate501inter3));
  inv1  gate2567(.a(s_289), .O(gate501inter4));
  nand2 gate2568(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2569(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2570(.a(G1264), .O(gate501inter7));
  inv1  gate2571(.a(G1265), .O(gate501inter8));
  nand2 gate2572(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2573(.a(s_289), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2574(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2575(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2576(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1541(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1542(.a(gate503inter0), .b(s_142), .O(gate503inter1));
  and2  gate1543(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1544(.a(s_142), .O(gate503inter3));
  inv1  gate1545(.a(s_143), .O(gate503inter4));
  nand2 gate1546(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1547(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1548(.a(G1268), .O(gate503inter7));
  inv1  gate1549(.a(G1269), .O(gate503inter8));
  nand2 gate1550(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1551(.a(s_143), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1552(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1553(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1554(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1345(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1346(.a(gate505inter0), .b(s_114), .O(gate505inter1));
  and2  gate1347(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1348(.a(s_114), .O(gate505inter3));
  inv1  gate1349(.a(s_115), .O(gate505inter4));
  nand2 gate1350(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1351(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1352(.a(G1272), .O(gate505inter7));
  inv1  gate1353(.a(G1273), .O(gate505inter8));
  nand2 gate1354(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1355(.a(s_115), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1356(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1357(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1358(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1835(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1836(.a(gate508inter0), .b(s_184), .O(gate508inter1));
  and2  gate1837(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1838(.a(s_184), .O(gate508inter3));
  inv1  gate1839(.a(s_185), .O(gate508inter4));
  nand2 gate1840(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1841(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1842(.a(G1278), .O(gate508inter7));
  inv1  gate1843(.a(G1279), .O(gate508inter8));
  nand2 gate1844(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1845(.a(s_185), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1846(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1847(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1848(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2801(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2802(.a(gate509inter0), .b(s_322), .O(gate509inter1));
  and2  gate2803(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2804(.a(s_322), .O(gate509inter3));
  inv1  gate2805(.a(s_323), .O(gate509inter4));
  nand2 gate2806(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2807(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2808(.a(G1280), .O(gate509inter7));
  inv1  gate2809(.a(G1281), .O(gate509inter8));
  nand2 gate2810(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2811(.a(s_323), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2812(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2813(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2814(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1219(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1220(.a(gate510inter0), .b(s_96), .O(gate510inter1));
  and2  gate1221(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1222(.a(s_96), .O(gate510inter3));
  inv1  gate1223(.a(s_97), .O(gate510inter4));
  nand2 gate1224(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1225(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1226(.a(G1282), .O(gate510inter7));
  inv1  gate1227(.a(G1283), .O(gate510inter8));
  nand2 gate1228(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1229(.a(s_97), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1230(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1231(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1232(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate715(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate716(.a(gate511inter0), .b(s_24), .O(gate511inter1));
  and2  gate717(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate718(.a(s_24), .O(gate511inter3));
  inv1  gate719(.a(s_25), .O(gate511inter4));
  nand2 gate720(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate721(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate722(.a(G1284), .O(gate511inter7));
  inv1  gate723(.a(G1285), .O(gate511inter8));
  nand2 gate724(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate725(.a(s_25), .b(gate511inter3), .O(gate511inter10));
  nor2  gate726(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate727(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate728(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1947(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1948(.a(gate512inter0), .b(s_200), .O(gate512inter1));
  and2  gate1949(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1950(.a(s_200), .O(gate512inter3));
  inv1  gate1951(.a(s_201), .O(gate512inter4));
  nand2 gate1952(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1953(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1954(.a(G1286), .O(gate512inter7));
  inv1  gate1955(.a(G1287), .O(gate512inter8));
  nand2 gate1956(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1957(.a(s_201), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1958(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1959(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1960(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate547(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate548(.a(gate513inter0), .b(s_0), .O(gate513inter1));
  and2  gate549(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate550(.a(s_0), .O(gate513inter3));
  inv1  gate551(.a(s_1), .O(gate513inter4));
  nand2 gate552(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate553(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate554(.a(G1288), .O(gate513inter7));
  inv1  gate555(.a(G1289), .O(gate513inter8));
  nand2 gate556(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate557(.a(s_1), .b(gate513inter3), .O(gate513inter10));
  nor2  gate558(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate559(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate560(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule