module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
input s_382,s_383;//RE__ALLOW(00,01,10,11);
input s_384,s_385;//RE__ALLOW(00,01,10,11);
input s_386,s_387;//RE__ALLOW(00,01,10,11);
input s_388,s_389;//RE__ALLOW(00,01,10,11);
input s_390,s_391;//RE__ALLOW(00,01,10,11);
input s_392,s_393;//RE__ALLOW(00,01,10,11);
input s_394,s_395;//RE__ALLOW(00,01,10,11);
input s_396,s_397;//RE__ALLOW(00,01,10,11);
input s_398,s_399;//RE__ALLOW(00,01,10,11);
input s_400,s_401;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1331(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1332(.a(gate9inter0), .b(s_112), .O(gate9inter1));
  and2  gate1333(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1334(.a(s_112), .O(gate9inter3));
  inv1  gate1335(.a(s_113), .O(gate9inter4));
  nand2 gate1336(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1337(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1338(.a(G1), .O(gate9inter7));
  inv1  gate1339(.a(G2), .O(gate9inter8));
  nand2 gate1340(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1341(.a(s_113), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1342(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1343(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1344(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2773(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2774(.a(gate12inter0), .b(s_318), .O(gate12inter1));
  and2  gate2775(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2776(.a(s_318), .O(gate12inter3));
  inv1  gate2777(.a(s_319), .O(gate12inter4));
  nand2 gate2778(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2779(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2780(.a(G7), .O(gate12inter7));
  inv1  gate2781(.a(G8), .O(gate12inter8));
  nand2 gate2782(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2783(.a(s_319), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2784(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2785(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2786(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1135(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1136(.a(gate15inter0), .b(s_84), .O(gate15inter1));
  and2  gate1137(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1138(.a(s_84), .O(gate15inter3));
  inv1  gate1139(.a(s_85), .O(gate15inter4));
  nand2 gate1140(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1141(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1142(.a(G13), .O(gate15inter7));
  inv1  gate1143(.a(G14), .O(gate15inter8));
  nand2 gate1144(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1145(.a(s_85), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1146(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1147(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1148(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2633(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2634(.a(gate21inter0), .b(s_298), .O(gate21inter1));
  and2  gate2635(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2636(.a(s_298), .O(gate21inter3));
  inv1  gate2637(.a(s_299), .O(gate21inter4));
  nand2 gate2638(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2639(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2640(.a(G25), .O(gate21inter7));
  inv1  gate2641(.a(G26), .O(gate21inter8));
  nand2 gate2642(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2643(.a(s_299), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2644(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2645(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2646(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2787(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2788(.a(gate22inter0), .b(s_320), .O(gate22inter1));
  and2  gate2789(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2790(.a(s_320), .O(gate22inter3));
  inv1  gate2791(.a(s_321), .O(gate22inter4));
  nand2 gate2792(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2793(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2794(.a(G27), .O(gate22inter7));
  inv1  gate2795(.a(G28), .O(gate22inter8));
  nand2 gate2796(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2797(.a(s_321), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2798(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2799(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2800(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1919(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1920(.a(gate23inter0), .b(s_196), .O(gate23inter1));
  and2  gate1921(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1922(.a(s_196), .O(gate23inter3));
  inv1  gate1923(.a(s_197), .O(gate23inter4));
  nand2 gate1924(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1925(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1926(.a(G29), .O(gate23inter7));
  inv1  gate1927(.a(G30), .O(gate23inter8));
  nand2 gate1928(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1929(.a(s_197), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1930(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1931(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1932(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate3319(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate3320(.a(gate24inter0), .b(s_396), .O(gate24inter1));
  and2  gate3321(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate3322(.a(s_396), .O(gate24inter3));
  inv1  gate3323(.a(s_397), .O(gate24inter4));
  nand2 gate3324(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate3325(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate3326(.a(G31), .O(gate24inter7));
  inv1  gate3327(.a(G32), .O(gate24inter8));
  nand2 gate3328(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate3329(.a(s_397), .b(gate24inter3), .O(gate24inter10));
  nor2  gate3330(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate3331(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate3332(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate561(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate562(.a(gate25inter0), .b(s_2), .O(gate25inter1));
  and2  gate563(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate564(.a(s_2), .O(gate25inter3));
  inv1  gate565(.a(s_3), .O(gate25inter4));
  nand2 gate566(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate567(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate568(.a(G1), .O(gate25inter7));
  inv1  gate569(.a(G5), .O(gate25inter8));
  nand2 gate570(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate571(.a(s_3), .b(gate25inter3), .O(gate25inter10));
  nor2  gate572(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate573(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate574(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2129(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2130(.a(gate27inter0), .b(s_226), .O(gate27inter1));
  and2  gate2131(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2132(.a(s_226), .O(gate27inter3));
  inv1  gate2133(.a(s_227), .O(gate27inter4));
  nand2 gate2134(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2135(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2136(.a(G2), .O(gate27inter7));
  inv1  gate2137(.a(G6), .O(gate27inter8));
  nand2 gate2138(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2139(.a(s_227), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2140(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2141(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2142(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate2227(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2228(.a(gate28inter0), .b(s_240), .O(gate28inter1));
  and2  gate2229(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2230(.a(s_240), .O(gate28inter3));
  inv1  gate2231(.a(s_241), .O(gate28inter4));
  nand2 gate2232(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2233(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2234(.a(G10), .O(gate28inter7));
  inv1  gate2235(.a(G14), .O(gate28inter8));
  nand2 gate2236(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2237(.a(s_241), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2238(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2239(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2240(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1079(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1080(.a(gate30inter0), .b(s_76), .O(gate30inter1));
  and2  gate1081(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1082(.a(s_76), .O(gate30inter3));
  inv1  gate1083(.a(s_77), .O(gate30inter4));
  nand2 gate1084(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1085(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1086(.a(G11), .O(gate30inter7));
  inv1  gate1087(.a(G15), .O(gate30inter8));
  nand2 gate1088(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1089(.a(s_77), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1090(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1091(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1092(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2087(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2088(.a(gate34inter0), .b(s_220), .O(gate34inter1));
  and2  gate2089(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2090(.a(s_220), .O(gate34inter3));
  inv1  gate2091(.a(s_221), .O(gate34inter4));
  nand2 gate2092(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2093(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2094(.a(G25), .O(gate34inter7));
  inv1  gate2095(.a(G29), .O(gate34inter8));
  nand2 gate2096(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2097(.a(s_221), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2098(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2099(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2100(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate575(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate576(.a(gate36inter0), .b(s_4), .O(gate36inter1));
  and2  gate577(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate578(.a(s_4), .O(gate36inter3));
  inv1  gate579(.a(s_5), .O(gate36inter4));
  nand2 gate580(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate581(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate582(.a(G26), .O(gate36inter7));
  inv1  gate583(.a(G30), .O(gate36inter8));
  nand2 gate584(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate585(.a(s_5), .b(gate36inter3), .O(gate36inter10));
  nor2  gate586(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate587(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate588(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate2549(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2550(.a(gate37inter0), .b(s_286), .O(gate37inter1));
  and2  gate2551(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2552(.a(s_286), .O(gate37inter3));
  inv1  gate2553(.a(s_287), .O(gate37inter4));
  nand2 gate2554(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2555(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2556(.a(G19), .O(gate37inter7));
  inv1  gate2557(.a(G23), .O(gate37inter8));
  nand2 gate2558(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2559(.a(s_287), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2560(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2561(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2562(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate3053(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate3054(.a(gate39inter0), .b(s_358), .O(gate39inter1));
  and2  gate3055(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate3056(.a(s_358), .O(gate39inter3));
  inv1  gate3057(.a(s_359), .O(gate39inter4));
  nand2 gate3058(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate3059(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate3060(.a(G20), .O(gate39inter7));
  inv1  gate3061(.a(G24), .O(gate39inter8));
  nand2 gate3062(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate3063(.a(s_359), .b(gate39inter3), .O(gate39inter10));
  nor2  gate3064(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate3065(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate3066(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate2479(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2480(.a(gate40inter0), .b(s_276), .O(gate40inter1));
  and2  gate2481(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2482(.a(s_276), .O(gate40inter3));
  inv1  gate2483(.a(s_277), .O(gate40inter4));
  nand2 gate2484(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2485(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2486(.a(G28), .O(gate40inter7));
  inv1  gate2487(.a(G32), .O(gate40inter8));
  nand2 gate2488(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2489(.a(s_277), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2490(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2491(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2492(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2017(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2018(.a(gate41inter0), .b(s_210), .O(gate41inter1));
  and2  gate2019(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2020(.a(s_210), .O(gate41inter3));
  inv1  gate2021(.a(s_211), .O(gate41inter4));
  nand2 gate2022(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2023(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2024(.a(G1), .O(gate41inter7));
  inv1  gate2025(.a(G266), .O(gate41inter8));
  nand2 gate2026(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2027(.a(s_211), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2028(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2029(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2030(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2591(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2592(.a(gate44inter0), .b(s_292), .O(gate44inter1));
  and2  gate2593(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2594(.a(s_292), .O(gate44inter3));
  inv1  gate2595(.a(s_293), .O(gate44inter4));
  nand2 gate2596(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2597(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2598(.a(G4), .O(gate44inter7));
  inv1  gate2599(.a(G269), .O(gate44inter8));
  nand2 gate2600(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2601(.a(s_293), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2602(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2603(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2604(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1513(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1514(.a(gate46inter0), .b(s_138), .O(gate46inter1));
  and2  gate1515(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1516(.a(s_138), .O(gate46inter3));
  inv1  gate1517(.a(s_139), .O(gate46inter4));
  nand2 gate1518(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1519(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1520(.a(G6), .O(gate46inter7));
  inv1  gate1521(.a(G272), .O(gate46inter8));
  nand2 gate1522(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1523(.a(s_139), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1524(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1525(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1526(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1415(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1416(.a(gate50inter0), .b(s_124), .O(gate50inter1));
  and2  gate1417(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1418(.a(s_124), .O(gate50inter3));
  inv1  gate1419(.a(s_125), .O(gate50inter4));
  nand2 gate1420(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1421(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1422(.a(G10), .O(gate50inter7));
  inv1  gate1423(.a(G278), .O(gate50inter8));
  nand2 gate1424(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1425(.a(s_125), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1426(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1427(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1428(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate883(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate884(.a(gate51inter0), .b(s_48), .O(gate51inter1));
  and2  gate885(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate886(.a(s_48), .O(gate51inter3));
  inv1  gate887(.a(s_49), .O(gate51inter4));
  nand2 gate888(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate889(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate890(.a(G11), .O(gate51inter7));
  inv1  gate891(.a(G281), .O(gate51inter8));
  nand2 gate892(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate893(.a(s_49), .b(gate51inter3), .O(gate51inter10));
  nor2  gate894(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate895(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate896(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1905(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1906(.a(gate53inter0), .b(s_194), .O(gate53inter1));
  and2  gate1907(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1908(.a(s_194), .O(gate53inter3));
  inv1  gate1909(.a(s_195), .O(gate53inter4));
  nand2 gate1910(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1911(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1912(.a(G13), .O(gate53inter7));
  inv1  gate1913(.a(G284), .O(gate53inter8));
  nand2 gate1914(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1915(.a(s_195), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1916(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1917(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1918(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate2185(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2186(.a(gate54inter0), .b(s_234), .O(gate54inter1));
  and2  gate2187(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2188(.a(s_234), .O(gate54inter3));
  inv1  gate2189(.a(s_235), .O(gate54inter4));
  nand2 gate2190(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2191(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2192(.a(G14), .O(gate54inter7));
  inv1  gate2193(.a(G284), .O(gate54inter8));
  nand2 gate2194(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2195(.a(s_235), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2196(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2197(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2198(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2899(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2900(.a(gate61inter0), .b(s_336), .O(gate61inter1));
  and2  gate2901(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2902(.a(s_336), .O(gate61inter3));
  inv1  gate2903(.a(s_337), .O(gate61inter4));
  nand2 gate2904(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2905(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2906(.a(G21), .O(gate61inter7));
  inv1  gate2907(.a(G296), .O(gate61inter8));
  nand2 gate2908(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2909(.a(s_337), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2910(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2911(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2912(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate2073(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2074(.a(gate63inter0), .b(s_218), .O(gate63inter1));
  and2  gate2075(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2076(.a(s_218), .O(gate63inter3));
  inv1  gate2077(.a(s_219), .O(gate63inter4));
  nand2 gate2078(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2079(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2080(.a(G23), .O(gate63inter7));
  inv1  gate2081(.a(G299), .O(gate63inter8));
  nand2 gate2082(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2083(.a(s_219), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2084(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2085(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2086(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2969(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2970(.a(gate68inter0), .b(s_346), .O(gate68inter1));
  and2  gate2971(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2972(.a(s_346), .O(gate68inter3));
  inv1  gate2973(.a(s_347), .O(gate68inter4));
  nand2 gate2974(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2975(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2976(.a(G28), .O(gate68inter7));
  inv1  gate2977(.a(G305), .O(gate68inter8));
  nand2 gate2978(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2979(.a(s_347), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2980(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2981(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2982(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate2409(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2410(.a(gate69inter0), .b(s_266), .O(gate69inter1));
  and2  gate2411(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2412(.a(s_266), .O(gate69inter3));
  inv1  gate2413(.a(s_267), .O(gate69inter4));
  nand2 gate2414(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2415(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2416(.a(G29), .O(gate69inter7));
  inv1  gate2417(.a(G308), .O(gate69inter8));
  nand2 gate2418(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2419(.a(s_267), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2420(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2421(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2422(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2269(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2270(.a(gate70inter0), .b(s_246), .O(gate70inter1));
  and2  gate2271(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2272(.a(s_246), .O(gate70inter3));
  inv1  gate2273(.a(s_247), .O(gate70inter4));
  nand2 gate2274(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2275(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2276(.a(G30), .O(gate70inter7));
  inv1  gate2277(.a(G308), .O(gate70inter8));
  nand2 gate2278(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2279(.a(s_247), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2280(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2281(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2282(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate3221(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate3222(.a(gate72inter0), .b(s_382), .O(gate72inter1));
  and2  gate3223(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate3224(.a(s_382), .O(gate72inter3));
  inv1  gate3225(.a(s_383), .O(gate72inter4));
  nand2 gate3226(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate3227(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate3228(.a(G32), .O(gate72inter7));
  inv1  gate3229(.a(G311), .O(gate72inter8));
  nand2 gate3230(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate3231(.a(s_383), .b(gate72inter3), .O(gate72inter10));
  nor2  gate3232(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate3233(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate3234(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1989(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1990(.a(gate73inter0), .b(s_206), .O(gate73inter1));
  and2  gate1991(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1992(.a(s_206), .O(gate73inter3));
  inv1  gate1993(.a(s_207), .O(gate73inter4));
  nand2 gate1994(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1995(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1996(.a(G1), .O(gate73inter7));
  inv1  gate1997(.a(G314), .O(gate73inter8));
  nand2 gate1998(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1999(.a(s_207), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2000(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2001(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2002(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate3123(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate3124(.a(gate74inter0), .b(s_368), .O(gate74inter1));
  and2  gate3125(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate3126(.a(s_368), .O(gate74inter3));
  inv1  gate3127(.a(s_369), .O(gate74inter4));
  nand2 gate3128(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate3129(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate3130(.a(G5), .O(gate74inter7));
  inv1  gate3131(.a(G314), .O(gate74inter8));
  nand2 gate3132(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate3133(.a(s_369), .b(gate74inter3), .O(gate74inter10));
  nor2  gate3134(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate3135(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate3136(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1009(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1010(.a(gate75inter0), .b(s_66), .O(gate75inter1));
  and2  gate1011(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1012(.a(s_66), .O(gate75inter3));
  inv1  gate1013(.a(s_67), .O(gate75inter4));
  nand2 gate1014(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1015(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1016(.a(G9), .O(gate75inter7));
  inv1  gate1017(.a(G317), .O(gate75inter8));
  nand2 gate1018(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1019(.a(s_67), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1020(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1021(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1022(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1807(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1808(.a(gate81inter0), .b(s_180), .O(gate81inter1));
  and2  gate1809(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1810(.a(s_180), .O(gate81inter3));
  inv1  gate1811(.a(s_181), .O(gate81inter4));
  nand2 gate1812(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1813(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1814(.a(G3), .O(gate81inter7));
  inv1  gate1815(.a(G326), .O(gate81inter8));
  nand2 gate1816(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1817(.a(s_181), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1818(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1819(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1820(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1345(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1346(.a(gate82inter0), .b(s_114), .O(gate82inter1));
  and2  gate1347(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1348(.a(s_114), .O(gate82inter3));
  inv1  gate1349(.a(s_115), .O(gate82inter4));
  nand2 gate1350(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1351(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1352(.a(G7), .O(gate82inter7));
  inv1  gate1353(.a(G326), .O(gate82inter8));
  nand2 gate1354(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1355(.a(s_115), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1356(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1357(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1358(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2493(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2494(.a(gate85inter0), .b(s_278), .O(gate85inter1));
  and2  gate2495(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2496(.a(s_278), .O(gate85inter3));
  inv1  gate2497(.a(s_279), .O(gate85inter4));
  nand2 gate2498(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2499(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2500(.a(G4), .O(gate85inter7));
  inv1  gate2501(.a(G332), .O(gate85inter8));
  nand2 gate2502(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2503(.a(s_279), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2504(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2505(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2506(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1751(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1752(.a(gate87inter0), .b(s_172), .O(gate87inter1));
  and2  gate1753(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1754(.a(s_172), .O(gate87inter3));
  inv1  gate1755(.a(s_173), .O(gate87inter4));
  nand2 gate1756(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1757(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1758(.a(G12), .O(gate87inter7));
  inv1  gate1759(.a(G335), .O(gate87inter8));
  nand2 gate1760(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1761(.a(s_173), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1762(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1763(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1764(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate743(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate744(.a(gate90inter0), .b(s_28), .O(gate90inter1));
  and2  gate745(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate746(.a(s_28), .O(gate90inter3));
  inv1  gate747(.a(s_29), .O(gate90inter4));
  nand2 gate748(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate749(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate750(.a(G21), .O(gate90inter7));
  inv1  gate751(.a(G338), .O(gate90inter8));
  nand2 gate752(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate753(.a(s_29), .b(gate90inter3), .O(gate90inter10));
  nor2  gate754(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate755(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate756(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2059(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2060(.a(gate92inter0), .b(s_216), .O(gate92inter1));
  and2  gate2061(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2062(.a(s_216), .O(gate92inter3));
  inv1  gate2063(.a(s_217), .O(gate92inter4));
  nand2 gate2064(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2065(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2066(.a(G29), .O(gate92inter7));
  inv1  gate2067(.a(G341), .O(gate92inter8));
  nand2 gate2068(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2069(.a(s_217), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2070(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2071(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2072(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate673(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate674(.a(gate94inter0), .b(s_18), .O(gate94inter1));
  and2  gate675(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate676(.a(s_18), .O(gate94inter3));
  inv1  gate677(.a(s_19), .O(gate94inter4));
  nand2 gate678(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate679(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate680(.a(G22), .O(gate94inter7));
  inv1  gate681(.a(G344), .O(gate94inter8));
  nand2 gate682(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate683(.a(s_19), .b(gate94inter3), .O(gate94inter10));
  nor2  gate684(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate685(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate686(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2241(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2242(.a(gate96inter0), .b(s_242), .O(gate96inter1));
  and2  gate2243(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2244(.a(s_242), .O(gate96inter3));
  inv1  gate2245(.a(s_243), .O(gate96inter4));
  nand2 gate2246(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2247(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2248(.a(G30), .O(gate96inter7));
  inv1  gate2249(.a(G347), .O(gate96inter8));
  nand2 gate2250(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2251(.a(s_243), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2252(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2253(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2254(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1275(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1276(.a(gate98inter0), .b(s_104), .O(gate98inter1));
  and2  gate1277(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1278(.a(s_104), .O(gate98inter3));
  inv1  gate1279(.a(s_105), .O(gate98inter4));
  nand2 gate1280(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1281(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1282(.a(G23), .O(gate98inter7));
  inv1  gate1283(.a(G350), .O(gate98inter8));
  nand2 gate1284(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1285(.a(s_105), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1286(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1287(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1288(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2213(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2214(.a(gate99inter0), .b(s_238), .O(gate99inter1));
  and2  gate2215(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2216(.a(s_238), .O(gate99inter3));
  inv1  gate2217(.a(s_239), .O(gate99inter4));
  nand2 gate2218(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2219(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2220(.a(G27), .O(gate99inter7));
  inv1  gate2221(.a(G353), .O(gate99inter8));
  nand2 gate2222(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2223(.a(s_239), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2224(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2225(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2226(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate3067(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate3068(.a(gate100inter0), .b(s_360), .O(gate100inter1));
  and2  gate3069(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate3070(.a(s_360), .O(gate100inter3));
  inv1  gate3071(.a(s_361), .O(gate100inter4));
  nand2 gate3072(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate3073(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate3074(.a(G31), .O(gate100inter7));
  inv1  gate3075(.a(G353), .O(gate100inter8));
  nand2 gate3076(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate3077(.a(s_361), .b(gate100inter3), .O(gate100inter10));
  nor2  gate3078(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate3079(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate3080(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate2101(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2102(.a(gate101inter0), .b(s_222), .O(gate101inter1));
  and2  gate2103(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2104(.a(s_222), .O(gate101inter3));
  inv1  gate2105(.a(s_223), .O(gate101inter4));
  nand2 gate2106(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2107(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2108(.a(G20), .O(gate101inter7));
  inv1  gate2109(.a(G356), .O(gate101inter8));
  nand2 gate2110(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2111(.a(s_223), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2112(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2113(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2114(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2381(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2382(.a(gate102inter0), .b(s_262), .O(gate102inter1));
  and2  gate2383(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2384(.a(s_262), .O(gate102inter3));
  inv1  gate2385(.a(s_263), .O(gate102inter4));
  nand2 gate2386(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2387(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2388(.a(G24), .O(gate102inter7));
  inv1  gate2389(.a(G356), .O(gate102inter8));
  nand2 gate2390(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2391(.a(s_263), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2392(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2393(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2394(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate981(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate982(.a(gate103inter0), .b(s_62), .O(gate103inter1));
  and2  gate983(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate984(.a(s_62), .O(gate103inter3));
  inv1  gate985(.a(s_63), .O(gate103inter4));
  nand2 gate986(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate987(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate988(.a(G28), .O(gate103inter7));
  inv1  gate989(.a(G359), .O(gate103inter8));
  nand2 gate990(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate991(.a(s_63), .b(gate103inter3), .O(gate103inter10));
  nor2  gate992(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate993(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate994(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1541(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1542(.a(gate106inter0), .b(s_142), .O(gate106inter1));
  and2  gate1543(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1544(.a(s_142), .O(gate106inter3));
  inv1  gate1545(.a(s_143), .O(gate106inter4));
  nand2 gate1546(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1547(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1548(.a(G364), .O(gate106inter7));
  inv1  gate1549(.a(G365), .O(gate106inter8));
  nand2 gate1550(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1551(.a(s_143), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1552(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1553(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1554(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1303(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1304(.a(gate107inter0), .b(s_108), .O(gate107inter1));
  and2  gate1305(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1306(.a(s_108), .O(gate107inter3));
  inv1  gate1307(.a(s_109), .O(gate107inter4));
  nand2 gate1308(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1309(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1310(.a(G366), .O(gate107inter7));
  inv1  gate1311(.a(G367), .O(gate107inter8));
  nand2 gate1312(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1313(.a(s_109), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1314(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1315(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1316(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate3109(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate3110(.a(gate108inter0), .b(s_366), .O(gate108inter1));
  and2  gate3111(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate3112(.a(s_366), .O(gate108inter3));
  inv1  gate3113(.a(s_367), .O(gate108inter4));
  nand2 gate3114(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate3115(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate3116(.a(G368), .O(gate108inter7));
  inv1  gate3117(.a(G369), .O(gate108inter8));
  nand2 gate3118(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate3119(.a(s_367), .b(gate108inter3), .O(gate108inter10));
  nor2  gate3120(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate3121(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate3122(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2423(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2424(.a(gate112inter0), .b(s_268), .O(gate112inter1));
  and2  gate2425(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2426(.a(s_268), .O(gate112inter3));
  inv1  gate2427(.a(s_269), .O(gate112inter4));
  nand2 gate2428(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2429(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2430(.a(G376), .O(gate112inter7));
  inv1  gate2431(.a(G377), .O(gate112inter8));
  nand2 gate2432(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2433(.a(s_269), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2434(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2435(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2436(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2731(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2732(.a(gate116inter0), .b(s_312), .O(gate116inter1));
  and2  gate2733(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2734(.a(s_312), .O(gate116inter3));
  inv1  gate2735(.a(s_313), .O(gate116inter4));
  nand2 gate2736(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2737(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2738(.a(G384), .O(gate116inter7));
  inv1  gate2739(.a(G385), .O(gate116inter8));
  nand2 gate2740(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2741(.a(s_313), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2742(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2743(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2744(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1121(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1122(.a(gate118inter0), .b(s_82), .O(gate118inter1));
  and2  gate1123(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1124(.a(s_82), .O(gate118inter3));
  inv1  gate1125(.a(s_83), .O(gate118inter4));
  nand2 gate1126(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1127(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1128(.a(G388), .O(gate118inter7));
  inv1  gate1129(.a(G389), .O(gate118inter8));
  nand2 gate1130(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1131(.a(s_83), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1132(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1133(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1134(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1821(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1822(.a(gate119inter0), .b(s_182), .O(gate119inter1));
  and2  gate1823(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1824(.a(s_182), .O(gate119inter3));
  inv1  gate1825(.a(s_183), .O(gate119inter4));
  nand2 gate1826(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1827(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1828(.a(G390), .O(gate119inter7));
  inv1  gate1829(.a(G391), .O(gate119inter8));
  nand2 gate1830(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1831(.a(s_183), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1832(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1833(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1834(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate2661(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2662(.a(gate120inter0), .b(s_302), .O(gate120inter1));
  and2  gate2663(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2664(.a(s_302), .O(gate120inter3));
  inv1  gate2665(.a(s_303), .O(gate120inter4));
  nand2 gate2666(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2667(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2668(.a(G392), .O(gate120inter7));
  inv1  gate2669(.a(G393), .O(gate120inter8));
  nand2 gate2670(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2671(.a(s_303), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2672(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2673(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2674(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1163(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1164(.a(gate127inter0), .b(s_88), .O(gate127inter1));
  and2  gate1165(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1166(.a(s_88), .O(gate127inter3));
  inv1  gate1167(.a(s_89), .O(gate127inter4));
  nand2 gate1168(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1169(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1170(.a(G406), .O(gate127inter7));
  inv1  gate1171(.a(G407), .O(gate127inter8));
  nand2 gate1172(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1173(.a(s_89), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1174(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1175(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1176(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1779(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1780(.a(gate129inter0), .b(s_176), .O(gate129inter1));
  and2  gate1781(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1782(.a(s_176), .O(gate129inter3));
  inv1  gate1783(.a(s_177), .O(gate129inter4));
  nand2 gate1784(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1785(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1786(.a(G410), .O(gate129inter7));
  inv1  gate1787(.a(G411), .O(gate129inter8));
  nand2 gate1788(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1789(.a(s_177), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1790(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1791(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1792(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate1709(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1710(.a(gate130inter0), .b(s_166), .O(gate130inter1));
  and2  gate1711(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1712(.a(s_166), .O(gate130inter3));
  inv1  gate1713(.a(s_167), .O(gate130inter4));
  nand2 gate1714(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1715(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1716(.a(G412), .O(gate130inter7));
  inv1  gate1717(.a(G413), .O(gate130inter8));
  nand2 gate1718(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1719(.a(s_167), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1720(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1721(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1722(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2801(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2802(.a(gate131inter0), .b(s_322), .O(gate131inter1));
  and2  gate2803(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2804(.a(s_322), .O(gate131inter3));
  inv1  gate2805(.a(s_323), .O(gate131inter4));
  nand2 gate2806(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2807(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2808(.a(G414), .O(gate131inter7));
  inv1  gate2809(.a(G415), .O(gate131inter8));
  nand2 gate2810(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2811(.a(s_323), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2812(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2813(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2814(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate897(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate898(.a(gate134inter0), .b(s_50), .O(gate134inter1));
  and2  gate899(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate900(.a(s_50), .O(gate134inter3));
  inv1  gate901(.a(s_51), .O(gate134inter4));
  nand2 gate902(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate903(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate904(.a(G420), .O(gate134inter7));
  inv1  gate905(.a(G421), .O(gate134inter8));
  nand2 gate906(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate907(.a(s_51), .b(gate134inter3), .O(gate134inter10));
  nor2  gate908(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate909(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate910(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2003(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2004(.a(gate137inter0), .b(s_208), .O(gate137inter1));
  and2  gate2005(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2006(.a(s_208), .O(gate137inter3));
  inv1  gate2007(.a(s_209), .O(gate137inter4));
  nand2 gate2008(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2009(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2010(.a(G426), .O(gate137inter7));
  inv1  gate2011(.a(G429), .O(gate137inter8));
  nand2 gate2012(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2013(.a(s_209), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2014(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2015(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2016(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2311(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2312(.a(gate139inter0), .b(s_252), .O(gate139inter1));
  and2  gate2313(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2314(.a(s_252), .O(gate139inter3));
  inv1  gate2315(.a(s_253), .O(gate139inter4));
  nand2 gate2316(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2317(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2318(.a(G438), .O(gate139inter7));
  inv1  gate2319(.a(G441), .O(gate139inter8));
  nand2 gate2320(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2321(.a(s_253), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2322(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2323(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2324(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2395(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2396(.a(gate141inter0), .b(s_264), .O(gate141inter1));
  and2  gate2397(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2398(.a(s_264), .O(gate141inter3));
  inv1  gate2399(.a(s_265), .O(gate141inter4));
  nand2 gate2400(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2401(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2402(.a(G450), .O(gate141inter7));
  inv1  gate2403(.a(G453), .O(gate141inter8));
  nand2 gate2404(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2405(.a(s_265), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2406(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2407(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2408(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2871(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2872(.a(gate143inter0), .b(s_332), .O(gate143inter1));
  and2  gate2873(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2874(.a(s_332), .O(gate143inter3));
  inv1  gate2875(.a(s_333), .O(gate143inter4));
  nand2 gate2876(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2877(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2878(.a(G462), .O(gate143inter7));
  inv1  gate2879(.a(G465), .O(gate143inter8));
  nand2 gate2880(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2881(.a(s_333), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2882(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2883(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2884(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate2717(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2718(.a(gate144inter0), .b(s_310), .O(gate144inter1));
  and2  gate2719(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2720(.a(s_310), .O(gate144inter3));
  inv1  gate2721(.a(s_311), .O(gate144inter4));
  nand2 gate2722(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2723(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2724(.a(G468), .O(gate144inter7));
  inv1  gate2725(.a(G471), .O(gate144inter8));
  nand2 gate2726(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2727(.a(s_311), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2728(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2729(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2730(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2997(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2998(.a(gate145inter0), .b(s_350), .O(gate145inter1));
  and2  gate2999(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate3000(.a(s_350), .O(gate145inter3));
  inv1  gate3001(.a(s_351), .O(gate145inter4));
  nand2 gate3002(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate3003(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate3004(.a(G474), .O(gate145inter7));
  inv1  gate3005(.a(G477), .O(gate145inter8));
  nand2 gate3006(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate3007(.a(s_351), .b(gate145inter3), .O(gate145inter10));
  nor2  gate3008(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate3009(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate3010(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate827(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate828(.a(gate147inter0), .b(s_40), .O(gate147inter1));
  and2  gate829(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate830(.a(s_40), .O(gate147inter3));
  inv1  gate831(.a(s_41), .O(gate147inter4));
  nand2 gate832(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate833(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate834(.a(G486), .O(gate147inter7));
  inv1  gate835(.a(G489), .O(gate147inter8));
  nand2 gate836(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate837(.a(s_41), .b(gate147inter3), .O(gate147inter10));
  nor2  gate838(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate839(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate840(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2605(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2606(.a(gate150inter0), .b(s_294), .O(gate150inter1));
  and2  gate2607(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2608(.a(s_294), .O(gate150inter3));
  inv1  gate2609(.a(s_295), .O(gate150inter4));
  nand2 gate2610(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2611(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2612(.a(G504), .O(gate150inter7));
  inv1  gate2613(.a(G507), .O(gate150inter8));
  nand2 gate2614(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2615(.a(s_295), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2616(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2617(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2618(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1429(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1430(.a(gate151inter0), .b(s_126), .O(gate151inter1));
  and2  gate1431(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1432(.a(s_126), .O(gate151inter3));
  inv1  gate1433(.a(s_127), .O(gate151inter4));
  nand2 gate1434(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1435(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1436(.a(G510), .O(gate151inter7));
  inv1  gate1437(.a(G513), .O(gate151inter8));
  nand2 gate1438(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1439(.a(s_127), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1440(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1441(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1442(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate3277(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate3278(.a(gate156inter0), .b(s_390), .O(gate156inter1));
  and2  gate3279(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate3280(.a(s_390), .O(gate156inter3));
  inv1  gate3281(.a(s_391), .O(gate156inter4));
  nand2 gate3282(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate3283(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate3284(.a(G435), .O(gate156inter7));
  inv1  gate3285(.a(G525), .O(gate156inter8));
  nand2 gate3286(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate3287(.a(s_391), .b(gate156inter3), .O(gate156inter10));
  nor2  gate3288(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate3289(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate3290(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1205(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1206(.a(gate157inter0), .b(s_94), .O(gate157inter1));
  and2  gate1207(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1208(.a(s_94), .O(gate157inter3));
  inv1  gate1209(.a(s_95), .O(gate157inter4));
  nand2 gate1210(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1211(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1212(.a(G438), .O(gate157inter7));
  inv1  gate1213(.a(G528), .O(gate157inter8));
  nand2 gate1214(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1215(.a(s_95), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1216(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1217(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1218(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1737(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1738(.a(gate158inter0), .b(s_170), .O(gate158inter1));
  and2  gate1739(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1740(.a(s_170), .O(gate158inter3));
  inv1  gate1741(.a(s_171), .O(gate158inter4));
  nand2 gate1742(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1743(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1744(.a(G441), .O(gate158inter7));
  inv1  gate1745(.a(G528), .O(gate158inter8));
  nand2 gate1746(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1747(.a(s_171), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1748(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1749(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1750(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2283(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2284(.a(gate160inter0), .b(s_248), .O(gate160inter1));
  and2  gate2285(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2286(.a(s_248), .O(gate160inter3));
  inv1  gate2287(.a(s_249), .O(gate160inter4));
  nand2 gate2288(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2289(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2290(.a(G447), .O(gate160inter7));
  inv1  gate2291(.a(G531), .O(gate160inter8));
  nand2 gate2292(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2293(.a(s_249), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2294(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2295(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2296(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1471(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1472(.a(gate162inter0), .b(s_132), .O(gate162inter1));
  and2  gate1473(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1474(.a(s_132), .O(gate162inter3));
  inv1  gate1475(.a(s_133), .O(gate162inter4));
  nand2 gate1476(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1477(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1478(.a(G453), .O(gate162inter7));
  inv1  gate1479(.a(G534), .O(gate162inter8));
  nand2 gate1480(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1481(.a(s_133), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1482(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1483(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1484(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate687(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate688(.a(gate163inter0), .b(s_20), .O(gate163inter1));
  and2  gate689(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate690(.a(s_20), .O(gate163inter3));
  inv1  gate691(.a(s_21), .O(gate163inter4));
  nand2 gate692(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate693(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate694(.a(G456), .O(gate163inter7));
  inv1  gate695(.a(G537), .O(gate163inter8));
  nand2 gate696(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate697(.a(s_21), .b(gate163inter3), .O(gate163inter10));
  nor2  gate698(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate699(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate700(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1289(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1290(.a(gate164inter0), .b(s_106), .O(gate164inter1));
  and2  gate1291(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1292(.a(s_106), .O(gate164inter3));
  inv1  gate1293(.a(s_107), .O(gate164inter4));
  nand2 gate1294(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1295(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1296(.a(G459), .O(gate164inter7));
  inv1  gate1297(.a(G537), .O(gate164inter8));
  nand2 gate1298(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1299(.a(s_107), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1300(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1301(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1302(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2885(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2886(.a(gate166inter0), .b(s_334), .O(gate166inter1));
  and2  gate2887(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2888(.a(s_334), .O(gate166inter3));
  inv1  gate2889(.a(s_335), .O(gate166inter4));
  nand2 gate2890(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2891(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2892(.a(G465), .O(gate166inter7));
  inv1  gate2893(.a(G540), .O(gate166inter8));
  nand2 gate2894(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2895(.a(s_335), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2896(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2897(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2898(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1457(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1458(.a(gate169inter0), .b(s_130), .O(gate169inter1));
  and2  gate1459(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1460(.a(s_130), .O(gate169inter3));
  inv1  gate1461(.a(s_131), .O(gate169inter4));
  nand2 gate1462(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1463(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1464(.a(G474), .O(gate169inter7));
  inv1  gate1465(.a(G546), .O(gate169inter8));
  nand2 gate1466(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1467(.a(s_131), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1468(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1469(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1470(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1317(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1318(.a(gate170inter0), .b(s_110), .O(gate170inter1));
  and2  gate1319(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1320(.a(s_110), .O(gate170inter3));
  inv1  gate1321(.a(s_111), .O(gate170inter4));
  nand2 gate1322(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1323(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1324(.a(G477), .O(gate170inter7));
  inv1  gate1325(.a(G546), .O(gate170inter8));
  nand2 gate1326(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1327(.a(s_111), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1328(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1329(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1330(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1555(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1556(.a(gate178inter0), .b(s_144), .O(gate178inter1));
  and2  gate1557(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1558(.a(s_144), .O(gate178inter3));
  inv1  gate1559(.a(s_145), .O(gate178inter4));
  nand2 gate1560(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1561(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1562(.a(G501), .O(gate178inter7));
  inv1  gate1563(.a(G558), .O(gate178inter8));
  nand2 gate1564(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1565(.a(s_145), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1566(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1567(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1568(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate2703(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2704(.a(gate179inter0), .b(s_308), .O(gate179inter1));
  and2  gate2705(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2706(.a(s_308), .O(gate179inter3));
  inv1  gate2707(.a(s_309), .O(gate179inter4));
  nand2 gate2708(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2709(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2710(.a(G504), .O(gate179inter7));
  inv1  gate2711(.a(G561), .O(gate179inter8));
  nand2 gate2712(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2713(.a(s_309), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2714(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2715(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2716(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate967(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate968(.a(gate183inter0), .b(s_60), .O(gate183inter1));
  and2  gate969(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate970(.a(s_60), .O(gate183inter3));
  inv1  gate971(.a(s_61), .O(gate183inter4));
  nand2 gate972(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate973(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate974(.a(G516), .O(gate183inter7));
  inv1  gate975(.a(G567), .O(gate183inter8));
  nand2 gate976(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate977(.a(s_61), .b(gate183inter3), .O(gate183inter10));
  nor2  gate978(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate979(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate980(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2171(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2172(.a(gate185inter0), .b(s_232), .O(gate185inter1));
  and2  gate2173(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2174(.a(s_232), .O(gate185inter3));
  inv1  gate2175(.a(s_233), .O(gate185inter4));
  nand2 gate2176(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2177(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2178(.a(G570), .O(gate185inter7));
  inv1  gate2179(.a(G571), .O(gate185inter8));
  nand2 gate2180(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2181(.a(s_233), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2182(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2183(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2184(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1849(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1850(.a(gate188inter0), .b(s_186), .O(gate188inter1));
  and2  gate1851(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1852(.a(s_186), .O(gate188inter3));
  inv1  gate1853(.a(s_187), .O(gate188inter4));
  nand2 gate1854(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1855(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1856(.a(G576), .O(gate188inter7));
  inv1  gate1857(.a(G577), .O(gate188inter8));
  nand2 gate1858(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1859(.a(s_187), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1860(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1861(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1862(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2115(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2116(.a(gate189inter0), .b(s_224), .O(gate189inter1));
  and2  gate2117(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2118(.a(s_224), .O(gate189inter3));
  inv1  gate2119(.a(s_225), .O(gate189inter4));
  nand2 gate2120(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2121(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2122(.a(G578), .O(gate189inter7));
  inv1  gate2123(.a(G579), .O(gate189inter8));
  nand2 gate2124(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2125(.a(s_225), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2126(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2127(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2128(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate785(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate786(.a(gate191inter0), .b(s_34), .O(gate191inter1));
  and2  gate787(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate788(.a(s_34), .O(gate191inter3));
  inv1  gate789(.a(s_35), .O(gate191inter4));
  nand2 gate790(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate791(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate792(.a(G582), .O(gate191inter7));
  inv1  gate793(.a(G583), .O(gate191inter8));
  nand2 gate794(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate795(.a(s_35), .b(gate191inter3), .O(gate191inter10));
  nor2  gate796(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate797(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate798(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate589(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate590(.a(gate192inter0), .b(s_6), .O(gate192inter1));
  and2  gate591(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate592(.a(s_6), .O(gate192inter3));
  inv1  gate593(.a(s_7), .O(gate192inter4));
  nand2 gate594(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate595(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate596(.a(G584), .O(gate192inter7));
  inv1  gate597(.a(G585), .O(gate192inter8));
  nand2 gate598(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate599(.a(s_7), .b(gate192inter3), .O(gate192inter10));
  nor2  gate600(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate601(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate602(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2437(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2438(.a(gate194inter0), .b(s_270), .O(gate194inter1));
  and2  gate2439(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2440(.a(s_270), .O(gate194inter3));
  inv1  gate2441(.a(s_271), .O(gate194inter4));
  nand2 gate2442(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2443(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2444(.a(G588), .O(gate194inter7));
  inv1  gate2445(.a(G589), .O(gate194inter8));
  nand2 gate2446(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2447(.a(s_271), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2448(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2449(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2450(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2745(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2746(.a(gate197inter0), .b(s_314), .O(gate197inter1));
  and2  gate2747(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2748(.a(s_314), .O(gate197inter3));
  inv1  gate2749(.a(s_315), .O(gate197inter4));
  nand2 gate2750(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2751(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2752(.a(G594), .O(gate197inter7));
  inv1  gate2753(.a(G595), .O(gate197inter8));
  nand2 gate2754(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2755(.a(s_315), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2756(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2757(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2758(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate3291(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate3292(.a(gate201inter0), .b(s_392), .O(gate201inter1));
  and2  gate3293(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate3294(.a(s_392), .O(gate201inter3));
  inv1  gate3295(.a(s_393), .O(gate201inter4));
  nand2 gate3296(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate3297(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate3298(.a(G602), .O(gate201inter7));
  inv1  gate3299(.a(G607), .O(gate201inter8));
  nand2 gate3300(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate3301(.a(s_393), .b(gate201inter3), .O(gate201inter10));
  nor2  gate3302(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate3303(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate3304(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2619(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2620(.a(gate203inter0), .b(s_296), .O(gate203inter1));
  and2  gate2621(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2622(.a(s_296), .O(gate203inter3));
  inv1  gate2623(.a(s_297), .O(gate203inter4));
  nand2 gate2624(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2625(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2626(.a(G602), .O(gate203inter7));
  inv1  gate2627(.a(G612), .O(gate203inter8));
  nand2 gate2628(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2629(.a(s_297), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2630(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2631(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2632(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate3249(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate3250(.a(gate204inter0), .b(s_386), .O(gate204inter1));
  and2  gate3251(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate3252(.a(s_386), .O(gate204inter3));
  inv1  gate3253(.a(s_387), .O(gate204inter4));
  nand2 gate3254(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate3255(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate3256(.a(G607), .O(gate204inter7));
  inv1  gate3257(.a(G617), .O(gate204inter8));
  nand2 gate3258(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate3259(.a(s_387), .b(gate204inter3), .O(gate204inter10));
  nor2  gate3260(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate3261(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate3262(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1191(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1192(.a(gate207inter0), .b(s_92), .O(gate207inter1));
  and2  gate1193(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1194(.a(s_92), .O(gate207inter3));
  inv1  gate1195(.a(s_93), .O(gate207inter4));
  nand2 gate1196(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1197(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1198(.a(G622), .O(gate207inter7));
  inv1  gate1199(.a(G632), .O(gate207inter8));
  nand2 gate1200(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1201(.a(s_93), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1202(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1203(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1204(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate3011(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate3012(.a(gate210inter0), .b(s_352), .O(gate210inter1));
  and2  gate3013(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate3014(.a(s_352), .O(gate210inter3));
  inv1  gate3015(.a(s_353), .O(gate210inter4));
  nand2 gate3016(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate3017(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate3018(.a(G607), .O(gate210inter7));
  inv1  gate3019(.a(G666), .O(gate210inter8));
  nand2 gate3020(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate3021(.a(s_353), .b(gate210inter3), .O(gate210inter10));
  nor2  gate3022(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate3023(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate3024(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate2353(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2354(.a(gate211inter0), .b(s_258), .O(gate211inter1));
  and2  gate2355(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2356(.a(s_258), .O(gate211inter3));
  inv1  gate2357(.a(s_259), .O(gate211inter4));
  nand2 gate2358(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2359(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2360(.a(G612), .O(gate211inter7));
  inv1  gate2361(.a(G669), .O(gate211inter8));
  nand2 gate2362(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2363(.a(s_259), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2364(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2365(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2366(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2913(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2914(.a(gate212inter0), .b(s_338), .O(gate212inter1));
  and2  gate2915(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2916(.a(s_338), .O(gate212inter3));
  inv1  gate2917(.a(s_339), .O(gate212inter4));
  nand2 gate2918(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2919(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2920(.a(G617), .O(gate212inter7));
  inv1  gate2921(.a(G669), .O(gate212inter8));
  nand2 gate2922(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2923(.a(s_339), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2924(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2925(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2926(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2199(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2200(.a(gate214inter0), .b(s_236), .O(gate214inter1));
  and2  gate2201(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2202(.a(s_236), .O(gate214inter3));
  inv1  gate2203(.a(s_237), .O(gate214inter4));
  nand2 gate2204(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2205(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2206(.a(G612), .O(gate214inter7));
  inv1  gate2207(.a(G672), .O(gate214inter8));
  nand2 gate2208(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2209(.a(s_237), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2210(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2211(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2212(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1863(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1864(.a(gate215inter0), .b(s_188), .O(gate215inter1));
  and2  gate1865(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1866(.a(s_188), .O(gate215inter3));
  inv1  gate1867(.a(s_189), .O(gate215inter4));
  nand2 gate1868(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1869(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1870(.a(G607), .O(gate215inter7));
  inv1  gate1871(.a(G675), .O(gate215inter8));
  nand2 gate1872(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1873(.a(s_189), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1874(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1875(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1876(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2157(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2158(.a(gate219inter0), .b(s_230), .O(gate219inter1));
  and2  gate2159(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2160(.a(s_230), .O(gate219inter3));
  inv1  gate2161(.a(s_231), .O(gate219inter4));
  nand2 gate2162(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2163(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2164(.a(G632), .O(gate219inter7));
  inv1  gate2165(.a(G681), .O(gate219inter8));
  nand2 gate2166(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2167(.a(s_231), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2168(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2169(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2170(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1569(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1570(.a(gate220inter0), .b(s_146), .O(gate220inter1));
  and2  gate1571(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1572(.a(s_146), .O(gate220inter3));
  inv1  gate1573(.a(s_147), .O(gate220inter4));
  nand2 gate1574(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1575(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1576(.a(G637), .O(gate220inter7));
  inv1  gate1577(.a(G681), .O(gate220inter8));
  nand2 gate1578(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1579(.a(s_147), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1580(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1581(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1582(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1051(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1052(.a(gate221inter0), .b(s_72), .O(gate221inter1));
  and2  gate1053(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1054(.a(s_72), .O(gate221inter3));
  inv1  gate1055(.a(s_73), .O(gate221inter4));
  nand2 gate1056(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1057(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1058(.a(G622), .O(gate221inter7));
  inv1  gate1059(.a(G684), .O(gate221inter8));
  nand2 gate1060(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1061(.a(s_73), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1062(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1063(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1064(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1947(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1948(.a(gate223inter0), .b(s_200), .O(gate223inter1));
  and2  gate1949(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1950(.a(s_200), .O(gate223inter3));
  inv1  gate1951(.a(s_201), .O(gate223inter4));
  nand2 gate1952(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1953(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1954(.a(G627), .O(gate223inter7));
  inv1  gate1955(.a(G687), .O(gate223inter8));
  nand2 gate1956(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1957(.a(s_201), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1958(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1959(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1960(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate911(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate912(.a(gate224inter0), .b(s_52), .O(gate224inter1));
  and2  gate913(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate914(.a(s_52), .O(gate224inter3));
  inv1  gate915(.a(s_53), .O(gate224inter4));
  nand2 gate916(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate917(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate918(.a(G637), .O(gate224inter7));
  inv1  gate919(.a(G687), .O(gate224inter8));
  nand2 gate920(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate921(.a(s_53), .b(gate224inter3), .O(gate224inter10));
  nor2  gate922(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate923(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate924(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2675(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2676(.a(gate227inter0), .b(s_304), .O(gate227inter1));
  and2  gate2677(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2678(.a(s_304), .O(gate227inter3));
  inv1  gate2679(.a(s_305), .O(gate227inter4));
  nand2 gate2680(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2681(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2682(.a(G694), .O(gate227inter7));
  inv1  gate2683(.a(G695), .O(gate227inter8));
  nand2 gate2684(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2685(.a(s_305), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2686(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2687(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2688(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate771(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate772(.a(gate228inter0), .b(s_32), .O(gate228inter1));
  and2  gate773(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate774(.a(s_32), .O(gate228inter3));
  inv1  gate775(.a(s_33), .O(gate228inter4));
  nand2 gate776(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate777(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate778(.a(G696), .O(gate228inter7));
  inv1  gate779(.a(G697), .O(gate228inter8));
  nand2 gate780(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate781(.a(s_33), .b(gate228inter3), .O(gate228inter10));
  nor2  gate782(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate783(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate784(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2325(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2326(.a(gate232inter0), .b(s_254), .O(gate232inter1));
  and2  gate2327(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2328(.a(s_254), .O(gate232inter3));
  inv1  gate2329(.a(s_255), .O(gate232inter4));
  nand2 gate2330(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2331(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2332(.a(G704), .O(gate232inter7));
  inv1  gate2333(.a(G705), .O(gate232inter8));
  nand2 gate2334(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2335(.a(s_255), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2336(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2337(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2338(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2465(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2466(.a(gate234inter0), .b(s_274), .O(gate234inter1));
  and2  gate2467(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2468(.a(s_274), .O(gate234inter3));
  inv1  gate2469(.a(s_275), .O(gate234inter4));
  nand2 gate2470(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2471(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2472(.a(G245), .O(gate234inter7));
  inv1  gate2473(.a(G721), .O(gate234inter8));
  nand2 gate2474(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2475(.a(s_275), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2476(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2477(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2478(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate841(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate842(.a(gate235inter0), .b(s_42), .O(gate235inter1));
  and2  gate843(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate844(.a(s_42), .O(gate235inter3));
  inv1  gate845(.a(s_43), .O(gate235inter4));
  nand2 gate846(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate847(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate848(.a(G248), .O(gate235inter7));
  inv1  gate849(.a(G724), .O(gate235inter8));
  nand2 gate850(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate851(.a(s_43), .b(gate235inter3), .O(gate235inter10));
  nor2  gate852(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate853(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate854(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1373(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1374(.a(gate238inter0), .b(s_118), .O(gate238inter1));
  and2  gate1375(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1376(.a(s_118), .O(gate238inter3));
  inv1  gate1377(.a(s_119), .O(gate238inter4));
  nand2 gate1378(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1379(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1380(.a(G257), .O(gate238inter7));
  inv1  gate1381(.a(G709), .O(gate238inter8));
  nand2 gate1382(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1383(.a(s_119), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1384(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1385(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1386(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2507(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2508(.a(gate239inter0), .b(s_280), .O(gate239inter1));
  and2  gate2509(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2510(.a(s_280), .O(gate239inter3));
  inv1  gate2511(.a(s_281), .O(gate239inter4));
  nand2 gate2512(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2513(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2514(.a(G260), .O(gate239inter7));
  inv1  gate2515(.a(G712), .O(gate239inter8));
  nand2 gate2516(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2517(.a(s_281), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2518(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2519(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2520(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1933(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1934(.a(gate241inter0), .b(s_198), .O(gate241inter1));
  and2  gate1935(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1936(.a(s_198), .O(gate241inter3));
  inv1  gate1937(.a(s_199), .O(gate241inter4));
  nand2 gate1938(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1939(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1940(.a(G242), .O(gate241inter7));
  inv1  gate1941(.a(G730), .O(gate241inter8));
  nand2 gate1942(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1943(.a(s_199), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1944(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1945(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1946(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2941(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2942(.a(gate243inter0), .b(s_342), .O(gate243inter1));
  and2  gate2943(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2944(.a(s_342), .O(gate243inter3));
  inv1  gate2945(.a(s_343), .O(gate243inter4));
  nand2 gate2946(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2947(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2948(.a(G245), .O(gate243inter7));
  inv1  gate2949(.a(G733), .O(gate243inter8));
  nand2 gate2950(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2951(.a(s_343), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2952(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2953(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2954(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate995(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate996(.a(gate245inter0), .b(s_64), .O(gate245inter1));
  and2  gate997(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate998(.a(s_64), .O(gate245inter3));
  inv1  gate999(.a(s_65), .O(gate245inter4));
  nand2 gate1000(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1001(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1002(.a(G248), .O(gate245inter7));
  inv1  gate1003(.a(G736), .O(gate245inter8));
  nand2 gate1004(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1005(.a(s_65), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1006(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1007(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1008(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2535(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2536(.a(gate247inter0), .b(s_284), .O(gate247inter1));
  and2  gate2537(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2538(.a(s_284), .O(gate247inter3));
  inv1  gate2539(.a(s_285), .O(gate247inter4));
  nand2 gate2540(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2541(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2542(.a(G251), .O(gate247inter7));
  inv1  gate2543(.a(G739), .O(gate247inter8));
  nand2 gate2544(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2545(.a(s_285), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2546(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2547(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2548(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1681(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1682(.a(gate248inter0), .b(s_162), .O(gate248inter1));
  and2  gate1683(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1684(.a(s_162), .O(gate248inter3));
  inv1  gate1685(.a(s_163), .O(gate248inter4));
  nand2 gate1686(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1687(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1688(.a(G727), .O(gate248inter7));
  inv1  gate1689(.a(G739), .O(gate248inter8));
  nand2 gate1690(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1691(.a(s_163), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1692(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1693(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1694(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1527(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1528(.a(gate250inter0), .b(s_140), .O(gate250inter1));
  and2  gate1529(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1530(.a(s_140), .O(gate250inter3));
  inv1  gate1531(.a(s_141), .O(gate250inter4));
  nand2 gate1532(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1533(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1534(.a(G706), .O(gate250inter7));
  inv1  gate1535(.a(G742), .O(gate250inter8));
  nand2 gate1536(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1537(.a(s_141), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1538(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1539(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1540(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate925(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate926(.a(gate251inter0), .b(s_54), .O(gate251inter1));
  and2  gate927(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate928(.a(s_54), .O(gate251inter3));
  inv1  gate929(.a(s_55), .O(gate251inter4));
  nand2 gate930(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate931(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate932(.a(G257), .O(gate251inter7));
  inv1  gate933(.a(G745), .O(gate251inter8));
  nand2 gate934(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate935(.a(s_55), .b(gate251inter3), .O(gate251inter10));
  nor2  gate936(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate937(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate938(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1499(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1500(.a(gate252inter0), .b(s_136), .O(gate252inter1));
  and2  gate1501(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1502(.a(s_136), .O(gate252inter3));
  inv1  gate1503(.a(s_137), .O(gate252inter4));
  nand2 gate1504(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1505(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1506(.a(G709), .O(gate252inter7));
  inv1  gate1507(.a(G745), .O(gate252inter8));
  nand2 gate1508(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1509(.a(s_137), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1510(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1511(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1512(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1667(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1668(.a(gate254inter0), .b(s_160), .O(gate254inter1));
  and2  gate1669(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1670(.a(s_160), .O(gate254inter3));
  inv1  gate1671(.a(s_161), .O(gate254inter4));
  nand2 gate1672(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1673(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1674(.a(G712), .O(gate254inter7));
  inv1  gate1675(.a(G748), .O(gate254inter8));
  nand2 gate1676(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1677(.a(s_161), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1678(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1679(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1680(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate2815(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2816(.a(gate255inter0), .b(s_324), .O(gate255inter1));
  and2  gate2817(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2818(.a(s_324), .O(gate255inter3));
  inv1  gate2819(.a(s_325), .O(gate255inter4));
  nand2 gate2820(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2821(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2822(.a(G263), .O(gate255inter7));
  inv1  gate2823(.a(G751), .O(gate255inter8));
  nand2 gate2824(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2825(.a(s_325), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2826(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2827(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2828(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate3039(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate3040(.a(gate256inter0), .b(s_356), .O(gate256inter1));
  and2  gate3041(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate3042(.a(s_356), .O(gate256inter3));
  inv1  gate3043(.a(s_357), .O(gate256inter4));
  nand2 gate3044(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate3045(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate3046(.a(G715), .O(gate256inter7));
  inv1  gate3047(.a(G751), .O(gate256inter8));
  nand2 gate3048(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate3049(.a(s_357), .b(gate256inter3), .O(gate256inter10));
  nor2  gate3050(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate3051(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate3052(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate3263(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate3264(.a(gate257inter0), .b(s_388), .O(gate257inter1));
  and2  gate3265(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate3266(.a(s_388), .O(gate257inter3));
  inv1  gate3267(.a(s_389), .O(gate257inter4));
  nand2 gate3268(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate3269(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate3270(.a(G754), .O(gate257inter7));
  inv1  gate3271(.a(G755), .O(gate257inter8));
  nand2 gate3272(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate3273(.a(s_389), .b(gate257inter3), .O(gate257inter10));
  nor2  gate3274(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate3275(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate3276(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1177(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1178(.a(gate258inter0), .b(s_90), .O(gate258inter1));
  and2  gate1179(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1180(.a(s_90), .O(gate258inter3));
  inv1  gate1181(.a(s_91), .O(gate258inter4));
  nand2 gate1182(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1183(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1184(.a(G756), .O(gate258inter7));
  inv1  gate1185(.a(G757), .O(gate258inter8));
  nand2 gate1186(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1187(.a(s_91), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1188(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1189(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1190(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate2521(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2522(.a(gate259inter0), .b(s_282), .O(gate259inter1));
  and2  gate2523(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2524(.a(s_282), .O(gate259inter3));
  inv1  gate2525(.a(s_283), .O(gate259inter4));
  nand2 gate2526(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2527(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2528(.a(G758), .O(gate259inter7));
  inv1  gate2529(.a(G759), .O(gate259inter8));
  nand2 gate2530(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2531(.a(s_283), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2532(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2533(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2534(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1961(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1962(.a(gate261inter0), .b(s_202), .O(gate261inter1));
  and2  gate1963(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1964(.a(s_202), .O(gate261inter3));
  inv1  gate1965(.a(s_203), .O(gate261inter4));
  nand2 gate1966(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1967(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1968(.a(G762), .O(gate261inter7));
  inv1  gate1969(.a(G763), .O(gate261inter8));
  nand2 gate1970(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1971(.a(s_203), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1972(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1973(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1974(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate3137(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate3138(.a(gate262inter0), .b(s_370), .O(gate262inter1));
  and2  gate3139(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate3140(.a(s_370), .O(gate262inter3));
  inv1  gate3141(.a(s_371), .O(gate262inter4));
  nand2 gate3142(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate3143(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate3144(.a(G764), .O(gate262inter7));
  inv1  gate3145(.a(G765), .O(gate262inter8));
  nand2 gate3146(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate3147(.a(s_371), .b(gate262inter3), .O(gate262inter10));
  nor2  gate3148(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate3149(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate3150(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1247(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1248(.a(gate264inter0), .b(s_100), .O(gate264inter1));
  and2  gate1249(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1250(.a(s_100), .O(gate264inter3));
  inv1  gate1251(.a(s_101), .O(gate264inter4));
  nand2 gate1252(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1253(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1254(.a(G768), .O(gate264inter7));
  inv1  gate1255(.a(G769), .O(gate264inter8));
  nand2 gate1256(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1257(.a(s_101), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1258(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1259(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1260(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate2563(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2564(.a(gate265inter0), .b(s_288), .O(gate265inter1));
  and2  gate2565(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2566(.a(s_288), .O(gate265inter3));
  inv1  gate2567(.a(s_289), .O(gate265inter4));
  nand2 gate2568(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2569(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2570(.a(G642), .O(gate265inter7));
  inv1  gate2571(.a(G770), .O(gate265inter8));
  nand2 gate2572(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2573(.a(s_289), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2574(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2575(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2576(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1485(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1486(.a(gate266inter0), .b(s_134), .O(gate266inter1));
  and2  gate1487(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1488(.a(s_134), .O(gate266inter3));
  inv1  gate1489(.a(s_135), .O(gate266inter4));
  nand2 gate1490(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1491(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1492(.a(G645), .O(gate266inter7));
  inv1  gate1493(.a(G773), .O(gate266inter8));
  nand2 gate1494(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1495(.a(s_135), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1496(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1497(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1498(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate3333(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate3334(.a(gate267inter0), .b(s_398), .O(gate267inter1));
  and2  gate3335(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate3336(.a(s_398), .O(gate267inter3));
  inv1  gate3337(.a(s_399), .O(gate267inter4));
  nand2 gate3338(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate3339(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate3340(.a(G648), .O(gate267inter7));
  inv1  gate3341(.a(G776), .O(gate267inter8));
  nand2 gate3342(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate3343(.a(s_399), .b(gate267inter3), .O(gate267inter10));
  nor2  gate3344(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate3345(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate3346(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate3179(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate3180(.a(gate270inter0), .b(s_376), .O(gate270inter1));
  and2  gate3181(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate3182(.a(s_376), .O(gate270inter3));
  inv1  gate3183(.a(s_377), .O(gate270inter4));
  nand2 gate3184(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate3185(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate3186(.a(G657), .O(gate270inter7));
  inv1  gate3187(.a(G785), .O(gate270inter8));
  nand2 gate3188(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate3189(.a(s_377), .b(gate270inter3), .O(gate270inter10));
  nor2  gate3190(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate3191(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate3192(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2843(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2844(.a(gate273inter0), .b(s_328), .O(gate273inter1));
  and2  gate2845(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2846(.a(s_328), .O(gate273inter3));
  inv1  gate2847(.a(s_329), .O(gate273inter4));
  nand2 gate2848(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2849(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2850(.a(G642), .O(gate273inter7));
  inv1  gate2851(.a(G794), .O(gate273inter8));
  nand2 gate2852(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2853(.a(s_329), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2854(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2855(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2856(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate3025(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate3026(.a(gate276inter0), .b(s_354), .O(gate276inter1));
  and2  gate3027(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate3028(.a(s_354), .O(gate276inter3));
  inv1  gate3029(.a(s_355), .O(gate276inter4));
  nand2 gate3030(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate3031(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate3032(.a(G773), .O(gate276inter7));
  inv1  gate3033(.a(G797), .O(gate276inter8));
  nand2 gate3034(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate3035(.a(s_355), .b(gate276inter3), .O(gate276inter10));
  nor2  gate3036(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate3037(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate3038(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate3347(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate3348(.a(gate278inter0), .b(s_400), .O(gate278inter1));
  and2  gate3349(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate3350(.a(s_400), .O(gate278inter3));
  inv1  gate3351(.a(s_401), .O(gate278inter4));
  nand2 gate3352(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate3353(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate3354(.a(G776), .O(gate278inter7));
  inv1  gate3355(.a(G800), .O(gate278inter8));
  nand2 gate3356(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate3357(.a(s_401), .b(gate278inter3), .O(gate278inter10));
  nor2  gate3358(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate3359(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate3360(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1639(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1640(.a(gate279inter0), .b(s_156), .O(gate279inter1));
  and2  gate1641(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1642(.a(s_156), .O(gate279inter3));
  inv1  gate1643(.a(s_157), .O(gate279inter4));
  nand2 gate1644(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1645(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1646(.a(G651), .O(gate279inter7));
  inv1  gate1647(.a(G803), .O(gate279inter8));
  nand2 gate1648(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1649(.a(s_157), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1650(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1651(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1652(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1065(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1066(.a(gate280inter0), .b(s_74), .O(gate280inter1));
  and2  gate1067(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1068(.a(s_74), .O(gate280inter3));
  inv1  gate1069(.a(s_75), .O(gate280inter4));
  nand2 gate1070(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1071(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1072(.a(G779), .O(gate280inter7));
  inv1  gate1073(.a(G803), .O(gate280inter8));
  nand2 gate1074(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1075(.a(s_75), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1076(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1077(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1078(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2857(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2858(.a(gate282inter0), .b(s_330), .O(gate282inter1));
  and2  gate2859(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2860(.a(s_330), .O(gate282inter3));
  inv1  gate2861(.a(s_331), .O(gate282inter4));
  nand2 gate2862(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2863(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2864(.a(G782), .O(gate282inter7));
  inv1  gate2865(.a(G806), .O(gate282inter8));
  nand2 gate2866(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2867(.a(s_331), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2868(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2869(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2870(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate939(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate940(.a(gate283inter0), .b(s_56), .O(gate283inter1));
  and2  gate941(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate942(.a(s_56), .O(gate283inter3));
  inv1  gate943(.a(s_57), .O(gate283inter4));
  nand2 gate944(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate945(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate946(.a(G657), .O(gate283inter7));
  inv1  gate947(.a(G809), .O(gate283inter8));
  nand2 gate948(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate949(.a(s_57), .b(gate283inter3), .O(gate283inter10));
  nor2  gate950(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate951(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate952(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate701(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate702(.a(gate285inter0), .b(s_22), .O(gate285inter1));
  and2  gate703(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate704(.a(s_22), .O(gate285inter3));
  inv1  gate705(.a(s_23), .O(gate285inter4));
  nand2 gate706(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate707(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate708(.a(G660), .O(gate285inter7));
  inv1  gate709(.a(G812), .O(gate285inter8));
  nand2 gate710(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate711(.a(s_23), .b(gate285inter3), .O(gate285inter10));
  nor2  gate712(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate713(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate714(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate3081(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate3082(.a(gate293inter0), .b(s_362), .O(gate293inter1));
  and2  gate3083(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate3084(.a(s_362), .O(gate293inter3));
  inv1  gate3085(.a(s_363), .O(gate293inter4));
  nand2 gate3086(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate3087(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate3088(.a(G828), .O(gate293inter7));
  inv1  gate3089(.a(G829), .O(gate293inter8));
  nand2 gate3090(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate3091(.a(s_363), .b(gate293inter3), .O(gate293inter10));
  nor2  gate3092(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate3093(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate3094(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate547(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate548(.a(gate294inter0), .b(s_0), .O(gate294inter1));
  and2  gate549(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate550(.a(s_0), .O(gate294inter3));
  inv1  gate551(.a(s_1), .O(gate294inter4));
  nand2 gate552(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate553(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate554(.a(G832), .O(gate294inter7));
  inv1  gate555(.a(G833), .O(gate294inter8));
  nand2 gate556(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate557(.a(s_1), .b(gate294inter3), .O(gate294inter10));
  nor2  gate558(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate559(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate560(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate3305(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate3306(.a(gate295inter0), .b(s_394), .O(gate295inter1));
  and2  gate3307(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate3308(.a(s_394), .O(gate295inter3));
  inv1  gate3309(.a(s_395), .O(gate295inter4));
  nand2 gate3310(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate3311(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate3312(.a(G830), .O(gate295inter7));
  inv1  gate3313(.a(G831), .O(gate295inter8));
  nand2 gate3314(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate3315(.a(s_395), .b(gate295inter3), .O(gate295inter10));
  nor2  gate3316(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate3317(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate3318(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate3165(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate3166(.a(gate388inter0), .b(s_374), .O(gate388inter1));
  and2  gate3167(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate3168(.a(s_374), .O(gate388inter3));
  inv1  gate3169(.a(s_375), .O(gate388inter4));
  nand2 gate3170(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate3171(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate3172(.a(G2), .O(gate388inter7));
  inv1  gate3173(.a(G1039), .O(gate388inter8));
  nand2 gate3174(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate3175(.a(s_375), .b(gate388inter3), .O(gate388inter10));
  nor2  gate3176(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate3177(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate3178(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate953(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate954(.a(gate390inter0), .b(s_58), .O(gate390inter1));
  and2  gate955(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate956(.a(s_58), .O(gate390inter3));
  inv1  gate957(.a(s_59), .O(gate390inter4));
  nand2 gate958(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate959(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate960(.a(G4), .O(gate390inter7));
  inv1  gate961(.a(G1045), .O(gate390inter8));
  nand2 gate962(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate963(.a(s_59), .b(gate390inter3), .O(gate390inter10));
  nor2  gate964(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate965(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate966(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1401(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1402(.a(gate396inter0), .b(s_122), .O(gate396inter1));
  and2  gate1403(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1404(.a(s_122), .O(gate396inter3));
  inv1  gate1405(.a(s_123), .O(gate396inter4));
  nand2 gate1406(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1407(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1408(.a(G10), .O(gate396inter7));
  inv1  gate1409(.a(G1063), .O(gate396inter8));
  nand2 gate1410(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1411(.a(s_123), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1412(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1413(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1414(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1149(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1150(.a(gate399inter0), .b(s_86), .O(gate399inter1));
  and2  gate1151(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1152(.a(s_86), .O(gate399inter3));
  inv1  gate1153(.a(s_87), .O(gate399inter4));
  nand2 gate1154(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1155(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1156(.a(G13), .O(gate399inter7));
  inv1  gate1157(.a(G1072), .O(gate399inter8));
  nand2 gate1158(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1159(.a(s_87), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1160(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1161(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1162(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1611(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1612(.a(gate403inter0), .b(s_152), .O(gate403inter1));
  and2  gate1613(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1614(.a(s_152), .O(gate403inter3));
  inv1  gate1615(.a(s_153), .O(gate403inter4));
  nand2 gate1616(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1617(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1618(.a(G17), .O(gate403inter7));
  inv1  gate1619(.a(G1084), .O(gate403inter8));
  nand2 gate1620(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1621(.a(s_153), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1622(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1623(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1624(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2297(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2298(.a(gate406inter0), .b(s_250), .O(gate406inter1));
  and2  gate2299(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2300(.a(s_250), .O(gate406inter3));
  inv1  gate2301(.a(s_251), .O(gate406inter4));
  nand2 gate2302(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2303(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2304(.a(G20), .O(gate406inter7));
  inv1  gate2305(.a(G1093), .O(gate406inter8));
  nand2 gate2306(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2307(.a(s_251), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2308(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2309(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2310(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1261(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1262(.a(gate408inter0), .b(s_102), .O(gate408inter1));
  and2  gate1263(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1264(.a(s_102), .O(gate408inter3));
  inv1  gate1265(.a(s_103), .O(gate408inter4));
  nand2 gate1266(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1267(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1268(.a(G22), .O(gate408inter7));
  inv1  gate1269(.a(G1099), .O(gate408inter8));
  nand2 gate1270(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1271(.a(s_103), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1272(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1273(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1274(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate855(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate856(.a(gate410inter0), .b(s_44), .O(gate410inter1));
  and2  gate857(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate858(.a(s_44), .O(gate410inter3));
  inv1  gate859(.a(s_45), .O(gate410inter4));
  nand2 gate860(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate861(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate862(.a(G24), .O(gate410inter7));
  inv1  gate863(.a(G1105), .O(gate410inter8));
  nand2 gate864(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate865(.a(s_45), .b(gate410inter3), .O(gate410inter10));
  nor2  gate866(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate867(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate868(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1597(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1598(.a(gate411inter0), .b(s_150), .O(gate411inter1));
  and2  gate1599(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1600(.a(s_150), .O(gate411inter3));
  inv1  gate1601(.a(s_151), .O(gate411inter4));
  nand2 gate1602(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1603(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1604(.a(G25), .O(gate411inter7));
  inv1  gate1605(.a(G1108), .O(gate411inter8));
  nand2 gate1606(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1607(.a(s_151), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1608(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1609(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1610(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1723(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1724(.a(gate412inter0), .b(s_168), .O(gate412inter1));
  and2  gate1725(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1726(.a(s_168), .O(gate412inter3));
  inv1  gate1727(.a(s_169), .O(gate412inter4));
  nand2 gate1728(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1729(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1730(.a(G26), .O(gate412inter7));
  inv1  gate1731(.a(G1111), .O(gate412inter8));
  nand2 gate1732(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1733(.a(s_169), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1734(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1735(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1736(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate2955(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2956(.a(gate413inter0), .b(s_344), .O(gate413inter1));
  and2  gate2957(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2958(.a(s_344), .O(gate413inter3));
  inv1  gate2959(.a(s_345), .O(gate413inter4));
  nand2 gate2960(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2961(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2962(.a(G27), .O(gate413inter7));
  inv1  gate2963(.a(G1114), .O(gate413inter8));
  nand2 gate2964(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2965(.a(s_345), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2966(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2967(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2968(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate603(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate604(.a(gate417inter0), .b(s_8), .O(gate417inter1));
  and2  gate605(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate606(.a(s_8), .O(gate417inter3));
  inv1  gate607(.a(s_9), .O(gate417inter4));
  nand2 gate608(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate609(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate610(.a(G31), .O(gate417inter7));
  inv1  gate611(.a(G1126), .O(gate417inter8));
  nand2 gate612(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate613(.a(s_9), .b(gate417inter3), .O(gate417inter10));
  nor2  gate614(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate615(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate616(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2143(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2144(.a(gate419inter0), .b(s_228), .O(gate419inter1));
  and2  gate2145(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2146(.a(s_228), .O(gate419inter3));
  inv1  gate2147(.a(s_229), .O(gate419inter4));
  nand2 gate2148(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2149(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2150(.a(G1), .O(gate419inter7));
  inv1  gate2151(.a(G1132), .O(gate419inter8));
  nand2 gate2152(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2153(.a(s_229), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2154(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2155(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2156(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2367(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2368(.a(gate422inter0), .b(s_260), .O(gate422inter1));
  and2  gate2369(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2370(.a(s_260), .O(gate422inter3));
  inv1  gate2371(.a(s_261), .O(gate422inter4));
  nand2 gate2372(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2373(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2374(.a(G1039), .O(gate422inter7));
  inv1  gate2375(.a(G1135), .O(gate422inter8));
  nand2 gate2376(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2377(.a(s_261), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2378(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2379(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2380(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate813(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate814(.a(gate423inter0), .b(s_38), .O(gate423inter1));
  and2  gate815(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate816(.a(s_38), .O(gate423inter3));
  inv1  gate817(.a(s_39), .O(gate423inter4));
  nand2 gate818(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate819(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate820(.a(G3), .O(gate423inter7));
  inv1  gate821(.a(G1138), .O(gate423inter8));
  nand2 gate822(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate823(.a(s_39), .b(gate423inter3), .O(gate423inter10));
  nor2  gate824(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate825(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate826(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate3235(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate3236(.a(gate425inter0), .b(s_384), .O(gate425inter1));
  and2  gate3237(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate3238(.a(s_384), .O(gate425inter3));
  inv1  gate3239(.a(s_385), .O(gate425inter4));
  nand2 gate3240(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate3241(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate3242(.a(G4), .O(gate425inter7));
  inv1  gate3243(.a(G1141), .O(gate425inter8));
  nand2 gate3244(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate3245(.a(s_385), .b(gate425inter3), .O(gate425inter10));
  nor2  gate3246(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate3247(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate3248(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate3095(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate3096(.a(gate426inter0), .b(s_364), .O(gate426inter1));
  and2  gate3097(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate3098(.a(s_364), .O(gate426inter3));
  inv1  gate3099(.a(s_365), .O(gate426inter4));
  nand2 gate3100(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate3101(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate3102(.a(G1045), .O(gate426inter7));
  inv1  gate3103(.a(G1141), .O(gate426inter8));
  nand2 gate3104(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate3105(.a(s_365), .b(gate426inter3), .O(gate426inter10));
  nor2  gate3106(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate3107(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate3108(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1107(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1108(.a(gate427inter0), .b(s_80), .O(gate427inter1));
  and2  gate1109(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1110(.a(s_80), .O(gate427inter3));
  inv1  gate1111(.a(s_81), .O(gate427inter4));
  nand2 gate1112(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1113(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1114(.a(G5), .O(gate427inter7));
  inv1  gate1115(.a(G1144), .O(gate427inter8));
  nand2 gate1116(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1117(.a(s_81), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1118(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1119(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1120(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1835(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1836(.a(gate430inter0), .b(s_184), .O(gate430inter1));
  and2  gate1837(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1838(.a(s_184), .O(gate430inter3));
  inv1  gate1839(.a(s_185), .O(gate430inter4));
  nand2 gate1840(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1841(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1842(.a(G1051), .O(gate430inter7));
  inv1  gate1843(.a(G1147), .O(gate430inter8));
  nand2 gate1844(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1845(.a(s_185), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1846(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1847(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1848(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1583(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1584(.a(gate432inter0), .b(s_148), .O(gate432inter1));
  and2  gate1585(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1586(.a(s_148), .O(gate432inter3));
  inv1  gate1587(.a(s_149), .O(gate432inter4));
  nand2 gate1588(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1589(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1590(.a(G1054), .O(gate432inter7));
  inv1  gate1591(.a(G1150), .O(gate432inter8));
  nand2 gate1592(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1593(.a(s_149), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1594(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1595(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1596(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1793(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1794(.a(gate434inter0), .b(s_178), .O(gate434inter1));
  and2  gate1795(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1796(.a(s_178), .O(gate434inter3));
  inv1  gate1797(.a(s_179), .O(gate434inter4));
  nand2 gate1798(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1799(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1800(.a(G1057), .O(gate434inter7));
  inv1  gate1801(.a(G1153), .O(gate434inter8));
  nand2 gate1802(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1803(.a(s_179), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1804(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1805(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1806(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate869(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate870(.a(gate437inter0), .b(s_46), .O(gate437inter1));
  and2  gate871(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate872(.a(s_46), .O(gate437inter3));
  inv1  gate873(.a(s_47), .O(gate437inter4));
  nand2 gate874(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate875(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate876(.a(G10), .O(gate437inter7));
  inv1  gate877(.a(G1159), .O(gate437inter8));
  nand2 gate878(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate879(.a(s_47), .b(gate437inter3), .O(gate437inter10));
  nor2  gate880(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate881(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate882(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate715(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate716(.a(gate438inter0), .b(s_24), .O(gate438inter1));
  and2  gate717(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate718(.a(s_24), .O(gate438inter3));
  inv1  gate719(.a(s_25), .O(gate438inter4));
  nand2 gate720(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate721(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate722(.a(G1063), .O(gate438inter7));
  inv1  gate723(.a(G1159), .O(gate438inter8));
  nand2 gate724(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate725(.a(s_25), .b(gate438inter3), .O(gate438inter10));
  nor2  gate726(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate727(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate728(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1219(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1220(.a(gate443inter0), .b(s_96), .O(gate443inter1));
  and2  gate1221(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1222(.a(s_96), .O(gate443inter3));
  inv1  gate1223(.a(s_97), .O(gate443inter4));
  nand2 gate1224(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1225(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1226(.a(G13), .O(gate443inter7));
  inv1  gate1227(.a(G1168), .O(gate443inter8));
  nand2 gate1228(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1229(.a(s_97), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1230(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1231(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1232(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2577(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2578(.a(gate448inter0), .b(s_290), .O(gate448inter1));
  and2  gate2579(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2580(.a(s_290), .O(gate448inter3));
  inv1  gate2581(.a(s_291), .O(gate448inter4));
  nand2 gate2582(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2583(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2584(.a(G1078), .O(gate448inter7));
  inv1  gate2585(.a(G1174), .O(gate448inter8));
  nand2 gate2586(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2587(.a(s_291), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2588(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2589(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2590(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate3193(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate3194(.a(gate453inter0), .b(s_378), .O(gate453inter1));
  and2  gate3195(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate3196(.a(s_378), .O(gate453inter3));
  inv1  gate3197(.a(s_379), .O(gate453inter4));
  nand2 gate3198(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate3199(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate3200(.a(G18), .O(gate453inter7));
  inv1  gate3201(.a(G1183), .O(gate453inter8));
  nand2 gate3202(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate3203(.a(s_379), .b(gate453inter3), .O(gate453inter10));
  nor2  gate3204(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate3205(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate3206(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1093(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1094(.a(gate457inter0), .b(s_78), .O(gate457inter1));
  and2  gate1095(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1096(.a(s_78), .O(gate457inter3));
  inv1  gate1097(.a(s_79), .O(gate457inter4));
  nand2 gate1098(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1099(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1100(.a(G20), .O(gate457inter7));
  inv1  gate1101(.a(G1189), .O(gate457inter8));
  nand2 gate1102(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1103(.a(s_79), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1104(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1105(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1106(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2927(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2928(.a(gate459inter0), .b(s_340), .O(gate459inter1));
  and2  gate2929(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2930(.a(s_340), .O(gate459inter3));
  inv1  gate2931(.a(s_341), .O(gate459inter4));
  nand2 gate2932(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2933(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2934(.a(G21), .O(gate459inter7));
  inv1  gate2935(.a(G1192), .O(gate459inter8));
  nand2 gate2936(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2937(.a(s_341), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2938(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2939(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2940(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate3207(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate3208(.a(gate460inter0), .b(s_380), .O(gate460inter1));
  and2  gate3209(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate3210(.a(s_380), .O(gate460inter3));
  inv1  gate3211(.a(s_381), .O(gate460inter4));
  nand2 gate3212(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate3213(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate3214(.a(G1096), .O(gate460inter7));
  inv1  gate3215(.a(G1192), .O(gate460inter8));
  nand2 gate3216(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate3217(.a(s_381), .b(gate460inter3), .O(gate460inter10));
  nor2  gate3218(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate3219(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate3220(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate659(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate660(.a(gate461inter0), .b(s_16), .O(gate461inter1));
  and2  gate661(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate662(.a(s_16), .O(gate461inter3));
  inv1  gate663(.a(s_17), .O(gate461inter4));
  nand2 gate664(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate665(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate666(.a(G22), .O(gate461inter7));
  inv1  gate667(.a(G1195), .O(gate461inter8));
  nand2 gate668(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate669(.a(s_17), .b(gate461inter3), .O(gate461inter10));
  nor2  gate670(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate671(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate672(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate1891(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1892(.a(gate462inter0), .b(s_192), .O(gate462inter1));
  and2  gate1893(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1894(.a(s_192), .O(gate462inter3));
  inv1  gate1895(.a(s_193), .O(gate462inter4));
  nand2 gate1896(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1897(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1898(.a(G1099), .O(gate462inter7));
  inv1  gate1899(.a(G1195), .O(gate462inter8));
  nand2 gate1900(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1901(.a(s_193), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1902(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1903(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1904(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1037(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1038(.a(gate463inter0), .b(s_70), .O(gate463inter1));
  and2  gate1039(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1040(.a(s_70), .O(gate463inter3));
  inv1  gate1041(.a(s_71), .O(gate463inter4));
  nand2 gate1042(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1043(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1044(.a(G23), .O(gate463inter7));
  inv1  gate1045(.a(G1198), .O(gate463inter8));
  nand2 gate1046(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1047(.a(s_71), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1048(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1049(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1050(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1359(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1360(.a(gate465inter0), .b(s_116), .O(gate465inter1));
  and2  gate1361(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1362(.a(s_116), .O(gate465inter3));
  inv1  gate1363(.a(s_117), .O(gate465inter4));
  nand2 gate1364(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1365(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1366(.a(G24), .O(gate465inter7));
  inv1  gate1367(.a(G1201), .O(gate465inter8));
  nand2 gate1368(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1369(.a(s_117), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1370(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1371(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1372(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1023(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1024(.a(gate466inter0), .b(s_68), .O(gate466inter1));
  and2  gate1025(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1026(.a(s_68), .O(gate466inter3));
  inv1  gate1027(.a(s_69), .O(gate466inter4));
  nand2 gate1028(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1029(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1030(.a(G1105), .O(gate466inter7));
  inv1  gate1031(.a(G1201), .O(gate466inter8));
  nand2 gate1032(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1033(.a(s_69), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1034(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1035(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1036(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate3151(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate3152(.a(gate471inter0), .b(s_372), .O(gate471inter1));
  and2  gate3153(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate3154(.a(s_372), .O(gate471inter3));
  inv1  gate3155(.a(s_373), .O(gate471inter4));
  nand2 gate3156(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate3157(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate3158(.a(G27), .O(gate471inter7));
  inv1  gate3159(.a(G1210), .O(gate471inter8));
  nand2 gate3160(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate3161(.a(s_373), .b(gate471inter3), .O(gate471inter10));
  nor2  gate3162(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate3163(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate3164(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate757(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate758(.a(gate472inter0), .b(s_30), .O(gate472inter1));
  and2  gate759(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate760(.a(s_30), .O(gate472inter3));
  inv1  gate761(.a(s_31), .O(gate472inter4));
  nand2 gate762(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate763(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate764(.a(G1114), .O(gate472inter7));
  inv1  gate765(.a(G1210), .O(gate472inter8));
  nand2 gate766(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate767(.a(s_31), .b(gate472inter3), .O(gate472inter10));
  nor2  gate768(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate769(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate770(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate617(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate618(.a(gate474inter0), .b(s_10), .O(gate474inter1));
  and2  gate619(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate620(.a(s_10), .O(gate474inter3));
  inv1  gate621(.a(s_11), .O(gate474inter4));
  nand2 gate622(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate623(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate624(.a(G1117), .O(gate474inter7));
  inv1  gate625(.a(G1213), .O(gate474inter8));
  nand2 gate626(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate627(.a(s_11), .b(gate474inter3), .O(gate474inter10));
  nor2  gate628(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate629(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate630(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate645(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate646(.a(gate475inter0), .b(s_14), .O(gate475inter1));
  and2  gate647(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate648(.a(s_14), .O(gate475inter3));
  inv1  gate649(.a(s_15), .O(gate475inter4));
  nand2 gate650(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate651(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate652(.a(G29), .O(gate475inter7));
  inv1  gate653(.a(G1216), .O(gate475inter8));
  nand2 gate654(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate655(.a(s_15), .b(gate475inter3), .O(gate475inter10));
  nor2  gate656(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate657(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate658(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1625(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1626(.a(gate478inter0), .b(s_154), .O(gate478inter1));
  and2  gate1627(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1628(.a(s_154), .O(gate478inter3));
  inv1  gate1629(.a(s_155), .O(gate478inter4));
  nand2 gate1630(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1631(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1632(.a(G1123), .O(gate478inter7));
  inv1  gate1633(.a(G1219), .O(gate478inter8));
  nand2 gate1634(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1635(.a(s_155), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1636(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1637(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1638(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2339(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2340(.a(gate479inter0), .b(s_256), .O(gate479inter1));
  and2  gate2341(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2342(.a(s_256), .O(gate479inter3));
  inv1  gate2343(.a(s_257), .O(gate479inter4));
  nand2 gate2344(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2345(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2346(.a(G31), .O(gate479inter7));
  inv1  gate2347(.a(G1222), .O(gate479inter8));
  nand2 gate2348(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2349(.a(s_257), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2350(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2351(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2352(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1695(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1696(.a(gate481inter0), .b(s_164), .O(gate481inter1));
  and2  gate1697(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1698(.a(s_164), .O(gate481inter3));
  inv1  gate1699(.a(s_165), .O(gate481inter4));
  nand2 gate1700(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1701(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1702(.a(G32), .O(gate481inter7));
  inv1  gate1703(.a(G1225), .O(gate481inter8));
  nand2 gate1704(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1705(.a(s_165), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1706(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1707(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1708(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate2031(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2032(.a(gate482inter0), .b(s_212), .O(gate482inter1));
  and2  gate2033(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2034(.a(s_212), .O(gate482inter3));
  inv1  gate2035(.a(s_213), .O(gate482inter4));
  nand2 gate2036(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2037(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2038(.a(G1129), .O(gate482inter7));
  inv1  gate2039(.a(G1225), .O(gate482inter8));
  nand2 gate2040(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2041(.a(s_213), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2042(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2043(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2044(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1877(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1878(.a(gate483inter0), .b(s_190), .O(gate483inter1));
  and2  gate1879(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1880(.a(s_190), .O(gate483inter3));
  inv1  gate1881(.a(s_191), .O(gate483inter4));
  nand2 gate1882(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1883(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1884(.a(G1228), .O(gate483inter7));
  inv1  gate1885(.a(G1229), .O(gate483inter8));
  nand2 gate1886(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1887(.a(s_191), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1888(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1889(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1890(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate2647(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2648(.a(gate487inter0), .b(s_300), .O(gate487inter1));
  and2  gate2649(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2650(.a(s_300), .O(gate487inter3));
  inv1  gate2651(.a(s_301), .O(gate487inter4));
  nand2 gate2652(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2653(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2654(.a(G1236), .O(gate487inter7));
  inv1  gate2655(.a(G1237), .O(gate487inter8));
  nand2 gate2656(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2657(.a(s_301), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2658(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2659(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2660(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1443(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1444(.a(gate489inter0), .b(s_128), .O(gate489inter1));
  and2  gate1445(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1446(.a(s_128), .O(gate489inter3));
  inv1  gate1447(.a(s_129), .O(gate489inter4));
  nand2 gate1448(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1449(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1450(.a(G1240), .O(gate489inter7));
  inv1  gate1451(.a(G1241), .O(gate489inter8));
  nand2 gate1452(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1453(.a(s_129), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1454(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1455(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1456(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1387(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1388(.a(gate491inter0), .b(s_120), .O(gate491inter1));
  and2  gate1389(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1390(.a(s_120), .O(gate491inter3));
  inv1  gate1391(.a(s_121), .O(gate491inter4));
  nand2 gate1392(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1393(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1394(.a(G1244), .O(gate491inter7));
  inv1  gate1395(.a(G1245), .O(gate491inter8));
  nand2 gate1396(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1397(.a(s_121), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1398(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1399(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1400(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate2983(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2984(.a(gate492inter0), .b(s_348), .O(gate492inter1));
  and2  gate2985(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2986(.a(s_348), .O(gate492inter3));
  inv1  gate2987(.a(s_349), .O(gate492inter4));
  nand2 gate2988(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2989(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2990(.a(G1246), .O(gate492inter7));
  inv1  gate2991(.a(G1247), .O(gate492inter8));
  nand2 gate2992(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2993(.a(s_349), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2994(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2995(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2996(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2689(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2690(.a(gate493inter0), .b(s_306), .O(gate493inter1));
  and2  gate2691(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2692(.a(s_306), .O(gate493inter3));
  inv1  gate2693(.a(s_307), .O(gate493inter4));
  nand2 gate2694(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2695(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2696(.a(G1248), .O(gate493inter7));
  inv1  gate2697(.a(G1249), .O(gate493inter8));
  nand2 gate2698(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2699(.a(s_307), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2700(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2701(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2702(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1233(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1234(.a(gate494inter0), .b(s_98), .O(gate494inter1));
  and2  gate1235(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1236(.a(s_98), .O(gate494inter3));
  inv1  gate1237(.a(s_99), .O(gate494inter4));
  nand2 gate1238(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1239(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1240(.a(G1250), .O(gate494inter7));
  inv1  gate1241(.a(G1251), .O(gate494inter8));
  nand2 gate1242(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1243(.a(s_99), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1244(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1245(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1246(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate631(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate632(.a(gate498inter0), .b(s_12), .O(gate498inter1));
  and2  gate633(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate634(.a(s_12), .O(gate498inter3));
  inv1  gate635(.a(s_13), .O(gate498inter4));
  nand2 gate636(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate637(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate638(.a(G1258), .O(gate498inter7));
  inv1  gate639(.a(G1259), .O(gate498inter8));
  nand2 gate640(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate641(.a(s_13), .b(gate498inter3), .O(gate498inter10));
  nor2  gate642(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate643(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate644(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate2451(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2452(.a(gate499inter0), .b(s_272), .O(gate499inter1));
  and2  gate2453(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2454(.a(s_272), .O(gate499inter3));
  inv1  gate2455(.a(s_273), .O(gate499inter4));
  nand2 gate2456(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2457(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2458(.a(G1260), .O(gate499inter7));
  inv1  gate2459(.a(G1261), .O(gate499inter8));
  nand2 gate2460(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2461(.a(s_273), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2462(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2463(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2464(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate729(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate730(.a(gate500inter0), .b(s_26), .O(gate500inter1));
  and2  gate731(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate732(.a(s_26), .O(gate500inter3));
  inv1  gate733(.a(s_27), .O(gate500inter4));
  nand2 gate734(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate735(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate736(.a(G1262), .O(gate500inter7));
  inv1  gate737(.a(G1263), .O(gate500inter8));
  nand2 gate738(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate739(.a(s_27), .b(gate500inter3), .O(gate500inter10));
  nor2  gate740(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate741(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate742(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2829(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2830(.a(gate501inter0), .b(s_326), .O(gate501inter1));
  and2  gate2831(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2832(.a(s_326), .O(gate501inter3));
  inv1  gate2833(.a(s_327), .O(gate501inter4));
  nand2 gate2834(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2835(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2836(.a(G1264), .O(gate501inter7));
  inv1  gate2837(.a(G1265), .O(gate501inter8));
  nand2 gate2838(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2839(.a(s_327), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2840(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2841(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2842(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1765(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1766(.a(gate502inter0), .b(s_174), .O(gate502inter1));
  and2  gate1767(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1768(.a(s_174), .O(gate502inter3));
  inv1  gate1769(.a(s_175), .O(gate502inter4));
  nand2 gate1770(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1771(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1772(.a(G1266), .O(gate502inter7));
  inv1  gate1773(.a(G1267), .O(gate502inter8));
  nand2 gate1774(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1775(.a(s_175), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1776(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1777(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1778(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1653(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1654(.a(gate503inter0), .b(s_158), .O(gate503inter1));
  and2  gate1655(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1656(.a(s_158), .O(gate503inter3));
  inv1  gate1657(.a(s_159), .O(gate503inter4));
  nand2 gate1658(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1659(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1660(.a(G1268), .O(gate503inter7));
  inv1  gate1661(.a(G1269), .O(gate503inter8));
  nand2 gate1662(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1663(.a(s_159), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1664(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1665(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1666(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate799(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate800(.a(gate505inter0), .b(s_36), .O(gate505inter1));
  and2  gate801(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate802(.a(s_36), .O(gate505inter3));
  inv1  gate803(.a(s_37), .O(gate505inter4));
  nand2 gate804(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate805(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate806(.a(G1272), .O(gate505inter7));
  inv1  gate807(.a(G1273), .O(gate505inter8));
  nand2 gate808(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate809(.a(s_37), .b(gate505inter3), .O(gate505inter10));
  nor2  gate810(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate811(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate812(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1975(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1976(.a(gate506inter0), .b(s_204), .O(gate506inter1));
  and2  gate1977(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1978(.a(s_204), .O(gate506inter3));
  inv1  gate1979(.a(s_205), .O(gate506inter4));
  nand2 gate1980(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1981(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1982(.a(G1274), .O(gate506inter7));
  inv1  gate1983(.a(G1275), .O(gate506inter8));
  nand2 gate1984(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1985(.a(s_205), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1986(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1987(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1988(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2045(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2046(.a(gate511inter0), .b(s_214), .O(gate511inter1));
  and2  gate2047(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2048(.a(s_214), .O(gate511inter3));
  inv1  gate2049(.a(s_215), .O(gate511inter4));
  nand2 gate2050(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2051(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2052(.a(G1284), .O(gate511inter7));
  inv1  gate2053(.a(G1285), .O(gate511inter8));
  nand2 gate2054(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2055(.a(s_215), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2056(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2057(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2058(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2255(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2256(.a(gate513inter0), .b(s_244), .O(gate513inter1));
  and2  gate2257(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2258(.a(s_244), .O(gate513inter3));
  inv1  gate2259(.a(s_245), .O(gate513inter4));
  nand2 gate2260(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2261(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2262(.a(G1288), .O(gate513inter7));
  inv1  gate2263(.a(G1289), .O(gate513inter8));
  nand2 gate2264(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2265(.a(s_245), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2266(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2267(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2268(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate2759(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2760(.a(gate514inter0), .b(s_316), .O(gate514inter1));
  and2  gate2761(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2762(.a(s_316), .O(gate514inter3));
  inv1  gate2763(.a(s_317), .O(gate514inter4));
  nand2 gate2764(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2765(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2766(.a(G1290), .O(gate514inter7));
  inv1  gate2767(.a(G1291), .O(gate514inter8));
  nand2 gate2768(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2769(.a(s_317), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2770(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2771(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2772(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule