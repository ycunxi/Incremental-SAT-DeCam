module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2801(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2802(.a(gate15inter0), .b(s_322), .O(gate15inter1));
  and2  gate2803(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2804(.a(s_322), .O(gate15inter3));
  inv1  gate2805(.a(s_323), .O(gate15inter4));
  nand2 gate2806(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2807(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2808(.a(G13), .O(gate15inter7));
  inv1  gate2809(.a(G14), .O(gate15inter8));
  nand2 gate2810(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2811(.a(s_323), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2812(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2813(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2814(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2073(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2074(.a(gate16inter0), .b(s_218), .O(gate16inter1));
  and2  gate2075(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2076(.a(s_218), .O(gate16inter3));
  inv1  gate2077(.a(s_219), .O(gate16inter4));
  nand2 gate2078(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2079(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2080(.a(G15), .O(gate16inter7));
  inv1  gate2081(.a(G16), .O(gate16inter8));
  nand2 gate2082(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2083(.a(s_219), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2084(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2085(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2086(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate799(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate800(.a(gate17inter0), .b(s_36), .O(gate17inter1));
  and2  gate801(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate802(.a(s_36), .O(gate17inter3));
  inv1  gate803(.a(s_37), .O(gate17inter4));
  nand2 gate804(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate805(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate806(.a(G17), .O(gate17inter7));
  inv1  gate807(.a(G18), .O(gate17inter8));
  nand2 gate808(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate809(.a(s_37), .b(gate17inter3), .O(gate17inter10));
  nor2  gate810(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate811(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate812(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1303(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1304(.a(gate20inter0), .b(s_108), .O(gate20inter1));
  and2  gate1305(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1306(.a(s_108), .O(gate20inter3));
  inv1  gate1307(.a(s_109), .O(gate20inter4));
  nand2 gate1308(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1309(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1310(.a(G23), .O(gate20inter7));
  inv1  gate1311(.a(G24), .O(gate20inter8));
  nand2 gate1312(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1313(.a(s_109), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1314(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1315(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1316(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1583(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1584(.a(gate22inter0), .b(s_148), .O(gate22inter1));
  and2  gate1585(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1586(.a(s_148), .O(gate22inter3));
  inv1  gate1587(.a(s_149), .O(gate22inter4));
  nand2 gate1588(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1589(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1590(.a(G27), .O(gate22inter7));
  inv1  gate1591(.a(G28), .O(gate22inter8));
  nand2 gate1592(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1593(.a(s_149), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1594(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1595(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1596(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1191(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1192(.a(gate24inter0), .b(s_92), .O(gate24inter1));
  and2  gate1193(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1194(.a(s_92), .O(gate24inter3));
  inv1  gate1195(.a(s_93), .O(gate24inter4));
  nand2 gate1196(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1197(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1198(.a(G31), .O(gate24inter7));
  inv1  gate1199(.a(G32), .O(gate24inter8));
  nand2 gate1200(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1201(.a(s_93), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1202(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1203(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1204(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2731(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2732(.a(gate26inter0), .b(s_312), .O(gate26inter1));
  and2  gate2733(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2734(.a(s_312), .O(gate26inter3));
  inv1  gate2735(.a(s_313), .O(gate26inter4));
  nand2 gate2736(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2737(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2738(.a(G9), .O(gate26inter7));
  inv1  gate2739(.a(G13), .O(gate26inter8));
  nand2 gate2740(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2741(.a(s_313), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2742(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2743(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2744(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2591(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2592(.a(gate28inter0), .b(s_292), .O(gate28inter1));
  and2  gate2593(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2594(.a(s_292), .O(gate28inter3));
  inv1  gate2595(.a(s_293), .O(gate28inter4));
  nand2 gate2596(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2597(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2598(.a(G10), .O(gate28inter7));
  inv1  gate2599(.a(G14), .O(gate28inter8));
  nand2 gate2600(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2601(.a(s_293), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2602(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2603(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2604(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2493(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2494(.a(gate32inter0), .b(s_278), .O(gate32inter1));
  and2  gate2495(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2496(.a(s_278), .O(gate32inter3));
  inv1  gate2497(.a(s_279), .O(gate32inter4));
  nand2 gate2498(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2499(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2500(.a(G12), .O(gate32inter7));
  inv1  gate2501(.a(G16), .O(gate32inter8));
  nand2 gate2502(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2503(.a(s_279), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2504(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2505(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2506(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1919(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1920(.a(gate37inter0), .b(s_196), .O(gate37inter1));
  and2  gate1921(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1922(.a(s_196), .O(gate37inter3));
  inv1  gate1923(.a(s_197), .O(gate37inter4));
  nand2 gate1924(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1925(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1926(.a(G19), .O(gate37inter7));
  inv1  gate1927(.a(G23), .O(gate37inter8));
  nand2 gate1928(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1929(.a(s_197), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1930(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1931(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1932(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2675(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2676(.a(gate39inter0), .b(s_304), .O(gate39inter1));
  and2  gate2677(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2678(.a(s_304), .O(gate39inter3));
  inv1  gate2679(.a(s_305), .O(gate39inter4));
  nand2 gate2680(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2681(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2682(.a(G20), .O(gate39inter7));
  inv1  gate2683(.a(G24), .O(gate39inter8));
  nand2 gate2684(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2685(.a(s_305), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2686(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2687(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2688(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1275(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1276(.a(gate42inter0), .b(s_104), .O(gate42inter1));
  and2  gate1277(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1278(.a(s_104), .O(gate42inter3));
  inv1  gate1279(.a(s_105), .O(gate42inter4));
  nand2 gate1280(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1281(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1282(.a(G2), .O(gate42inter7));
  inv1  gate1283(.a(G266), .O(gate42inter8));
  nand2 gate1284(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1285(.a(s_105), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1286(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1287(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1288(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1835(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1836(.a(gate43inter0), .b(s_184), .O(gate43inter1));
  and2  gate1837(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1838(.a(s_184), .O(gate43inter3));
  inv1  gate1839(.a(s_185), .O(gate43inter4));
  nand2 gate1840(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1841(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1842(.a(G3), .O(gate43inter7));
  inv1  gate1843(.a(G269), .O(gate43inter8));
  nand2 gate1844(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1845(.a(s_185), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1846(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1847(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1848(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1527(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1528(.a(gate44inter0), .b(s_140), .O(gate44inter1));
  and2  gate1529(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1530(.a(s_140), .O(gate44inter3));
  inv1  gate1531(.a(s_141), .O(gate44inter4));
  nand2 gate1532(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1533(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1534(.a(G4), .O(gate44inter7));
  inv1  gate1535(.a(G269), .O(gate44inter8));
  nand2 gate1536(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1537(.a(s_141), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1538(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1539(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1540(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1653(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1654(.a(gate48inter0), .b(s_158), .O(gate48inter1));
  and2  gate1655(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1656(.a(s_158), .O(gate48inter3));
  inv1  gate1657(.a(s_159), .O(gate48inter4));
  nand2 gate1658(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1659(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1660(.a(G8), .O(gate48inter7));
  inv1  gate1661(.a(G275), .O(gate48inter8));
  nand2 gate1662(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1663(.a(s_159), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1664(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1665(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1666(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1695(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1696(.a(gate50inter0), .b(s_164), .O(gate50inter1));
  and2  gate1697(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1698(.a(s_164), .O(gate50inter3));
  inv1  gate1699(.a(s_165), .O(gate50inter4));
  nand2 gate1700(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1701(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1702(.a(G10), .O(gate50inter7));
  inv1  gate1703(.a(G278), .O(gate50inter8));
  nand2 gate1704(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1705(.a(s_165), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1706(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1707(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1708(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate939(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate940(.a(gate54inter0), .b(s_56), .O(gate54inter1));
  and2  gate941(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate942(.a(s_56), .O(gate54inter3));
  inv1  gate943(.a(s_57), .O(gate54inter4));
  nand2 gate944(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate945(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate946(.a(G14), .O(gate54inter7));
  inv1  gate947(.a(G284), .O(gate54inter8));
  nand2 gate948(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate949(.a(s_57), .b(gate54inter3), .O(gate54inter10));
  nor2  gate950(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate951(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate952(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1863(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1864(.a(gate55inter0), .b(s_188), .O(gate55inter1));
  and2  gate1865(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1866(.a(s_188), .O(gate55inter3));
  inv1  gate1867(.a(s_189), .O(gate55inter4));
  nand2 gate1868(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1869(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1870(.a(G15), .O(gate55inter7));
  inv1  gate1871(.a(G287), .O(gate55inter8));
  nand2 gate1872(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1873(.a(s_189), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1874(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1875(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1876(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate2395(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2396(.a(gate57inter0), .b(s_264), .O(gate57inter1));
  and2  gate2397(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2398(.a(s_264), .O(gate57inter3));
  inv1  gate2399(.a(s_265), .O(gate57inter4));
  nand2 gate2400(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2401(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2402(.a(G17), .O(gate57inter7));
  inv1  gate2403(.a(G290), .O(gate57inter8));
  nand2 gate2404(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2405(.a(s_265), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2406(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2407(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2408(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2619(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2620(.a(gate60inter0), .b(s_296), .O(gate60inter1));
  and2  gate2621(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2622(.a(s_296), .O(gate60inter3));
  inv1  gate2623(.a(s_297), .O(gate60inter4));
  nand2 gate2624(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2625(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2626(.a(G20), .O(gate60inter7));
  inv1  gate2627(.a(G293), .O(gate60inter8));
  nand2 gate2628(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2629(.a(s_297), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2630(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2631(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2632(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1765(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1766(.a(gate61inter0), .b(s_174), .O(gate61inter1));
  and2  gate1767(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1768(.a(s_174), .O(gate61inter3));
  inv1  gate1769(.a(s_175), .O(gate61inter4));
  nand2 gate1770(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1771(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1772(.a(G21), .O(gate61inter7));
  inv1  gate1773(.a(G296), .O(gate61inter8));
  nand2 gate1774(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1775(.a(s_175), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1776(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1777(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1778(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1163(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1164(.a(gate62inter0), .b(s_88), .O(gate62inter1));
  and2  gate1165(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1166(.a(s_88), .O(gate62inter3));
  inv1  gate1167(.a(s_89), .O(gate62inter4));
  nand2 gate1168(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1169(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1170(.a(G22), .O(gate62inter7));
  inv1  gate1171(.a(G296), .O(gate62inter8));
  nand2 gate1172(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1173(.a(s_89), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1174(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1175(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1176(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1177(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1178(.a(gate64inter0), .b(s_90), .O(gate64inter1));
  and2  gate1179(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1180(.a(s_90), .O(gate64inter3));
  inv1  gate1181(.a(s_91), .O(gate64inter4));
  nand2 gate1182(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1183(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1184(.a(G24), .O(gate64inter7));
  inv1  gate1185(.a(G299), .O(gate64inter8));
  nand2 gate1186(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1187(.a(s_91), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1188(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1189(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1190(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate645(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate646(.a(gate68inter0), .b(s_14), .O(gate68inter1));
  and2  gate647(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate648(.a(s_14), .O(gate68inter3));
  inv1  gate649(.a(s_15), .O(gate68inter4));
  nand2 gate650(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate651(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate652(.a(G28), .O(gate68inter7));
  inv1  gate653(.a(G305), .O(gate68inter8));
  nand2 gate654(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate655(.a(s_15), .b(gate68inter3), .O(gate68inter10));
  nor2  gate656(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate657(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate658(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2871(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2872(.a(gate72inter0), .b(s_332), .O(gate72inter1));
  and2  gate2873(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2874(.a(s_332), .O(gate72inter3));
  inv1  gate2875(.a(s_333), .O(gate72inter4));
  nand2 gate2876(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2877(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2878(.a(G32), .O(gate72inter7));
  inv1  gate2879(.a(G311), .O(gate72inter8));
  nand2 gate2880(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2881(.a(s_333), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2882(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2883(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2884(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate911(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate912(.a(gate73inter0), .b(s_52), .O(gate73inter1));
  and2  gate913(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate914(.a(s_52), .O(gate73inter3));
  inv1  gate915(.a(s_53), .O(gate73inter4));
  nand2 gate916(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate917(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate918(.a(G1), .O(gate73inter7));
  inv1  gate919(.a(G314), .O(gate73inter8));
  nand2 gate920(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate921(.a(s_53), .b(gate73inter3), .O(gate73inter10));
  nor2  gate922(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate923(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate924(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2003(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2004(.a(gate76inter0), .b(s_208), .O(gate76inter1));
  and2  gate2005(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2006(.a(s_208), .O(gate76inter3));
  inv1  gate2007(.a(s_209), .O(gate76inter4));
  nand2 gate2008(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2009(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2010(.a(G13), .O(gate76inter7));
  inv1  gate2011(.a(G317), .O(gate76inter8));
  nand2 gate2012(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2013(.a(s_209), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2014(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2015(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2016(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1639(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1640(.a(gate78inter0), .b(s_156), .O(gate78inter1));
  and2  gate1641(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1642(.a(s_156), .O(gate78inter3));
  inv1  gate1643(.a(s_157), .O(gate78inter4));
  nand2 gate1644(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1645(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1646(.a(G6), .O(gate78inter7));
  inv1  gate1647(.a(G320), .O(gate78inter8));
  nand2 gate1648(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1649(.a(s_157), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1650(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1651(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1652(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2199(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2200(.a(gate79inter0), .b(s_236), .O(gate79inter1));
  and2  gate2201(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2202(.a(s_236), .O(gate79inter3));
  inv1  gate2203(.a(s_237), .O(gate79inter4));
  nand2 gate2204(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2205(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2206(.a(G10), .O(gate79inter7));
  inv1  gate2207(.a(G323), .O(gate79inter8));
  nand2 gate2208(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2209(.a(s_237), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2210(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2211(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2212(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1989(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1990(.a(gate82inter0), .b(s_206), .O(gate82inter1));
  and2  gate1991(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1992(.a(s_206), .O(gate82inter3));
  inv1  gate1993(.a(s_207), .O(gate82inter4));
  nand2 gate1994(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1995(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1996(.a(G7), .O(gate82inter7));
  inv1  gate1997(.a(G326), .O(gate82inter8));
  nand2 gate1998(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1999(.a(s_207), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2000(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2001(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2002(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1219(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1220(.a(gate83inter0), .b(s_96), .O(gate83inter1));
  and2  gate1221(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1222(.a(s_96), .O(gate83inter3));
  inv1  gate1223(.a(s_97), .O(gate83inter4));
  nand2 gate1224(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1225(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1226(.a(G11), .O(gate83inter7));
  inv1  gate1227(.a(G329), .O(gate83inter8));
  nand2 gate1228(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1229(.a(s_97), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1230(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1231(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1232(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1891(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1892(.a(gate85inter0), .b(s_192), .O(gate85inter1));
  and2  gate1893(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1894(.a(s_192), .O(gate85inter3));
  inv1  gate1895(.a(s_193), .O(gate85inter4));
  nand2 gate1896(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1897(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1898(.a(G4), .O(gate85inter7));
  inv1  gate1899(.a(G332), .O(gate85inter8));
  nand2 gate1900(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1901(.a(s_193), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1902(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1903(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1904(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2759(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2760(.a(gate87inter0), .b(s_316), .O(gate87inter1));
  and2  gate2761(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2762(.a(s_316), .O(gate87inter3));
  inv1  gate2763(.a(s_317), .O(gate87inter4));
  nand2 gate2764(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2765(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2766(.a(G12), .O(gate87inter7));
  inv1  gate2767(.a(G335), .O(gate87inter8));
  nand2 gate2768(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2769(.a(s_317), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2770(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2771(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2772(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1569(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1570(.a(gate93inter0), .b(s_146), .O(gate93inter1));
  and2  gate1571(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1572(.a(s_146), .O(gate93inter3));
  inv1  gate1573(.a(s_147), .O(gate93inter4));
  nand2 gate1574(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1575(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1576(.a(G18), .O(gate93inter7));
  inv1  gate1577(.a(G344), .O(gate93inter8));
  nand2 gate1578(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1579(.a(s_147), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1580(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1581(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1582(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1961(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1962(.a(gate94inter0), .b(s_202), .O(gate94inter1));
  and2  gate1963(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1964(.a(s_202), .O(gate94inter3));
  inv1  gate1965(.a(s_203), .O(gate94inter4));
  nand2 gate1966(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1967(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1968(.a(G22), .O(gate94inter7));
  inv1  gate1969(.a(G344), .O(gate94inter8));
  nand2 gate1970(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1971(.a(s_203), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1972(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1973(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1974(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1149(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1150(.a(gate95inter0), .b(s_86), .O(gate95inter1));
  and2  gate1151(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1152(.a(s_86), .O(gate95inter3));
  inv1  gate1153(.a(s_87), .O(gate95inter4));
  nand2 gate1154(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1155(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1156(.a(G26), .O(gate95inter7));
  inv1  gate1157(.a(G347), .O(gate95inter8));
  nand2 gate1158(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1159(.a(s_87), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1160(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1161(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1162(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2311(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2312(.a(gate100inter0), .b(s_252), .O(gate100inter1));
  and2  gate2313(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2314(.a(s_252), .O(gate100inter3));
  inv1  gate2315(.a(s_253), .O(gate100inter4));
  nand2 gate2316(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2317(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2318(.a(G31), .O(gate100inter7));
  inv1  gate2319(.a(G353), .O(gate100inter8));
  nand2 gate2320(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2321(.a(s_253), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2322(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2323(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2324(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1079(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1080(.a(gate101inter0), .b(s_76), .O(gate101inter1));
  and2  gate1081(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1082(.a(s_76), .O(gate101inter3));
  inv1  gate1083(.a(s_77), .O(gate101inter4));
  nand2 gate1084(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1085(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1086(.a(G20), .O(gate101inter7));
  inv1  gate1087(.a(G356), .O(gate101inter8));
  nand2 gate1088(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1089(.a(s_77), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1090(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1091(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1092(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate715(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate716(.a(gate102inter0), .b(s_24), .O(gate102inter1));
  and2  gate717(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate718(.a(s_24), .O(gate102inter3));
  inv1  gate719(.a(s_25), .O(gate102inter4));
  nand2 gate720(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate721(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate722(.a(G24), .O(gate102inter7));
  inv1  gate723(.a(G356), .O(gate102inter8));
  nand2 gate724(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate725(.a(s_25), .b(gate102inter3), .O(gate102inter10));
  nor2  gate726(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate727(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate728(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate2465(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2466(.a(gate103inter0), .b(s_274), .O(gate103inter1));
  and2  gate2467(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2468(.a(s_274), .O(gate103inter3));
  inv1  gate2469(.a(s_275), .O(gate103inter4));
  nand2 gate2470(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2471(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2472(.a(G28), .O(gate103inter7));
  inv1  gate2473(.a(G359), .O(gate103inter8));
  nand2 gate2474(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2475(.a(s_275), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2476(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2477(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2478(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1051(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1052(.a(gate106inter0), .b(s_72), .O(gate106inter1));
  and2  gate1053(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1054(.a(s_72), .O(gate106inter3));
  inv1  gate1055(.a(s_73), .O(gate106inter4));
  nand2 gate1056(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1057(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1058(.a(G364), .O(gate106inter7));
  inv1  gate1059(.a(G365), .O(gate106inter8));
  nand2 gate1060(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1061(.a(s_73), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1062(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1063(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1064(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2255(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2256(.a(gate108inter0), .b(s_244), .O(gate108inter1));
  and2  gate2257(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2258(.a(s_244), .O(gate108inter3));
  inv1  gate2259(.a(s_245), .O(gate108inter4));
  nand2 gate2260(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2261(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2262(.a(G368), .O(gate108inter7));
  inv1  gate2263(.a(G369), .O(gate108inter8));
  nand2 gate2264(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2265(.a(s_245), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2266(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2267(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2268(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2563(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2564(.a(gate112inter0), .b(s_288), .O(gate112inter1));
  and2  gate2565(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2566(.a(s_288), .O(gate112inter3));
  inv1  gate2567(.a(s_289), .O(gate112inter4));
  nand2 gate2568(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2569(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2570(.a(G376), .O(gate112inter7));
  inv1  gate2571(.a(G377), .O(gate112inter8));
  nand2 gate2572(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2573(.a(s_289), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2574(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2575(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2576(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2913(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2914(.a(gate115inter0), .b(s_338), .O(gate115inter1));
  and2  gate2915(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2916(.a(s_338), .O(gate115inter3));
  inv1  gate2917(.a(s_339), .O(gate115inter4));
  nand2 gate2918(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2919(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2920(.a(G382), .O(gate115inter7));
  inv1  gate2921(.a(G383), .O(gate115inter8));
  nand2 gate2922(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2923(.a(s_339), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2924(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2925(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2926(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate897(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate898(.a(gate122inter0), .b(s_50), .O(gate122inter1));
  and2  gate899(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate900(.a(s_50), .O(gate122inter3));
  inv1  gate901(.a(s_51), .O(gate122inter4));
  nand2 gate902(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate903(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate904(.a(G396), .O(gate122inter7));
  inv1  gate905(.a(G397), .O(gate122inter8));
  nand2 gate906(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate907(.a(s_51), .b(gate122inter3), .O(gate122inter10));
  nor2  gate908(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate909(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate910(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate659(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate660(.a(gate126inter0), .b(s_16), .O(gate126inter1));
  and2  gate661(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate662(.a(s_16), .O(gate126inter3));
  inv1  gate663(.a(s_17), .O(gate126inter4));
  nand2 gate664(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate665(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate666(.a(G404), .O(gate126inter7));
  inv1  gate667(.a(G405), .O(gate126inter8));
  nand2 gate668(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate669(.a(s_17), .b(gate126inter3), .O(gate126inter10));
  nor2  gate670(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate671(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate672(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2157(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2158(.a(gate128inter0), .b(s_230), .O(gate128inter1));
  and2  gate2159(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2160(.a(s_230), .O(gate128inter3));
  inv1  gate2161(.a(s_231), .O(gate128inter4));
  nand2 gate2162(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2163(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2164(.a(G408), .O(gate128inter7));
  inv1  gate2165(.a(G409), .O(gate128inter8));
  nand2 gate2166(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2167(.a(s_231), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2168(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2169(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2170(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate925(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate926(.a(gate132inter0), .b(s_54), .O(gate132inter1));
  and2  gate927(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate928(.a(s_54), .O(gate132inter3));
  inv1  gate929(.a(s_55), .O(gate132inter4));
  nand2 gate930(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate931(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate932(.a(G416), .O(gate132inter7));
  inv1  gate933(.a(G417), .O(gate132inter8));
  nand2 gate934(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate935(.a(s_55), .b(gate132inter3), .O(gate132inter10));
  nor2  gate936(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate937(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate938(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1681(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1682(.a(gate133inter0), .b(s_162), .O(gate133inter1));
  and2  gate1683(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1684(.a(s_162), .O(gate133inter3));
  inv1  gate1685(.a(s_163), .O(gate133inter4));
  nand2 gate1686(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1687(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1688(.a(G418), .O(gate133inter7));
  inv1  gate1689(.a(G419), .O(gate133inter8));
  nand2 gate1690(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1691(.a(s_163), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1692(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1693(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1694(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1597(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1598(.a(gate134inter0), .b(s_150), .O(gate134inter1));
  and2  gate1599(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1600(.a(s_150), .O(gate134inter3));
  inv1  gate1601(.a(s_151), .O(gate134inter4));
  nand2 gate1602(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1603(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1604(.a(G420), .O(gate134inter7));
  inv1  gate1605(.a(G421), .O(gate134inter8));
  nand2 gate1606(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1607(.a(s_151), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1608(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1609(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1610(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate617(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate618(.a(gate140inter0), .b(s_10), .O(gate140inter1));
  and2  gate619(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate620(.a(s_10), .O(gate140inter3));
  inv1  gate621(.a(s_11), .O(gate140inter4));
  nand2 gate622(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate623(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate624(.a(G444), .O(gate140inter7));
  inv1  gate625(.a(G447), .O(gate140inter8));
  nand2 gate626(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate627(.a(s_11), .b(gate140inter3), .O(gate140inter10));
  nor2  gate628(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate629(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate630(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1359(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1360(.a(gate143inter0), .b(s_116), .O(gate143inter1));
  and2  gate1361(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1362(.a(s_116), .O(gate143inter3));
  inv1  gate1363(.a(s_117), .O(gate143inter4));
  nand2 gate1364(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1365(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1366(.a(G462), .O(gate143inter7));
  inv1  gate1367(.a(G465), .O(gate143inter8));
  nand2 gate1368(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1369(.a(s_117), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1370(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1371(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1372(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate2507(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2508(.a(gate144inter0), .b(s_280), .O(gate144inter1));
  and2  gate2509(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2510(.a(s_280), .O(gate144inter3));
  inv1  gate2511(.a(s_281), .O(gate144inter4));
  nand2 gate2512(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2513(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2514(.a(G468), .O(gate144inter7));
  inv1  gate2515(.a(G471), .O(gate144inter8));
  nand2 gate2516(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2517(.a(s_281), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2518(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2519(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2520(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate869(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate870(.a(gate148inter0), .b(s_46), .O(gate148inter1));
  and2  gate871(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate872(.a(s_46), .O(gate148inter3));
  inv1  gate873(.a(s_47), .O(gate148inter4));
  nand2 gate874(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate875(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate876(.a(G492), .O(gate148inter7));
  inv1  gate877(.a(G495), .O(gate148inter8));
  nand2 gate878(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate879(.a(s_47), .b(gate148inter3), .O(gate148inter10));
  nor2  gate880(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate881(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate882(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate589(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate590(.a(gate150inter0), .b(s_6), .O(gate150inter1));
  and2  gate591(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate592(.a(s_6), .O(gate150inter3));
  inv1  gate593(.a(s_7), .O(gate150inter4));
  nand2 gate594(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate595(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate596(.a(G504), .O(gate150inter7));
  inv1  gate597(.a(G507), .O(gate150inter8));
  nand2 gate598(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate599(.a(s_7), .b(gate150inter3), .O(gate150inter10));
  nor2  gate600(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate601(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate602(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1667(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1668(.a(gate154inter0), .b(s_160), .O(gate154inter1));
  and2  gate1669(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1670(.a(s_160), .O(gate154inter3));
  inv1  gate1671(.a(s_161), .O(gate154inter4));
  nand2 gate1672(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1673(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1674(.a(G429), .O(gate154inter7));
  inv1  gate1675(.a(G522), .O(gate154inter8));
  nand2 gate1676(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1677(.a(s_161), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1678(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1679(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1680(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2773(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2774(.a(gate160inter0), .b(s_318), .O(gate160inter1));
  and2  gate2775(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2776(.a(s_318), .O(gate160inter3));
  inv1  gate2777(.a(s_319), .O(gate160inter4));
  nand2 gate2778(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2779(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2780(.a(G447), .O(gate160inter7));
  inv1  gate2781(.a(G531), .O(gate160inter8));
  nand2 gate2782(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2783(.a(s_319), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2784(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2785(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2786(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1513(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1514(.a(gate165inter0), .b(s_138), .O(gate165inter1));
  and2  gate1515(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1516(.a(s_138), .O(gate165inter3));
  inv1  gate1517(.a(s_139), .O(gate165inter4));
  nand2 gate1518(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1519(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1520(.a(G462), .O(gate165inter7));
  inv1  gate1521(.a(G540), .O(gate165inter8));
  nand2 gate1522(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1523(.a(s_139), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1524(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1525(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1526(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate2549(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2550(.a(gate166inter0), .b(s_286), .O(gate166inter1));
  and2  gate2551(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2552(.a(s_286), .O(gate166inter3));
  inv1  gate2553(.a(s_287), .O(gate166inter4));
  nand2 gate2554(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2555(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2556(.a(G465), .O(gate166inter7));
  inv1  gate2557(.a(G540), .O(gate166inter8));
  nand2 gate2558(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2559(.a(s_287), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2560(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2561(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2562(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2241(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2242(.a(gate167inter0), .b(s_242), .O(gate167inter1));
  and2  gate2243(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2244(.a(s_242), .O(gate167inter3));
  inv1  gate2245(.a(s_243), .O(gate167inter4));
  nand2 gate2246(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2247(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2248(.a(G468), .O(gate167inter7));
  inv1  gate2249(.a(G543), .O(gate167inter8));
  nand2 gate2250(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2251(.a(s_243), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2252(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2253(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2254(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1093(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1094(.a(gate173inter0), .b(s_78), .O(gate173inter1));
  and2  gate1095(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1096(.a(s_78), .O(gate173inter3));
  inv1  gate1097(.a(s_79), .O(gate173inter4));
  nand2 gate1098(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1099(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1100(.a(G486), .O(gate173inter7));
  inv1  gate1101(.a(G552), .O(gate173inter8));
  nand2 gate1102(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1103(.a(s_79), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1104(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1105(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1106(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1457(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1458(.a(gate175inter0), .b(s_130), .O(gate175inter1));
  and2  gate1459(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1460(.a(s_130), .O(gate175inter3));
  inv1  gate1461(.a(s_131), .O(gate175inter4));
  nand2 gate1462(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1463(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1464(.a(G492), .O(gate175inter7));
  inv1  gate1465(.a(G555), .O(gate175inter8));
  nand2 gate1466(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1467(.a(s_131), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1468(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1469(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1470(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate2577(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2578(.a(gate176inter0), .b(s_290), .O(gate176inter1));
  and2  gate2579(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2580(.a(s_290), .O(gate176inter3));
  inv1  gate2581(.a(s_291), .O(gate176inter4));
  nand2 gate2582(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2583(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2584(.a(G495), .O(gate176inter7));
  inv1  gate2585(.a(G555), .O(gate176inter8));
  nand2 gate2586(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2587(.a(s_291), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2588(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2589(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2590(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate2843(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2844(.a(gate177inter0), .b(s_328), .O(gate177inter1));
  and2  gate2845(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2846(.a(s_328), .O(gate177inter3));
  inv1  gate2847(.a(s_329), .O(gate177inter4));
  nand2 gate2848(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2849(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2850(.a(G498), .O(gate177inter7));
  inv1  gate2851(.a(G558), .O(gate177inter8));
  nand2 gate2852(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2853(.a(s_329), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2854(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2855(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2856(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2647(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2648(.a(gate179inter0), .b(s_300), .O(gate179inter1));
  and2  gate2649(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2650(.a(s_300), .O(gate179inter3));
  inv1  gate2651(.a(s_301), .O(gate179inter4));
  nand2 gate2652(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2653(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2654(.a(G504), .O(gate179inter7));
  inv1  gate2655(.a(G561), .O(gate179inter8));
  nand2 gate2656(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2657(.a(s_301), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2658(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2659(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2660(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1009(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1010(.a(gate181inter0), .b(s_66), .O(gate181inter1));
  and2  gate1011(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1012(.a(s_66), .O(gate181inter3));
  inv1  gate1013(.a(s_67), .O(gate181inter4));
  nand2 gate1014(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1015(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1016(.a(G510), .O(gate181inter7));
  inv1  gate1017(.a(G564), .O(gate181inter8));
  nand2 gate1018(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1019(.a(s_67), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1020(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1021(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1022(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1247(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1248(.a(gate186inter0), .b(s_100), .O(gate186inter1));
  and2  gate1249(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1250(.a(s_100), .O(gate186inter3));
  inv1  gate1251(.a(s_101), .O(gate186inter4));
  nand2 gate1252(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1253(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1254(.a(G572), .O(gate186inter7));
  inv1  gate1255(.a(G573), .O(gate186inter8));
  nand2 gate1256(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1257(.a(s_101), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1258(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1259(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1260(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate757(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate758(.a(gate188inter0), .b(s_30), .O(gate188inter1));
  and2  gate759(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate760(.a(s_30), .O(gate188inter3));
  inv1  gate761(.a(s_31), .O(gate188inter4));
  nand2 gate762(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate763(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate764(.a(G576), .O(gate188inter7));
  inv1  gate765(.a(G577), .O(gate188inter8));
  nand2 gate766(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate767(.a(s_31), .b(gate188inter3), .O(gate188inter10));
  nor2  gate768(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate769(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate770(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1611(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1612(.a(gate189inter0), .b(s_152), .O(gate189inter1));
  and2  gate1613(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1614(.a(s_152), .O(gate189inter3));
  inv1  gate1615(.a(s_153), .O(gate189inter4));
  nand2 gate1616(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1617(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1618(.a(G578), .O(gate189inter7));
  inv1  gate1619(.a(G579), .O(gate189inter8));
  nand2 gate1620(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1621(.a(s_153), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1622(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1623(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1624(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate701(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate702(.a(gate190inter0), .b(s_22), .O(gate190inter1));
  and2  gate703(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate704(.a(s_22), .O(gate190inter3));
  inv1  gate705(.a(s_23), .O(gate190inter4));
  nand2 gate706(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate707(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate708(.a(G580), .O(gate190inter7));
  inv1  gate709(.a(G581), .O(gate190inter8));
  nand2 gate710(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate711(.a(s_23), .b(gate190inter3), .O(gate190inter10));
  nor2  gate712(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate713(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate714(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2045(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2046(.a(gate192inter0), .b(s_214), .O(gate192inter1));
  and2  gate2047(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2048(.a(s_214), .O(gate192inter3));
  inv1  gate2049(.a(s_215), .O(gate192inter4));
  nand2 gate2050(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2051(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2052(.a(G584), .O(gate192inter7));
  inv1  gate2053(.a(G585), .O(gate192inter8));
  nand2 gate2054(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2055(.a(s_215), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2056(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2057(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2058(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate2535(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2536(.a(gate199inter0), .b(s_284), .O(gate199inter1));
  and2  gate2537(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2538(.a(s_284), .O(gate199inter3));
  inv1  gate2539(.a(s_285), .O(gate199inter4));
  nand2 gate2540(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2541(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2542(.a(G598), .O(gate199inter7));
  inv1  gate2543(.a(G599), .O(gate199inter8));
  nand2 gate2544(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2545(.a(s_285), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2546(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2547(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2548(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate771(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate772(.a(gate200inter0), .b(s_32), .O(gate200inter1));
  and2  gate773(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate774(.a(s_32), .O(gate200inter3));
  inv1  gate775(.a(s_33), .O(gate200inter4));
  nand2 gate776(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate777(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate778(.a(G600), .O(gate200inter7));
  inv1  gate779(.a(G601), .O(gate200inter8));
  nand2 gate780(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate781(.a(s_33), .b(gate200inter3), .O(gate200inter10));
  nor2  gate782(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate783(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate784(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1737(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1738(.a(gate201inter0), .b(s_170), .O(gate201inter1));
  and2  gate1739(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1740(.a(s_170), .O(gate201inter3));
  inv1  gate1741(.a(s_171), .O(gate201inter4));
  nand2 gate1742(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1743(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1744(.a(G602), .O(gate201inter7));
  inv1  gate1745(.a(G607), .O(gate201inter8));
  nand2 gate1746(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1747(.a(s_171), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1748(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1749(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1750(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate855(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate856(.a(gate203inter0), .b(s_44), .O(gate203inter1));
  and2  gate857(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate858(.a(s_44), .O(gate203inter3));
  inv1  gate859(.a(s_45), .O(gate203inter4));
  nand2 gate860(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate861(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate862(.a(G602), .O(gate203inter7));
  inv1  gate863(.a(G612), .O(gate203inter8));
  nand2 gate864(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate865(.a(s_45), .b(gate203inter3), .O(gate203inter10));
  nor2  gate866(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate867(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate868(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2171(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2172(.a(gate208inter0), .b(s_232), .O(gate208inter1));
  and2  gate2173(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2174(.a(s_232), .O(gate208inter3));
  inv1  gate2175(.a(s_233), .O(gate208inter4));
  nand2 gate2176(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2177(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2178(.a(G627), .O(gate208inter7));
  inv1  gate2179(.a(G637), .O(gate208inter8));
  nand2 gate2180(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2181(.a(s_233), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2182(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2183(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2184(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1905(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1906(.a(gate213inter0), .b(s_194), .O(gate213inter1));
  and2  gate1907(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1908(.a(s_194), .O(gate213inter3));
  inv1  gate1909(.a(s_195), .O(gate213inter4));
  nand2 gate1910(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1911(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1912(.a(G602), .O(gate213inter7));
  inv1  gate1913(.a(G672), .O(gate213inter8));
  nand2 gate1914(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1915(.a(s_195), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1916(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1917(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1918(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2451(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2452(.a(gate214inter0), .b(s_272), .O(gate214inter1));
  and2  gate2453(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2454(.a(s_272), .O(gate214inter3));
  inv1  gate2455(.a(s_273), .O(gate214inter4));
  nand2 gate2456(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2457(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2458(.a(G612), .O(gate214inter7));
  inv1  gate2459(.a(G672), .O(gate214inter8));
  nand2 gate2460(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2461(.a(s_273), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2462(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2463(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2464(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2031(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2032(.a(gate215inter0), .b(s_212), .O(gate215inter1));
  and2  gate2033(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2034(.a(s_212), .O(gate215inter3));
  inv1  gate2035(.a(s_213), .O(gate215inter4));
  nand2 gate2036(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2037(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2038(.a(G607), .O(gate215inter7));
  inv1  gate2039(.a(G675), .O(gate215inter8));
  nand2 gate2040(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2041(.a(s_213), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2042(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2043(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2044(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2017(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2018(.a(gate220inter0), .b(s_210), .O(gate220inter1));
  and2  gate2019(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2020(.a(s_210), .O(gate220inter3));
  inv1  gate2021(.a(s_211), .O(gate220inter4));
  nand2 gate2022(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2023(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2024(.a(G637), .O(gate220inter7));
  inv1  gate2025(.a(G681), .O(gate220inter8));
  nand2 gate2026(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2027(.a(s_211), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2028(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2029(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2030(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1373(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1374(.a(gate221inter0), .b(s_118), .O(gate221inter1));
  and2  gate1375(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1376(.a(s_118), .O(gate221inter3));
  inv1  gate1377(.a(s_119), .O(gate221inter4));
  nand2 gate1378(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1379(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1380(.a(G622), .O(gate221inter7));
  inv1  gate1381(.a(G684), .O(gate221inter8));
  nand2 gate1382(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1383(.a(s_119), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1384(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1385(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1386(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2899(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2900(.a(gate223inter0), .b(s_336), .O(gate223inter1));
  and2  gate2901(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2902(.a(s_336), .O(gate223inter3));
  inv1  gate2903(.a(s_337), .O(gate223inter4));
  nand2 gate2904(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2905(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2906(.a(G627), .O(gate223inter7));
  inv1  gate2907(.a(G687), .O(gate223inter8));
  nand2 gate2908(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2909(.a(s_337), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2910(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2911(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2912(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate953(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate954(.a(gate225inter0), .b(s_58), .O(gate225inter1));
  and2  gate955(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate956(.a(s_58), .O(gate225inter3));
  inv1  gate957(.a(s_59), .O(gate225inter4));
  nand2 gate958(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate959(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate960(.a(G690), .O(gate225inter7));
  inv1  gate961(.a(G691), .O(gate225inter8));
  nand2 gate962(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate963(.a(s_59), .b(gate225inter3), .O(gate225inter10));
  nor2  gate964(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate965(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate966(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2227(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2228(.a(gate227inter0), .b(s_240), .O(gate227inter1));
  and2  gate2229(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2230(.a(s_240), .O(gate227inter3));
  inv1  gate2231(.a(s_241), .O(gate227inter4));
  nand2 gate2232(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2233(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2234(.a(G694), .O(gate227inter7));
  inv1  gate2235(.a(G695), .O(gate227inter8));
  nand2 gate2236(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2237(.a(s_241), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2238(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2239(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2240(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1807(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1808(.a(gate228inter0), .b(s_180), .O(gate228inter1));
  and2  gate1809(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1810(.a(s_180), .O(gate228inter3));
  inv1  gate1811(.a(s_181), .O(gate228inter4));
  nand2 gate1812(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1813(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1814(.a(G696), .O(gate228inter7));
  inv1  gate1815(.a(G697), .O(gate228inter8));
  nand2 gate1816(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1817(.a(s_181), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1818(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1819(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1820(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1261(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1262(.a(gate229inter0), .b(s_102), .O(gate229inter1));
  and2  gate1263(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1264(.a(s_102), .O(gate229inter3));
  inv1  gate1265(.a(s_103), .O(gate229inter4));
  nand2 gate1266(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1267(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1268(.a(G698), .O(gate229inter7));
  inv1  gate1269(.a(G699), .O(gate229inter8));
  nand2 gate1270(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1271(.a(s_103), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1272(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1273(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1274(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1023(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1024(.a(gate230inter0), .b(s_68), .O(gate230inter1));
  and2  gate1025(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1026(.a(s_68), .O(gate230inter3));
  inv1  gate1027(.a(s_69), .O(gate230inter4));
  nand2 gate1028(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1029(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1030(.a(G700), .O(gate230inter7));
  inv1  gate1031(.a(G701), .O(gate230inter8));
  nand2 gate1032(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1033(.a(s_69), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1034(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1035(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1036(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1933(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1934(.a(gate231inter0), .b(s_198), .O(gate231inter1));
  and2  gate1935(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1936(.a(s_198), .O(gate231inter3));
  inv1  gate1937(.a(s_199), .O(gate231inter4));
  nand2 gate1938(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1939(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1940(.a(G702), .O(gate231inter7));
  inv1  gate1941(.a(G703), .O(gate231inter8));
  nand2 gate1942(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1943(.a(s_199), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1944(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1945(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1946(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2059(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2060(.a(gate234inter0), .b(s_216), .O(gate234inter1));
  and2  gate2061(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2062(.a(s_216), .O(gate234inter3));
  inv1  gate2063(.a(s_217), .O(gate234inter4));
  nand2 gate2064(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2065(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2066(.a(G245), .O(gate234inter7));
  inv1  gate2067(.a(G721), .O(gate234inter8));
  nand2 gate2068(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2069(.a(s_217), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2070(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2071(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2072(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1849(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1850(.a(gate235inter0), .b(s_186), .O(gate235inter1));
  and2  gate1851(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1852(.a(s_186), .O(gate235inter3));
  inv1  gate1853(.a(s_187), .O(gate235inter4));
  nand2 gate1854(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1855(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1856(.a(G248), .O(gate235inter7));
  inv1  gate1857(.a(G724), .O(gate235inter8));
  nand2 gate1858(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1859(.a(s_187), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1860(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1861(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1862(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate575(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate576(.a(gate237inter0), .b(s_4), .O(gate237inter1));
  and2  gate577(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate578(.a(s_4), .O(gate237inter3));
  inv1  gate579(.a(s_5), .O(gate237inter4));
  nand2 gate580(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate581(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate582(.a(G254), .O(gate237inter7));
  inv1  gate583(.a(G706), .O(gate237inter8));
  nand2 gate584(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate585(.a(s_5), .b(gate237inter3), .O(gate237inter10));
  nor2  gate586(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate587(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate588(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate547(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate548(.a(gate238inter0), .b(s_0), .O(gate238inter1));
  and2  gate549(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate550(.a(s_0), .O(gate238inter3));
  inv1  gate551(.a(s_1), .O(gate238inter4));
  nand2 gate552(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate553(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate554(.a(G257), .O(gate238inter7));
  inv1  gate555(.a(G709), .O(gate238inter8));
  nand2 gate556(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate557(.a(s_1), .b(gate238inter3), .O(gate238inter10));
  nor2  gate558(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate559(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate560(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate561(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate562(.a(gate239inter0), .b(s_2), .O(gate239inter1));
  and2  gate563(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate564(.a(s_2), .O(gate239inter3));
  inv1  gate565(.a(s_3), .O(gate239inter4));
  nand2 gate566(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate567(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate568(.a(G260), .O(gate239inter7));
  inv1  gate569(.a(G712), .O(gate239inter8));
  nand2 gate570(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate571(.a(s_3), .b(gate239inter3), .O(gate239inter10));
  nor2  gate572(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate573(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate574(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1877(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1878(.a(gate241inter0), .b(s_190), .O(gate241inter1));
  and2  gate1879(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1880(.a(s_190), .O(gate241inter3));
  inv1  gate1881(.a(s_191), .O(gate241inter4));
  nand2 gate1882(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1883(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1884(.a(G242), .O(gate241inter7));
  inv1  gate1885(.a(G730), .O(gate241inter8));
  nand2 gate1886(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1887(.a(s_191), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1888(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1889(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1890(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2787(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2788(.a(gate243inter0), .b(s_320), .O(gate243inter1));
  and2  gate2789(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2790(.a(s_320), .O(gate243inter3));
  inv1  gate2791(.a(s_321), .O(gate243inter4));
  nand2 gate2792(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2793(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2794(.a(G245), .O(gate243inter7));
  inv1  gate2795(.a(G733), .O(gate243inter8));
  nand2 gate2796(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2797(.a(s_321), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2798(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2799(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2800(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1723(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1724(.a(gate245inter0), .b(s_168), .O(gate245inter1));
  and2  gate1725(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1726(.a(s_168), .O(gate245inter3));
  inv1  gate1727(.a(s_169), .O(gate245inter4));
  nand2 gate1728(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1729(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1730(.a(G248), .O(gate245inter7));
  inv1  gate1731(.a(G736), .O(gate245inter8));
  nand2 gate1732(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1733(.a(s_169), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1734(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1735(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1736(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1429(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1430(.a(gate249inter0), .b(s_126), .O(gate249inter1));
  and2  gate1431(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1432(.a(s_126), .O(gate249inter3));
  inv1  gate1433(.a(s_127), .O(gate249inter4));
  nand2 gate1434(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1435(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1436(.a(G254), .O(gate249inter7));
  inv1  gate1437(.a(G742), .O(gate249inter8));
  nand2 gate1438(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1439(.a(s_127), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1440(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1441(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1442(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate813(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate814(.a(gate252inter0), .b(s_38), .O(gate252inter1));
  and2  gate815(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate816(.a(s_38), .O(gate252inter3));
  inv1  gate817(.a(s_39), .O(gate252inter4));
  nand2 gate818(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate819(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate820(.a(G709), .O(gate252inter7));
  inv1  gate821(.a(G745), .O(gate252inter8));
  nand2 gate822(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate823(.a(s_39), .b(gate252inter3), .O(gate252inter10));
  nor2  gate824(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate825(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate826(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1387(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1388(.a(gate256inter0), .b(s_120), .O(gate256inter1));
  and2  gate1389(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1390(.a(s_120), .O(gate256inter3));
  inv1  gate1391(.a(s_121), .O(gate256inter4));
  nand2 gate1392(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1393(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1394(.a(G715), .O(gate256inter7));
  inv1  gate1395(.a(G751), .O(gate256inter8));
  nand2 gate1396(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1397(.a(s_121), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1398(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1399(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1400(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate631(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate632(.a(gate259inter0), .b(s_12), .O(gate259inter1));
  and2  gate633(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate634(.a(s_12), .O(gate259inter3));
  inv1  gate635(.a(s_13), .O(gate259inter4));
  nand2 gate636(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate637(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate638(.a(G758), .O(gate259inter7));
  inv1  gate639(.a(G759), .O(gate259inter8));
  nand2 gate640(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate641(.a(s_13), .b(gate259inter3), .O(gate259inter10));
  nor2  gate642(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate643(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate644(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate2143(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2144(.a(gate260inter0), .b(s_228), .O(gate260inter1));
  and2  gate2145(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2146(.a(s_228), .O(gate260inter3));
  inv1  gate2147(.a(s_229), .O(gate260inter4));
  nand2 gate2148(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2149(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2150(.a(G760), .O(gate260inter7));
  inv1  gate2151(.a(G761), .O(gate260inter8));
  nand2 gate2152(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2153(.a(s_229), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2154(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2155(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2156(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate603(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate604(.a(gate264inter0), .b(s_8), .O(gate264inter1));
  and2  gate605(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate606(.a(s_8), .O(gate264inter3));
  inv1  gate607(.a(s_9), .O(gate264inter4));
  nand2 gate608(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate609(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate610(.a(G768), .O(gate264inter7));
  inv1  gate611(.a(G769), .O(gate264inter8));
  nand2 gate612(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate613(.a(s_9), .b(gate264inter3), .O(gate264inter10));
  nor2  gate614(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate615(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate616(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate729(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate730(.a(gate268inter0), .b(s_26), .O(gate268inter1));
  and2  gate731(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate732(.a(s_26), .O(gate268inter3));
  inv1  gate733(.a(s_27), .O(gate268inter4));
  nand2 gate734(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate735(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate736(.a(G651), .O(gate268inter7));
  inv1  gate737(.a(G779), .O(gate268inter8));
  nand2 gate738(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate739(.a(s_27), .b(gate268inter3), .O(gate268inter10));
  nor2  gate740(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate741(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate742(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2633(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2634(.a(gate269inter0), .b(s_298), .O(gate269inter1));
  and2  gate2635(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2636(.a(s_298), .O(gate269inter3));
  inv1  gate2637(.a(s_299), .O(gate269inter4));
  nand2 gate2638(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2639(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2640(.a(G654), .O(gate269inter7));
  inv1  gate2641(.a(G782), .O(gate269inter8));
  nand2 gate2642(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2643(.a(s_299), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2644(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2645(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2646(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1709(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1710(.a(gate272inter0), .b(s_166), .O(gate272inter1));
  and2  gate1711(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1712(.a(s_166), .O(gate272inter3));
  inv1  gate1713(.a(s_167), .O(gate272inter4));
  nand2 gate1714(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1715(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1716(.a(G663), .O(gate272inter7));
  inv1  gate1717(.a(G791), .O(gate272inter8));
  nand2 gate1718(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1719(.a(s_167), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1720(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1721(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1722(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1317(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1318(.a(gate273inter0), .b(s_110), .O(gate273inter1));
  and2  gate1319(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1320(.a(s_110), .O(gate273inter3));
  inv1  gate1321(.a(s_111), .O(gate273inter4));
  nand2 gate1322(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1323(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1324(.a(G642), .O(gate273inter7));
  inv1  gate1325(.a(G794), .O(gate273inter8));
  nand2 gate1326(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1327(.a(s_111), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1328(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1329(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1330(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2339(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2340(.a(gate276inter0), .b(s_256), .O(gate276inter1));
  and2  gate2341(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2342(.a(s_256), .O(gate276inter3));
  inv1  gate2343(.a(s_257), .O(gate276inter4));
  nand2 gate2344(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2345(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2346(.a(G773), .O(gate276inter7));
  inv1  gate2347(.a(G797), .O(gate276inter8));
  nand2 gate2348(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2349(.a(s_257), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2350(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2351(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2352(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1499(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1500(.a(gate281inter0), .b(s_136), .O(gate281inter1));
  and2  gate1501(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1502(.a(s_136), .O(gate281inter3));
  inv1  gate1503(.a(s_137), .O(gate281inter4));
  nand2 gate1504(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1505(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1506(.a(G654), .O(gate281inter7));
  inv1  gate1507(.a(G806), .O(gate281inter8));
  nand2 gate1508(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1509(.a(s_137), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1510(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1511(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1512(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate967(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate968(.a(gate293inter0), .b(s_60), .O(gate293inter1));
  and2  gate969(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate970(.a(s_60), .O(gate293inter3));
  inv1  gate971(.a(s_61), .O(gate293inter4));
  nand2 gate972(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate973(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate974(.a(G828), .O(gate293inter7));
  inv1  gate975(.a(G829), .O(gate293inter8));
  nand2 gate976(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate977(.a(s_61), .b(gate293inter3), .O(gate293inter10));
  nor2  gate978(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate979(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate980(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate883(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate884(.a(gate294inter0), .b(s_48), .O(gate294inter1));
  and2  gate885(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate886(.a(s_48), .O(gate294inter3));
  inv1  gate887(.a(s_49), .O(gate294inter4));
  nand2 gate888(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate889(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate890(.a(G832), .O(gate294inter7));
  inv1  gate891(.a(G833), .O(gate294inter8));
  nand2 gate892(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate893(.a(s_49), .b(gate294inter3), .O(gate294inter10));
  nor2  gate894(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate895(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate896(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2717(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2718(.a(gate295inter0), .b(s_310), .O(gate295inter1));
  and2  gate2719(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2720(.a(s_310), .O(gate295inter3));
  inv1  gate2721(.a(s_311), .O(gate295inter4));
  nand2 gate2722(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2723(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2724(.a(G830), .O(gate295inter7));
  inv1  gate2725(.a(G831), .O(gate295inter8));
  nand2 gate2726(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2727(.a(s_311), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2728(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2729(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2730(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1121(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1122(.a(gate390inter0), .b(s_82), .O(gate390inter1));
  and2  gate1123(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1124(.a(s_82), .O(gate390inter3));
  inv1  gate1125(.a(s_83), .O(gate390inter4));
  nand2 gate1126(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1127(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1128(.a(G4), .O(gate390inter7));
  inv1  gate1129(.a(G1045), .O(gate390inter8));
  nand2 gate1130(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1131(.a(s_83), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1132(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1133(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1134(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate785(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate786(.a(gate392inter0), .b(s_34), .O(gate392inter1));
  and2  gate787(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate788(.a(s_34), .O(gate392inter3));
  inv1  gate789(.a(s_35), .O(gate392inter4));
  nand2 gate790(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate791(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate792(.a(G6), .O(gate392inter7));
  inv1  gate793(.a(G1051), .O(gate392inter8));
  nand2 gate794(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate795(.a(s_35), .b(gate392inter3), .O(gate392inter10));
  nor2  gate796(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate797(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate798(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate2605(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2606(.a(gate393inter0), .b(s_294), .O(gate393inter1));
  and2  gate2607(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2608(.a(s_294), .O(gate393inter3));
  inv1  gate2609(.a(s_295), .O(gate393inter4));
  nand2 gate2610(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2611(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2612(.a(G7), .O(gate393inter7));
  inv1  gate2613(.a(G1054), .O(gate393inter8));
  nand2 gate2614(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2615(.a(s_295), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2616(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2617(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2618(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate827(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate828(.a(gate399inter0), .b(s_40), .O(gate399inter1));
  and2  gate829(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate830(.a(s_40), .O(gate399inter3));
  inv1  gate831(.a(s_41), .O(gate399inter4));
  nand2 gate832(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate833(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate834(.a(G13), .O(gate399inter7));
  inv1  gate835(.a(G1072), .O(gate399inter8));
  nand2 gate836(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate837(.a(s_41), .b(gate399inter3), .O(gate399inter10));
  nor2  gate838(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate839(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate840(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1205(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1206(.a(gate400inter0), .b(s_94), .O(gate400inter1));
  and2  gate1207(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1208(.a(s_94), .O(gate400inter3));
  inv1  gate1209(.a(s_95), .O(gate400inter4));
  nand2 gate1210(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1211(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1212(.a(G14), .O(gate400inter7));
  inv1  gate1213(.a(G1075), .O(gate400inter8));
  nand2 gate1214(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1215(.a(s_95), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1216(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1217(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1218(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1541(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1542(.a(gate401inter0), .b(s_142), .O(gate401inter1));
  and2  gate1543(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1544(.a(s_142), .O(gate401inter3));
  inv1  gate1545(.a(s_143), .O(gate401inter4));
  nand2 gate1546(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1547(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1548(.a(G15), .O(gate401inter7));
  inv1  gate1549(.a(G1078), .O(gate401inter8));
  nand2 gate1550(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1551(.a(s_143), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1552(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1553(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1554(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate981(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate982(.a(gate404inter0), .b(s_62), .O(gate404inter1));
  and2  gate983(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate984(.a(s_62), .O(gate404inter3));
  inv1  gate985(.a(s_63), .O(gate404inter4));
  nand2 gate986(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate987(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate988(.a(G18), .O(gate404inter7));
  inv1  gate989(.a(G1087), .O(gate404inter8));
  nand2 gate990(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate991(.a(s_63), .b(gate404inter3), .O(gate404inter10));
  nor2  gate992(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate993(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate994(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate2423(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2424(.a(gate405inter0), .b(s_268), .O(gate405inter1));
  and2  gate2425(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2426(.a(s_268), .O(gate405inter3));
  inv1  gate2427(.a(s_269), .O(gate405inter4));
  nand2 gate2428(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2429(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2430(.a(G19), .O(gate405inter7));
  inv1  gate2431(.a(G1090), .O(gate405inter8));
  nand2 gate2432(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2433(.a(s_269), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2434(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2435(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2436(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2857(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2858(.a(gate406inter0), .b(s_330), .O(gate406inter1));
  and2  gate2859(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2860(.a(s_330), .O(gate406inter3));
  inv1  gate2861(.a(s_331), .O(gate406inter4));
  nand2 gate2862(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2863(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2864(.a(G20), .O(gate406inter7));
  inv1  gate2865(.a(G1093), .O(gate406inter8));
  nand2 gate2866(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2867(.a(s_331), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2868(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2869(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2870(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1415(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1416(.a(gate407inter0), .b(s_124), .O(gate407inter1));
  and2  gate1417(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1418(.a(s_124), .O(gate407inter3));
  inv1  gate1419(.a(s_125), .O(gate407inter4));
  nand2 gate1420(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1421(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1422(.a(G21), .O(gate407inter7));
  inv1  gate1423(.a(G1096), .O(gate407inter8));
  nand2 gate1424(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1425(.a(s_125), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1426(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1427(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1428(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate2087(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2088(.a(gate408inter0), .b(s_220), .O(gate408inter1));
  and2  gate2089(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2090(.a(s_220), .O(gate408inter3));
  inv1  gate2091(.a(s_221), .O(gate408inter4));
  nand2 gate2092(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2093(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2094(.a(G22), .O(gate408inter7));
  inv1  gate2095(.a(G1099), .O(gate408inter8));
  nand2 gate2096(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2097(.a(s_221), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2098(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2099(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2100(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1135(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1136(.a(gate411inter0), .b(s_84), .O(gate411inter1));
  and2  gate1137(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1138(.a(s_84), .O(gate411inter3));
  inv1  gate1139(.a(s_85), .O(gate411inter4));
  nand2 gate1140(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1141(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1142(.a(G25), .O(gate411inter7));
  inv1  gate1143(.a(G1108), .O(gate411inter8));
  nand2 gate1144(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1145(.a(s_85), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1146(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1147(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1148(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1751(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1752(.a(gate415inter0), .b(s_172), .O(gate415inter1));
  and2  gate1753(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1754(.a(s_172), .O(gate415inter3));
  inv1  gate1755(.a(s_173), .O(gate415inter4));
  nand2 gate1756(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1757(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1758(.a(G29), .O(gate415inter7));
  inv1  gate1759(.a(G1120), .O(gate415inter8));
  nand2 gate1760(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1761(.a(s_173), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1762(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1763(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1764(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2927(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2928(.a(gate417inter0), .b(s_340), .O(gate417inter1));
  and2  gate2929(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2930(.a(s_340), .O(gate417inter3));
  inv1  gate2931(.a(s_341), .O(gate417inter4));
  nand2 gate2932(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2933(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2934(.a(G31), .O(gate417inter7));
  inv1  gate2935(.a(G1126), .O(gate417inter8));
  nand2 gate2936(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2937(.a(s_341), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2938(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2939(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2940(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2661(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2662(.a(gate418inter0), .b(s_302), .O(gate418inter1));
  and2  gate2663(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2664(.a(s_302), .O(gate418inter3));
  inv1  gate2665(.a(s_303), .O(gate418inter4));
  nand2 gate2666(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2667(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2668(.a(G32), .O(gate418inter7));
  inv1  gate2669(.a(G1129), .O(gate418inter8));
  nand2 gate2670(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2671(.a(s_303), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2672(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2673(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2674(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1401(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1402(.a(gate422inter0), .b(s_122), .O(gate422inter1));
  and2  gate1403(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1404(.a(s_122), .O(gate422inter3));
  inv1  gate1405(.a(s_123), .O(gate422inter4));
  nand2 gate1406(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1407(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1408(.a(G1039), .O(gate422inter7));
  inv1  gate1409(.a(G1135), .O(gate422inter8));
  nand2 gate1410(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1411(.a(s_123), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1412(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1413(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1414(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate2115(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2116(.a(gate423inter0), .b(s_224), .O(gate423inter1));
  and2  gate2117(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2118(.a(s_224), .O(gate423inter3));
  inv1  gate2119(.a(s_225), .O(gate423inter4));
  nand2 gate2120(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2121(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2122(.a(G3), .O(gate423inter7));
  inv1  gate2123(.a(G1138), .O(gate423inter8));
  nand2 gate2124(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2125(.a(s_225), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2126(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2127(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2128(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2703(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2704(.a(gate424inter0), .b(s_308), .O(gate424inter1));
  and2  gate2705(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2706(.a(s_308), .O(gate424inter3));
  inv1  gate2707(.a(s_309), .O(gate424inter4));
  nand2 gate2708(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2709(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2710(.a(G1042), .O(gate424inter7));
  inv1  gate2711(.a(G1138), .O(gate424inter8));
  nand2 gate2712(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2713(.a(s_309), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2714(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2715(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2716(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate2213(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2214(.a(gate425inter0), .b(s_238), .O(gate425inter1));
  and2  gate2215(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2216(.a(s_238), .O(gate425inter3));
  inv1  gate2217(.a(s_239), .O(gate425inter4));
  nand2 gate2218(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2219(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2220(.a(G4), .O(gate425inter7));
  inv1  gate2221(.a(G1141), .O(gate425inter8));
  nand2 gate2222(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2223(.a(s_239), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2224(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2225(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2226(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate743(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate744(.a(gate426inter0), .b(s_28), .O(gate426inter1));
  and2  gate745(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate746(.a(s_28), .O(gate426inter3));
  inv1  gate747(.a(s_29), .O(gate426inter4));
  nand2 gate748(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate749(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate750(.a(G1045), .O(gate426inter7));
  inv1  gate751(.a(G1141), .O(gate426inter8));
  nand2 gate752(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate753(.a(s_29), .b(gate426inter3), .O(gate426inter10));
  nor2  gate754(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate755(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate756(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2297(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2298(.a(gate428inter0), .b(s_250), .O(gate428inter1));
  and2  gate2299(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2300(.a(s_250), .O(gate428inter3));
  inv1  gate2301(.a(s_251), .O(gate428inter4));
  nand2 gate2302(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2303(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2304(.a(G1048), .O(gate428inter7));
  inv1  gate2305(.a(G1144), .O(gate428inter8));
  nand2 gate2306(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2307(.a(s_251), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2308(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2309(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2310(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2885(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2886(.a(gate430inter0), .b(s_334), .O(gate430inter1));
  and2  gate2887(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2888(.a(s_334), .O(gate430inter3));
  inv1  gate2889(.a(s_335), .O(gate430inter4));
  nand2 gate2890(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2891(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2892(.a(G1051), .O(gate430inter7));
  inv1  gate2893(.a(G1147), .O(gate430inter8));
  nand2 gate2894(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2895(.a(s_335), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2896(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2897(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2898(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2185(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2186(.a(gate431inter0), .b(s_234), .O(gate431inter1));
  and2  gate2187(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2188(.a(s_234), .O(gate431inter3));
  inv1  gate2189(.a(s_235), .O(gate431inter4));
  nand2 gate2190(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2191(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2192(.a(G7), .O(gate431inter7));
  inv1  gate2193(.a(G1150), .O(gate431inter8));
  nand2 gate2194(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2195(.a(s_235), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2196(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2197(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2198(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate687(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate688(.a(gate432inter0), .b(s_20), .O(gate432inter1));
  and2  gate689(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate690(.a(s_20), .O(gate432inter3));
  inv1  gate691(.a(s_21), .O(gate432inter4));
  nand2 gate692(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate693(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate694(.a(G1054), .O(gate432inter7));
  inv1  gate695(.a(G1150), .O(gate432inter8));
  nand2 gate696(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate697(.a(s_21), .b(gate432inter3), .O(gate432inter10));
  nor2  gate698(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate699(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate700(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1345(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1346(.a(gate434inter0), .b(s_114), .O(gate434inter1));
  and2  gate1347(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1348(.a(s_114), .O(gate434inter3));
  inv1  gate1349(.a(s_115), .O(gate434inter4));
  nand2 gate1350(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1351(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1352(.a(G1057), .O(gate434inter7));
  inv1  gate1353(.a(G1153), .O(gate434inter8));
  nand2 gate1354(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1355(.a(s_115), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1356(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1357(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1358(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate2409(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2410(.a(gate436inter0), .b(s_266), .O(gate436inter1));
  and2  gate2411(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2412(.a(s_266), .O(gate436inter3));
  inv1  gate2413(.a(s_267), .O(gate436inter4));
  nand2 gate2414(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2415(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2416(.a(G1060), .O(gate436inter7));
  inv1  gate2417(.a(G1156), .O(gate436inter8));
  nand2 gate2418(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2419(.a(s_267), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2420(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2421(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2422(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate2479(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2480(.a(gate437inter0), .b(s_276), .O(gate437inter1));
  and2  gate2481(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2482(.a(s_276), .O(gate437inter3));
  inv1  gate2483(.a(s_277), .O(gate437inter4));
  nand2 gate2484(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2485(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2486(.a(G10), .O(gate437inter7));
  inv1  gate2487(.a(G1159), .O(gate437inter8));
  nand2 gate2488(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2489(.a(s_277), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2490(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2491(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2492(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1471(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1472(.a(gate439inter0), .b(s_132), .O(gate439inter1));
  and2  gate1473(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1474(.a(s_132), .O(gate439inter3));
  inv1  gate1475(.a(s_133), .O(gate439inter4));
  nand2 gate1476(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1477(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1478(.a(G11), .O(gate439inter7));
  inv1  gate1479(.a(G1162), .O(gate439inter8));
  nand2 gate1480(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1481(.a(s_133), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1482(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1483(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1484(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate2283(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2284(.a(gate440inter0), .b(s_248), .O(gate440inter1));
  and2  gate2285(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2286(.a(s_248), .O(gate440inter3));
  inv1  gate2287(.a(s_249), .O(gate440inter4));
  nand2 gate2288(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2289(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2290(.a(G1066), .O(gate440inter7));
  inv1  gate2291(.a(G1162), .O(gate440inter8));
  nand2 gate2292(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2293(.a(s_249), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2294(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2295(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2296(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1779(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1780(.a(gate441inter0), .b(s_176), .O(gate441inter1));
  and2  gate1781(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1782(.a(s_176), .O(gate441inter3));
  inv1  gate1783(.a(s_177), .O(gate441inter4));
  nand2 gate1784(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1785(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1786(.a(G12), .O(gate441inter7));
  inv1  gate1787(.a(G1165), .O(gate441inter8));
  nand2 gate1788(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1789(.a(s_177), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1790(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1791(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1792(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2815(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2816(.a(gate444inter0), .b(s_324), .O(gate444inter1));
  and2  gate2817(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2818(.a(s_324), .O(gate444inter3));
  inv1  gate2819(.a(s_325), .O(gate444inter4));
  nand2 gate2820(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2821(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2822(.a(G1072), .O(gate444inter7));
  inv1  gate2823(.a(G1168), .O(gate444inter8));
  nand2 gate2824(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2825(.a(s_325), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2826(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2827(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2828(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1485(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1486(.a(gate445inter0), .b(s_134), .O(gate445inter1));
  and2  gate1487(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1488(.a(s_134), .O(gate445inter3));
  inv1  gate1489(.a(s_135), .O(gate445inter4));
  nand2 gate1490(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1491(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1492(.a(G14), .O(gate445inter7));
  inv1  gate1493(.a(G1171), .O(gate445inter8));
  nand2 gate1494(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1495(.a(s_135), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1496(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1497(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1498(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1331(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1332(.a(gate448inter0), .b(s_112), .O(gate448inter1));
  and2  gate1333(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1334(.a(s_112), .O(gate448inter3));
  inv1  gate1335(.a(s_113), .O(gate448inter4));
  nand2 gate1336(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1337(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1338(.a(G1078), .O(gate448inter7));
  inv1  gate1339(.a(G1174), .O(gate448inter8));
  nand2 gate1340(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1341(.a(s_113), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1342(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1343(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1344(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1289(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1290(.a(gate449inter0), .b(s_106), .O(gate449inter1));
  and2  gate1291(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1292(.a(s_106), .O(gate449inter3));
  inv1  gate1293(.a(s_107), .O(gate449inter4));
  nand2 gate1294(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1295(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1296(.a(G16), .O(gate449inter7));
  inv1  gate1297(.a(G1177), .O(gate449inter8));
  nand2 gate1298(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1299(.a(s_107), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1300(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1301(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1302(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1625(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1626(.a(gate450inter0), .b(s_154), .O(gate450inter1));
  and2  gate1627(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1628(.a(s_154), .O(gate450inter3));
  inv1  gate1629(.a(s_155), .O(gate450inter4));
  nand2 gate1630(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1631(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1632(.a(G1081), .O(gate450inter7));
  inv1  gate1633(.a(G1177), .O(gate450inter8));
  nand2 gate1634(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1635(.a(s_155), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1636(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1637(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1638(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1443(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1444(.a(gate452inter0), .b(s_128), .O(gate452inter1));
  and2  gate1445(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1446(.a(s_128), .O(gate452inter3));
  inv1  gate1447(.a(s_129), .O(gate452inter4));
  nand2 gate1448(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1449(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1450(.a(G1084), .O(gate452inter7));
  inv1  gate1451(.a(G1180), .O(gate452inter8));
  nand2 gate1452(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1453(.a(s_129), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1454(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1455(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1456(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate2101(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2102(.a(gate453inter0), .b(s_222), .O(gate453inter1));
  and2  gate2103(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2104(.a(s_222), .O(gate453inter3));
  inv1  gate2105(.a(s_223), .O(gate453inter4));
  nand2 gate2106(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2107(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2108(.a(G18), .O(gate453inter7));
  inv1  gate2109(.a(G1183), .O(gate453inter8));
  nand2 gate2110(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2111(.a(s_223), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2112(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2113(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2114(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2829(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2830(.a(gate455inter0), .b(s_326), .O(gate455inter1));
  and2  gate2831(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2832(.a(s_326), .O(gate455inter3));
  inv1  gate2833(.a(s_327), .O(gate455inter4));
  nand2 gate2834(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2835(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2836(.a(G19), .O(gate455inter7));
  inv1  gate2837(.a(G1186), .O(gate455inter8));
  nand2 gate2838(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2839(.a(s_327), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2840(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2841(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2842(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate2437(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2438(.a(gate456inter0), .b(s_270), .O(gate456inter1));
  and2  gate2439(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2440(.a(s_270), .O(gate456inter3));
  inv1  gate2441(.a(s_271), .O(gate456inter4));
  nand2 gate2442(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2443(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2444(.a(G1090), .O(gate456inter7));
  inv1  gate2445(.a(G1186), .O(gate456inter8));
  nand2 gate2446(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2447(.a(s_271), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2448(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2449(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2450(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2129(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2130(.a(gate460inter0), .b(s_226), .O(gate460inter1));
  and2  gate2131(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2132(.a(s_226), .O(gate460inter3));
  inv1  gate2133(.a(s_227), .O(gate460inter4));
  nand2 gate2134(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2135(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2136(.a(G1096), .O(gate460inter7));
  inv1  gate2137(.a(G1192), .O(gate460inter8));
  nand2 gate2138(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2139(.a(s_227), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2140(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2141(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2142(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2521(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2522(.a(gate463inter0), .b(s_282), .O(gate463inter1));
  and2  gate2523(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2524(.a(s_282), .O(gate463inter3));
  inv1  gate2525(.a(s_283), .O(gate463inter4));
  nand2 gate2526(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2527(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2528(.a(G23), .O(gate463inter7));
  inv1  gate2529(.a(G1198), .O(gate463inter8));
  nand2 gate2530(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2531(.a(s_283), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2532(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2533(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2534(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate995(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate996(.a(gate464inter0), .b(s_64), .O(gate464inter1));
  and2  gate997(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate998(.a(s_64), .O(gate464inter3));
  inv1  gate999(.a(s_65), .O(gate464inter4));
  nand2 gate1000(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1001(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1002(.a(G1102), .O(gate464inter7));
  inv1  gate1003(.a(G1198), .O(gate464inter8));
  nand2 gate1004(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1005(.a(s_65), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1006(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1007(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1008(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1107(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1108(.a(gate469inter0), .b(s_80), .O(gate469inter1));
  and2  gate1109(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1110(.a(s_80), .O(gate469inter3));
  inv1  gate1111(.a(s_81), .O(gate469inter4));
  nand2 gate1112(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1113(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1114(.a(G26), .O(gate469inter7));
  inv1  gate1115(.a(G1207), .O(gate469inter8));
  nand2 gate1116(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1117(.a(s_81), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1118(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1119(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1120(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1975(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1976(.a(gate472inter0), .b(s_204), .O(gate472inter1));
  and2  gate1977(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1978(.a(s_204), .O(gate472inter3));
  inv1  gate1979(.a(s_205), .O(gate472inter4));
  nand2 gate1980(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1981(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1982(.a(G1114), .O(gate472inter7));
  inv1  gate1983(.a(G1210), .O(gate472inter8));
  nand2 gate1984(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1985(.a(s_205), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1986(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1987(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1988(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1555(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1556(.a(gate474inter0), .b(s_144), .O(gate474inter1));
  and2  gate1557(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1558(.a(s_144), .O(gate474inter3));
  inv1  gate1559(.a(s_145), .O(gate474inter4));
  nand2 gate1560(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1561(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1562(.a(G1117), .O(gate474inter7));
  inv1  gate1563(.a(G1213), .O(gate474inter8));
  nand2 gate1564(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1565(.a(s_145), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1566(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1567(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1568(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1947(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1948(.a(gate477inter0), .b(s_200), .O(gate477inter1));
  and2  gate1949(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1950(.a(s_200), .O(gate477inter3));
  inv1  gate1951(.a(s_201), .O(gate477inter4));
  nand2 gate1952(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1953(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1954(.a(G30), .O(gate477inter7));
  inv1  gate1955(.a(G1219), .O(gate477inter8));
  nand2 gate1956(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1957(.a(s_201), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1958(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1959(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1960(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1821(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1822(.a(gate478inter0), .b(s_182), .O(gate478inter1));
  and2  gate1823(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1824(.a(s_182), .O(gate478inter3));
  inv1  gate1825(.a(s_183), .O(gate478inter4));
  nand2 gate1826(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1827(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1828(.a(G1123), .O(gate478inter7));
  inv1  gate1829(.a(G1219), .O(gate478inter8));
  nand2 gate1830(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1831(.a(s_183), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1832(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1833(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1834(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1233(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1234(.a(gate479inter0), .b(s_98), .O(gate479inter1));
  and2  gate1235(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1236(.a(s_98), .O(gate479inter3));
  inv1  gate1237(.a(s_99), .O(gate479inter4));
  nand2 gate1238(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1239(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1240(.a(G31), .O(gate479inter7));
  inv1  gate1241(.a(G1222), .O(gate479inter8));
  nand2 gate1242(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1243(.a(s_99), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1244(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1245(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1246(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate2269(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2270(.a(gate487inter0), .b(s_246), .O(gate487inter1));
  and2  gate2271(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2272(.a(s_246), .O(gate487inter3));
  inv1  gate2273(.a(s_247), .O(gate487inter4));
  nand2 gate2274(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2275(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2276(.a(G1236), .O(gate487inter7));
  inv1  gate2277(.a(G1237), .O(gate487inter8));
  nand2 gate2278(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2279(.a(s_247), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2280(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2281(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2282(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1037(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1038(.a(gate488inter0), .b(s_70), .O(gate488inter1));
  and2  gate1039(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1040(.a(s_70), .O(gate488inter3));
  inv1  gate1041(.a(s_71), .O(gate488inter4));
  nand2 gate1042(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1043(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1044(.a(G1238), .O(gate488inter7));
  inv1  gate1045(.a(G1239), .O(gate488inter8));
  nand2 gate1046(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1047(.a(s_71), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1048(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1049(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1050(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2325(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2326(.a(gate490inter0), .b(s_254), .O(gate490inter1));
  and2  gate2327(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2328(.a(s_254), .O(gate490inter3));
  inv1  gate2329(.a(s_255), .O(gate490inter4));
  nand2 gate2330(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2331(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2332(.a(G1242), .O(gate490inter7));
  inv1  gate2333(.a(G1243), .O(gate490inter8));
  nand2 gate2334(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2335(.a(s_255), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2336(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2337(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2338(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2353(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2354(.a(gate493inter0), .b(s_258), .O(gate493inter1));
  and2  gate2355(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2356(.a(s_258), .O(gate493inter3));
  inv1  gate2357(.a(s_259), .O(gate493inter4));
  nand2 gate2358(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2359(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2360(.a(G1248), .O(gate493inter7));
  inv1  gate2361(.a(G1249), .O(gate493inter8));
  nand2 gate2362(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2363(.a(s_259), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2364(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2365(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2366(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate2367(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2368(.a(gate495inter0), .b(s_260), .O(gate495inter1));
  and2  gate2369(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2370(.a(s_260), .O(gate495inter3));
  inv1  gate2371(.a(s_261), .O(gate495inter4));
  nand2 gate2372(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2373(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2374(.a(G1252), .O(gate495inter7));
  inv1  gate2375(.a(G1253), .O(gate495inter8));
  nand2 gate2376(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2377(.a(s_261), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2378(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2379(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2380(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2745(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2746(.a(gate497inter0), .b(s_314), .O(gate497inter1));
  and2  gate2747(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2748(.a(s_314), .O(gate497inter3));
  inv1  gate2749(.a(s_315), .O(gate497inter4));
  nand2 gate2750(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2751(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2752(.a(G1256), .O(gate497inter7));
  inv1  gate2753(.a(G1257), .O(gate497inter8));
  nand2 gate2754(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2755(.a(s_315), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2756(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2757(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2758(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2689(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2690(.a(gate499inter0), .b(s_306), .O(gate499inter1));
  and2  gate2691(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2692(.a(s_306), .O(gate499inter3));
  inv1  gate2693(.a(s_307), .O(gate499inter4));
  nand2 gate2694(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2695(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2696(.a(G1260), .O(gate499inter7));
  inv1  gate2697(.a(G1261), .O(gate499inter8));
  nand2 gate2698(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2699(.a(s_307), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2700(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2701(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2702(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2381(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2382(.a(gate501inter0), .b(s_262), .O(gate501inter1));
  and2  gate2383(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2384(.a(s_262), .O(gate501inter3));
  inv1  gate2385(.a(s_263), .O(gate501inter4));
  nand2 gate2386(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2387(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2388(.a(G1264), .O(gate501inter7));
  inv1  gate2389(.a(G1265), .O(gate501inter8));
  nand2 gate2390(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2391(.a(s_263), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2392(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2393(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2394(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1793(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1794(.a(gate506inter0), .b(s_178), .O(gate506inter1));
  and2  gate1795(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1796(.a(s_178), .O(gate506inter3));
  inv1  gate1797(.a(s_179), .O(gate506inter4));
  nand2 gate1798(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1799(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1800(.a(G1274), .O(gate506inter7));
  inv1  gate1801(.a(G1275), .O(gate506inter8));
  nand2 gate1802(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1803(.a(s_179), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1804(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1805(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1806(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate841(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate842(.a(gate508inter0), .b(s_42), .O(gate508inter1));
  and2  gate843(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate844(.a(s_42), .O(gate508inter3));
  inv1  gate845(.a(s_43), .O(gate508inter4));
  nand2 gate846(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate847(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate848(.a(G1278), .O(gate508inter7));
  inv1  gate849(.a(G1279), .O(gate508inter8));
  nand2 gate850(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate851(.a(s_43), .b(gate508inter3), .O(gate508inter10));
  nor2  gate852(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate853(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate854(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate673(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate674(.a(gate509inter0), .b(s_18), .O(gate509inter1));
  and2  gate675(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate676(.a(s_18), .O(gate509inter3));
  inv1  gate677(.a(s_19), .O(gate509inter4));
  nand2 gate678(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate679(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate680(.a(G1280), .O(gate509inter7));
  inv1  gate681(.a(G1281), .O(gate509inter8));
  nand2 gate682(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate683(.a(s_19), .b(gate509inter3), .O(gate509inter10));
  nor2  gate684(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate685(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate686(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1065(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1066(.a(gate513inter0), .b(s_74), .O(gate513inter1));
  and2  gate1067(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1068(.a(s_74), .O(gate513inter3));
  inv1  gate1069(.a(s_75), .O(gate513inter4));
  nand2 gate1070(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1071(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1072(.a(G1288), .O(gate513inter7));
  inv1  gate1073(.a(G1289), .O(gate513inter8));
  nand2 gate1074(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1075(.a(s_75), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1076(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1077(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1078(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule