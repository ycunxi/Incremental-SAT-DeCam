module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );

  xor2  gate301(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate302(.a(gate2inter0), .b(s_14), .O(gate2inter1));
  and2  gate303(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate304(.a(s_14), .O(gate2inter3));
  inv1  gate305(.a(s_15), .O(gate2inter4));
  nand2 gate306(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate307(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate308(.a(N9), .O(gate2inter7));
  inv1  gate309(.a(N13), .O(gate2inter8));
  nand2 gate310(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate311(.a(s_15), .b(gate2inter3), .O(gate2inter10));
  nor2  gate312(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate313(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate314(.a(gate2inter12), .b(gate2inter1), .O(N251));
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate777(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate778(.a(gate4inter0), .b(s_82), .O(gate4inter1));
  and2  gate779(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate780(.a(s_82), .O(gate4inter3));
  inv1  gate781(.a(s_83), .O(gate4inter4));
  nand2 gate782(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate783(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate784(.a(N25), .O(gate4inter7));
  inv1  gate785(.a(N29), .O(gate4inter8));
  nand2 gate786(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate787(.a(s_83), .b(gate4inter3), .O(gate4inter10));
  nor2  gate788(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate789(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate790(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate721(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate722(.a(gate6inter0), .b(s_74), .O(gate6inter1));
  and2  gate723(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate724(.a(s_74), .O(gate6inter3));
  inv1  gate725(.a(s_75), .O(gate6inter4));
  nand2 gate726(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate727(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate728(.a(N41), .O(gate6inter7));
  inv1  gate729(.a(N45), .O(gate6inter8));
  nand2 gate730(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate731(.a(s_75), .b(gate6inter3), .O(gate6inter10));
  nor2  gate732(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate733(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate734(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate651(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate652(.a(gate8inter0), .b(s_64), .O(gate8inter1));
  and2  gate653(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate654(.a(s_64), .O(gate8inter3));
  inv1  gate655(.a(s_65), .O(gate8inter4));
  nand2 gate656(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate657(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate658(.a(N57), .O(gate8inter7));
  inv1  gate659(.a(N61), .O(gate8inter8));
  nand2 gate660(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate661(.a(s_65), .b(gate8inter3), .O(gate8inter10));
  nor2  gate662(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate663(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate664(.a(gate8inter12), .b(gate8inter1), .O(N257));
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );

  xor2  gate217(.a(N93), .b(N89), .O(gate12inter0));
  nand2 gate218(.a(gate12inter0), .b(s_2), .O(gate12inter1));
  and2  gate219(.a(N93), .b(N89), .O(gate12inter2));
  inv1  gate220(.a(s_2), .O(gate12inter3));
  inv1  gate221(.a(s_3), .O(gate12inter4));
  nand2 gate222(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate223(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate224(.a(N89), .O(gate12inter7));
  inv1  gate225(.a(N93), .O(gate12inter8));
  nand2 gate226(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate227(.a(s_3), .b(gate12inter3), .O(gate12inter10));
  nor2  gate228(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate229(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate230(.a(gate12inter12), .b(gate12inter1), .O(N261));

  xor2  gate833(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate834(.a(gate13inter0), .b(s_90), .O(gate13inter1));
  and2  gate835(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate836(.a(s_90), .O(gate13inter3));
  inv1  gate837(.a(s_91), .O(gate13inter4));
  nand2 gate838(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate839(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate840(.a(N97), .O(gate13inter7));
  inv1  gate841(.a(N101), .O(gate13inter8));
  nand2 gate842(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate843(.a(s_91), .b(gate13inter3), .O(gate13inter10));
  nor2  gate844(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate845(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate846(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate427(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate428(.a(gate25inter0), .b(s_32), .O(gate25inter1));
  and2  gate429(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate430(.a(s_32), .O(gate25inter3));
  inv1  gate431(.a(s_33), .O(gate25inter4));
  nand2 gate432(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate433(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate434(.a(N1), .O(gate25inter7));
  inv1  gate435(.a(N17), .O(gate25inter8));
  nand2 gate436(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate437(.a(s_33), .b(gate25inter3), .O(gate25inter10));
  nor2  gate438(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate439(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate440(.a(gate25inter12), .b(gate25inter1), .O(N274));

  xor2  gate371(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate372(.a(gate26inter0), .b(s_24), .O(gate26inter1));
  and2  gate373(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate374(.a(s_24), .O(gate26inter3));
  inv1  gate375(.a(s_25), .O(gate26inter4));
  nand2 gate376(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate377(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate378(.a(N33), .O(gate26inter7));
  inv1  gate379(.a(N49), .O(gate26inter8));
  nand2 gate380(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate381(.a(s_25), .b(gate26inter3), .O(gate26inter10));
  nor2  gate382(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate383(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate384(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );

  xor2  gate791(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate792(.a(gate28inter0), .b(s_84), .O(gate28inter1));
  and2  gate793(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate794(.a(s_84), .O(gate28inter3));
  inv1  gate795(.a(s_85), .O(gate28inter4));
  nand2 gate796(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate797(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate798(.a(N37), .O(gate28inter7));
  inv1  gate799(.a(N53), .O(gate28inter8));
  nand2 gate800(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate801(.a(s_85), .b(gate28inter3), .O(gate28inter10));
  nor2  gate802(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate803(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate804(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );

  xor2  gate273(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate274(.a(gate32inter0), .b(s_10), .O(gate32inter1));
  and2  gate275(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate276(.a(s_10), .O(gate32inter3));
  inv1  gate277(.a(s_11), .O(gate32inter4));
  nand2 gate278(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate279(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate280(.a(N45), .O(gate32inter7));
  inv1  gate281(.a(N61), .O(gate32inter8));
  nand2 gate282(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate283(.a(s_11), .b(gate32inter3), .O(gate32inter10));
  nor2  gate284(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate285(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate286(.a(gate32inter12), .b(gate32inter1), .O(N281));

  xor2  gate693(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate694(.a(gate33inter0), .b(s_70), .O(gate33inter1));
  and2  gate695(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate696(.a(s_70), .O(gate33inter3));
  inv1  gate697(.a(s_71), .O(gate33inter4));
  nand2 gate698(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate699(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate700(.a(N65), .O(gate33inter7));
  inv1  gate701(.a(N81), .O(gate33inter8));
  nand2 gate702(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate703(.a(s_71), .b(gate33inter3), .O(gate33inter10));
  nor2  gate704(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate705(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate706(.a(gate33inter12), .b(gate33inter1), .O(N282));
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );

  xor2  gate231(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate232(.a(gate36inter0), .b(s_4), .O(gate36inter1));
  and2  gate233(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate234(.a(s_4), .O(gate36inter3));
  inv1  gate235(.a(s_5), .O(gate36inter4));
  nand2 gate236(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate237(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate238(.a(N101), .O(gate36inter7));
  inv1  gate239(.a(N117), .O(gate36inter8));
  nand2 gate240(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate241(.a(s_5), .b(gate36inter3), .O(gate36inter10));
  nor2  gate242(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate243(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate244(.a(gate36inter12), .b(gate36inter1), .O(N285));
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );

  xor2  gate469(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate470(.a(gate40inter0), .b(s_38), .O(gate40inter1));
  and2  gate471(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate472(.a(s_38), .O(gate40inter3));
  inv1  gate473(.a(s_39), .O(gate40inter4));
  nand2 gate474(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate475(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate476(.a(N109), .O(gate40inter7));
  inv1  gate477(.a(N125), .O(gate40inter8));
  nand2 gate478(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate479(.a(s_39), .b(gate40inter3), .O(gate40inter10));
  nor2  gate480(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate481(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate482(.a(gate40inter12), .b(gate40inter1), .O(N289));
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate805(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate806(.a(gate42inter0), .b(s_86), .O(gate42inter1));
  and2  gate807(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate808(.a(s_86), .O(gate42inter3));
  inv1  gate809(.a(s_87), .O(gate42inter4));
  nand2 gate810(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate811(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate812(.a(N252), .O(gate42inter7));
  inv1  gate813(.a(N253), .O(gate42inter8));
  nand2 gate814(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate815(.a(s_87), .b(gate42inter3), .O(gate42inter10));
  nor2  gate816(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate817(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate818(.a(gate42inter12), .b(gate42inter1), .O(N293));
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );

  xor2  gate343(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate344(.a(gate46inter0), .b(s_20), .O(gate46inter1));
  and2  gate345(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate346(.a(s_20), .O(gate46inter3));
  inv1  gate347(.a(s_21), .O(gate46inter4));
  nand2 gate348(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate349(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate350(.a(N260), .O(gate46inter7));
  inv1  gate351(.a(N261), .O(gate46inter8));
  nand2 gate352(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate353(.a(s_21), .b(gate46inter3), .O(gate46inter10));
  nor2  gate354(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate355(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate356(.a(gate46inter12), .b(gate46inter1), .O(N305));

  xor2  gate819(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate820(.a(gate47inter0), .b(s_88), .O(gate47inter1));
  and2  gate821(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate822(.a(s_88), .O(gate47inter3));
  inv1  gate823(.a(s_89), .O(gate47inter4));
  nand2 gate824(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate825(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate826(.a(N262), .O(gate47inter7));
  inv1  gate827(.a(N263), .O(gate47inter8));
  nand2 gate828(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate829(.a(s_89), .b(gate47inter3), .O(gate47inter10));
  nor2  gate830(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate831(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate832(.a(gate47inter12), .b(gate47inter1), .O(N308));

  xor2  gate749(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate750(.a(gate48inter0), .b(s_78), .O(gate48inter1));
  and2  gate751(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate752(.a(s_78), .O(gate48inter3));
  inv1  gate753(.a(s_79), .O(gate48inter4));
  nand2 gate754(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate755(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate756(.a(N264), .O(gate48inter7));
  inv1  gate757(.a(N265), .O(gate48inter8));
  nand2 gate758(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate759(.a(s_79), .b(gate48inter3), .O(gate48inter10));
  nor2  gate760(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate761(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate762(.a(gate48inter12), .b(gate48inter1), .O(N311));

  xor2  gate735(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate736(.a(gate49inter0), .b(s_76), .O(gate49inter1));
  and2  gate737(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate738(.a(s_76), .O(gate49inter3));
  inv1  gate739(.a(s_77), .O(gate49inter4));
  nand2 gate740(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate741(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate742(.a(N274), .O(gate49inter7));
  inv1  gate743(.a(N275), .O(gate49inter8));
  nand2 gate744(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate745(.a(s_77), .b(gate49inter3), .O(gate49inter10));
  nor2  gate746(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate747(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate748(.a(gate49inter12), .b(gate49inter1), .O(N314));
xor2 gate50( .a(N276), .b(N277), .O(N315) );

  xor2  gate455(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate456(.a(gate51inter0), .b(s_36), .O(gate51inter1));
  and2  gate457(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate458(.a(s_36), .O(gate51inter3));
  inv1  gate459(.a(s_37), .O(gate51inter4));
  nand2 gate460(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate461(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate462(.a(N278), .O(gate51inter7));
  inv1  gate463(.a(N279), .O(gate51inter8));
  nand2 gate464(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate465(.a(s_37), .b(gate51inter3), .O(gate51inter10));
  nor2  gate466(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate467(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate468(.a(gate51inter12), .b(gate51inter1), .O(N316));

  xor2  gate525(.a(N281), .b(N280), .O(gate52inter0));
  nand2 gate526(.a(gate52inter0), .b(s_46), .O(gate52inter1));
  and2  gate527(.a(N281), .b(N280), .O(gate52inter2));
  inv1  gate528(.a(s_46), .O(gate52inter3));
  inv1  gate529(.a(s_47), .O(gate52inter4));
  nand2 gate530(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate531(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate532(.a(N280), .O(gate52inter7));
  inv1  gate533(.a(N281), .O(gate52inter8));
  nand2 gate534(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate535(.a(s_47), .b(gate52inter3), .O(gate52inter10));
  nor2  gate536(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate537(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate538(.a(gate52inter12), .b(gate52inter1), .O(N317));

  xor2  gate707(.a(N283), .b(N282), .O(gate53inter0));
  nand2 gate708(.a(gate53inter0), .b(s_72), .O(gate53inter1));
  and2  gate709(.a(N283), .b(N282), .O(gate53inter2));
  inv1  gate710(.a(s_72), .O(gate53inter3));
  inv1  gate711(.a(s_73), .O(gate53inter4));
  nand2 gate712(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate713(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate714(.a(N282), .O(gate53inter7));
  inv1  gate715(.a(N283), .O(gate53inter8));
  nand2 gate716(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate717(.a(s_73), .b(gate53inter3), .O(gate53inter10));
  nor2  gate718(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate719(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate720(.a(gate53inter12), .b(gate53inter1), .O(N318));

  xor2  gate567(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate568(.a(gate54inter0), .b(s_52), .O(gate54inter1));
  and2  gate569(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate570(.a(s_52), .O(gate54inter3));
  inv1  gate571(.a(s_53), .O(gate54inter4));
  nand2 gate572(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate573(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate574(.a(N284), .O(gate54inter7));
  inv1  gate575(.a(N285), .O(gate54inter8));
  nand2 gate576(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate577(.a(s_53), .b(gate54inter3), .O(gate54inter10));
  nor2  gate578(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate579(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate580(.a(gate54inter12), .b(gate54inter1), .O(N319));
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );

  xor2  gate399(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate400(.a(gate60inter0), .b(s_28), .O(gate60inter1));
  and2  gate401(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate402(.a(s_28), .O(gate60inter3));
  inv1  gate403(.a(s_29), .O(gate60inter4));
  nand2 gate404(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate405(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate406(.a(N293), .O(gate60inter7));
  inv1  gate407(.a(N299), .O(gate60inter8));
  nand2 gate408(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate409(.a(s_29), .b(gate60inter3), .O(gate60inter10));
  nor2  gate410(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate411(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate412(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate315(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate316(.a(gate62inter0), .b(s_16), .O(gate62inter1));
  and2  gate317(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate318(.a(s_16), .O(gate62inter3));
  inv1  gate319(.a(s_17), .O(gate62inter4));
  nand2 gate320(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate321(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate322(.a(N308), .O(gate62inter7));
  inv1  gate323(.a(N311), .O(gate62inter8));
  nand2 gate324(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate325(.a(s_17), .b(gate62inter3), .O(gate62inter10));
  nor2  gate326(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate327(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate328(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );

  xor2  gate595(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate596(.a(gate64inter0), .b(s_56), .O(gate64inter1));
  and2  gate597(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate598(.a(s_56), .O(gate64inter3));
  inv1  gate599(.a(s_57), .O(gate64inter4));
  nand2 gate600(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate601(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate602(.a(N305), .O(gate64inter7));
  inv1  gate603(.a(N311), .O(gate64inter8));
  nand2 gate604(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate605(.a(s_57), .b(gate64inter3), .O(gate64inter10));
  nor2  gate606(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate607(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate608(.a(gate64inter12), .b(gate64inter1), .O(N345));
xor2 gate65( .a(N266), .b(N342), .O(N346) );

  xor2  gate679(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate680(.a(gate66inter0), .b(s_68), .O(gate66inter1));
  and2  gate681(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate682(.a(s_68), .O(gate66inter3));
  inv1  gate683(.a(s_69), .O(gate66inter4));
  nand2 gate684(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate685(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate686(.a(N267), .O(gate66inter7));
  inv1  gate687(.a(N343), .O(gate66inter8));
  nand2 gate688(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate689(.a(s_69), .b(gate66inter3), .O(gate66inter10));
  nor2  gate690(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate691(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate692(.a(gate66inter12), .b(gate66inter1), .O(N347));
xor2 gate67( .a(N268), .b(N344), .O(N348) );

  xor2  gate665(.a(N345), .b(N269), .O(gate68inter0));
  nand2 gate666(.a(gate68inter0), .b(s_66), .O(gate68inter1));
  and2  gate667(.a(N345), .b(N269), .O(gate68inter2));
  inv1  gate668(.a(s_66), .O(gate68inter3));
  inv1  gate669(.a(s_67), .O(gate68inter4));
  nand2 gate670(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate671(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate672(.a(N269), .O(gate68inter7));
  inv1  gate673(.a(N345), .O(gate68inter8));
  nand2 gate674(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate675(.a(s_67), .b(gate68inter3), .O(gate68inter10));
  nor2  gate676(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate677(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate678(.a(gate68inter12), .b(gate68inter1), .O(N349));
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate287(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate288(.a(gate70inter0), .b(s_12), .O(gate70inter1));
  and2  gate289(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate290(.a(s_12), .O(gate70inter3));
  inv1  gate291(.a(s_13), .O(gate70inter4));
  nand2 gate292(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate293(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate294(.a(N271), .O(gate70inter7));
  inv1  gate295(.a(N339), .O(gate70inter8));
  nand2 gate296(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate297(.a(s_13), .b(gate70inter3), .O(gate70inter10));
  nor2  gate298(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate299(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate300(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );

  xor2  gate539(.a(N341), .b(N273), .O(gate72inter0));
  nand2 gate540(.a(gate72inter0), .b(s_48), .O(gate72inter1));
  and2  gate541(.a(N341), .b(N273), .O(gate72inter2));
  inv1  gate542(.a(s_48), .O(gate72inter3));
  inv1  gate543(.a(s_49), .O(gate72inter4));
  nand2 gate544(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate545(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate546(.a(N273), .O(gate72inter7));
  inv1  gate547(.a(N341), .O(gate72inter8));
  nand2 gate548(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate549(.a(s_49), .b(gate72inter3), .O(gate72inter10));
  nor2  gate550(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate551(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate552(.a(gate72inter12), .b(gate72inter1), .O(N353));
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );

  xor2  gate203(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate204(.a(gate76inter0), .b(s_0), .O(gate76inter1));
  and2  gate205(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate206(.a(s_0), .O(gate76inter3));
  inv1  gate207(.a(s_1), .O(gate76inter4));
  nand2 gate208(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate209(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate210(.a(N317), .O(gate76inter7));
  inv1  gate211(.a(N349), .O(gate76inter8));
  nand2 gate212(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate213(.a(s_1), .b(gate76inter3), .O(gate76inter10));
  nor2  gate214(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate215(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate216(.a(gate76inter12), .b(gate76inter1), .O(N393));

  xor2  gate497(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate498(.a(gate77inter0), .b(s_42), .O(gate77inter1));
  and2  gate499(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate500(.a(s_42), .O(gate77inter3));
  inv1  gate501(.a(s_43), .O(gate77inter4));
  nand2 gate502(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate503(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate504(.a(N318), .O(gate77inter7));
  inv1  gate505(.a(N350), .O(gate77inter8));
  nand2 gate506(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate507(.a(s_43), .b(gate77inter3), .O(gate77inter10));
  nor2  gate508(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate509(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate510(.a(gate77inter12), .b(gate77inter1), .O(N406));

  xor2  gate441(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate442(.a(gate78inter0), .b(s_34), .O(gate78inter1));
  and2  gate443(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate444(.a(s_34), .O(gate78inter3));
  inv1  gate445(.a(s_35), .O(gate78inter4));
  nand2 gate446(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate447(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate448(.a(N319), .O(gate78inter7));
  inv1  gate449(.a(N351), .O(gate78inter8));
  nand2 gate450(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate451(.a(s_35), .b(gate78inter3), .O(gate78inter10));
  nor2  gate452(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate453(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate454(.a(gate78inter12), .b(gate78inter1), .O(N419));
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate329(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate330(.a(gate172inter0), .b(s_18), .O(gate172inter1));
  and2  gate331(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate332(.a(s_18), .O(gate172inter3));
  inv1  gate333(.a(s_19), .O(gate172inter4));
  nand2 gate334(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate335(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate336(.a(N5), .O(gate172inter7));
  inv1  gate337(.a(N693), .O(gate172inter8));
  nand2 gate338(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate339(.a(s_19), .b(gate172inter3), .O(gate172inter10));
  nor2  gate340(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate341(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate342(.a(gate172inter12), .b(gate172inter1), .O(N725));

  xor2  gate763(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate764(.a(gate173inter0), .b(s_80), .O(gate173inter1));
  and2  gate765(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate766(.a(s_80), .O(gate173inter3));
  inv1  gate767(.a(s_81), .O(gate173inter4));
  nand2 gate768(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate769(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate770(.a(N9), .O(gate173inter7));
  inv1  gate771(.a(N694), .O(gate173inter8));
  nand2 gate772(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate773(.a(s_81), .b(gate173inter3), .O(gate173inter10));
  nor2  gate774(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate775(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate776(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate413(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate414(.a(gate176inter0), .b(s_30), .O(gate176inter1));
  and2  gate415(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate416(.a(s_30), .O(gate176inter3));
  inv1  gate417(.a(s_31), .O(gate176inter4));
  nand2 gate418(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate419(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate420(.a(N21), .O(gate176inter7));
  inv1  gate421(.a(N697), .O(gate176inter8));
  nand2 gate422(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate423(.a(s_31), .b(gate176inter3), .O(gate176inter10));
  nor2  gate424(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate425(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate426(.a(gate176inter12), .b(gate176inter1), .O(N729));

  xor2  gate581(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate582(.a(gate177inter0), .b(s_54), .O(gate177inter1));
  and2  gate583(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate584(.a(s_54), .O(gate177inter3));
  inv1  gate585(.a(s_55), .O(gate177inter4));
  nand2 gate586(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate587(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate588(.a(N25), .O(gate177inter7));
  inv1  gate589(.a(N698), .O(gate177inter8));
  nand2 gate590(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate591(.a(s_55), .b(gate177inter3), .O(gate177inter10));
  nor2  gate592(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate593(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate594(.a(gate177inter12), .b(gate177inter1), .O(N730));

  xor2  gate623(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate624(.a(gate178inter0), .b(s_60), .O(gate178inter1));
  and2  gate625(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate626(.a(s_60), .O(gate178inter3));
  inv1  gate627(.a(s_61), .O(gate178inter4));
  nand2 gate628(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate629(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate630(.a(N29), .O(gate178inter7));
  inv1  gate631(.a(N699), .O(gate178inter8));
  nand2 gate632(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate633(.a(s_61), .b(gate178inter3), .O(gate178inter10));
  nor2  gate634(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate635(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate636(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );

  xor2  gate385(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate386(.a(gate183inter0), .b(s_26), .O(gate183inter1));
  and2  gate387(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate388(.a(s_26), .O(gate183inter3));
  inv1  gate389(.a(s_27), .O(gate183inter4));
  nand2 gate390(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate391(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate392(.a(N49), .O(gate183inter7));
  inv1  gate393(.a(N704), .O(gate183inter8));
  nand2 gate394(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate395(.a(s_27), .b(gate183inter3), .O(gate183inter10));
  nor2  gate396(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate397(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate398(.a(gate183inter12), .b(gate183inter1), .O(N736));

  xor2  gate245(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate246(.a(gate184inter0), .b(s_6), .O(gate184inter1));
  and2  gate247(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate248(.a(s_6), .O(gate184inter3));
  inv1  gate249(.a(s_7), .O(gate184inter4));
  nand2 gate250(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate251(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate252(.a(N53), .O(gate184inter7));
  inv1  gate253(.a(N705), .O(gate184inter8));
  nand2 gate254(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate255(.a(s_7), .b(gate184inter3), .O(gate184inter10));
  nor2  gate256(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate257(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate258(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate483(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate484(.a(gate186inter0), .b(s_40), .O(gate186inter1));
  and2  gate485(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate486(.a(s_40), .O(gate186inter3));
  inv1  gate487(.a(s_41), .O(gate186inter4));
  nand2 gate488(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate489(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate490(.a(N61), .O(gate186inter7));
  inv1  gate491(.a(N707), .O(gate186inter8));
  nand2 gate492(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate493(.a(s_41), .b(gate186inter3), .O(gate186inter10));
  nor2  gate494(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate495(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate496(.a(gate186inter12), .b(gate186inter1), .O(N739));

  xor2  gate609(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate610(.a(gate187inter0), .b(s_58), .O(gate187inter1));
  and2  gate611(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate612(.a(s_58), .O(gate187inter3));
  inv1  gate613(.a(s_59), .O(gate187inter4));
  nand2 gate614(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate615(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate616(.a(N65), .O(gate187inter7));
  inv1  gate617(.a(N708), .O(gate187inter8));
  nand2 gate618(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate619(.a(s_59), .b(gate187inter3), .O(gate187inter10));
  nor2  gate620(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate621(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate622(.a(gate187inter12), .b(gate187inter1), .O(N740));

  xor2  gate511(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate512(.a(gate188inter0), .b(s_44), .O(gate188inter1));
  and2  gate513(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate514(.a(s_44), .O(gate188inter3));
  inv1  gate515(.a(s_45), .O(gate188inter4));
  nand2 gate516(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate517(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate518(.a(N69), .O(gate188inter7));
  inv1  gate519(.a(N709), .O(gate188inter8));
  nand2 gate520(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate521(.a(s_45), .b(gate188inter3), .O(gate188inter10));
  nor2  gate522(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate523(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate524(.a(gate188inter12), .b(gate188inter1), .O(N741));
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );

  xor2  gate637(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate638(.a(gate192inter0), .b(s_62), .O(gate192inter1));
  and2  gate639(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate640(.a(s_62), .O(gate192inter3));
  inv1  gate641(.a(s_63), .O(gate192inter4));
  nand2 gate642(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate643(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate644(.a(N85), .O(gate192inter7));
  inv1  gate645(.a(N713), .O(gate192inter8));
  nand2 gate646(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate647(.a(s_63), .b(gate192inter3), .O(gate192inter10));
  nor2  gate648(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate649(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate650(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );

  xor2  gate259(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate260(.a(gate195inter0), .b(s_8), .O(gate195inter1));
  and2  gate261(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate262(.a(s_8), .O(gate195inter3));
  inv1  gate263(.a(s_9), .O(gate195inter4));
  nand2 gate264(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate265(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate266(.a(N97), .O(gate195inter7));
  inv1  gate267(.a(N716), .O(gate195inter8));
  nand2 gate268(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate269(.a(s_9), .b(gate195inter3), .O(gate195inter10));
  nor2  gate270(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate271(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate272(.a(gate195inter12), .b(gate195inter1), .O(N748));
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );

  xor2  gate553(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate554(.a(gate199inter0), .b(s_50), .O(gate199inter1));
  and2  gate555(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate556(.a(s_50), .O(gate199inter3));
  inv1  gate557(.a(s_51), .O(gate199inter4));
  nand2 gate558(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate559(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate560(.a(N113), .O(gate199inter7));
  inv1  gate561(.a(N720), .O(gate199inter8));
  nand2 gate562(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate563(.a(s_51), .b(gate199inter3), .O(gate199inter10));
  nor2  gate564(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate565(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate566(.a(gate199inter12), .b(gate199inter1), .O(N752));
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );

  xor2  gate357(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate358(.a(gate202inter0), .b(s_22), .O(gate202inter1));
  and2  gate359(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate360(.a(s_22), .O(gate202inter3));
  inv1  gate361(.a(s_23), .O(gate202inter4));
  nand2 gate362(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate363(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate364(.a(N125), .O(gate202inter7));
  inv1  gate365(.a(N723), .O(gate202inter8));
  nand2 gate366(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate367(.a(s_23), .b(gate202inter3), .O(gate202inter10));
  nor2  gate368(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate369(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate370(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule