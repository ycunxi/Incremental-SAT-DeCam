module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate775inter0, gate775inter1, gate775inter2, gate775inter3, gate775inter4, gate775inter5, gate775inter6, gate775inter7, gate775inter8, gate775inter9, gate775inter10, gate775inter11, gate775inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate530inter0, gate530inter1, gate530inter2, gate530inter3, gate530inter4, gate530inter5, gate530inter6, gate530inter7, gate530inter8, gate530inter9, gate530inter10, gate530inter11, gate530inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate374inter0, gate374inter1, gate374inter2, gate374inter3, gate374inter4, gate374inter5, gate374inter6, gate374inter7, gate374inter8, gate374inter9, gate374inter10, gate374inter11, gate374inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate632inter0, gate632inter1, gate632inter2, gate632inter3, gate632inter4, gate632inter5, gate632inter6, gate632inter7, gate632inter8, gate632inter9, gate632inter10, gate632inter11, gate632inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate866inter0, gate866inter1, gate866inter2, gate866inter3, gate866inter4, gate866inter5, gate866inter6, gate866inter7, gate866inter8, gate866inter9, gate866inter10, gate866inter11, gate866inter12, gate586inter0, gate586inter1, gate586inter2, gate586inter3, gate586inter4, gate586inter5, gate586inter6, gate586inter7, gate586inter8, gate586inter9, gate586inter10, gate586inter11, gate586inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate605inter0, gate605inter1, gate605inter2, gate605inter3, gate605inter4, gate605inter5, gate605inter6, gate605inter7, gate605inter8, gate605inter9, gate605inter10, gate605inter11, gate605inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate528inter0, gate528inter1, gate528inter2, gate528inter3, gate528inter4, gate528inter5, gate528inter6, gate528inter7, gate528inter8, gate528inter9, gate528inter10, gate528inter11, gate528inter12, gate682inter0, gate682inter1, gate682inter2, gate682inter3, gate682inter4, gate682inter5, gate682inter6, gate682inter7, gate682inter8, gate682inter9, gate682inter10, gate682inter11, gate682inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate786inter0, gate786inter1, gate786inter2, gate786inter3, gate786inter4, gate786inter5, gate786inter6, gate786inter7, gate786inter8, gate786inter9, gate786inter10, gate786inter11, gate786inter12, gate539inter0, gate539inter1, gate539inter2, gate539inter3, gate539inter4, gate539inter5, gate539inter6, gate539inter7, gate539inter8, gate539inter9, gate539inter10, gate539inter11, gate539inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate536inter0, gate536inter1, gate536inter2, gate536inter3, gate536inter4, gate536inter5, gate536inter6, gate536inter7, gate536inter8, gate536inter9, gate536inter10, gate536inter11, gate536inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate618inter0, gate618inter1, gate618inter2, gate618inter3, gate618inter4, gate618inter5, gate618inter6, gate618inter7, gate618inter8, gate618inter9, gate618inter10, gate618inter11, gate618inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate550inter0, gate550inter1, gate550inter2, gate550inter3, gate550inter4, gate550inter5, gate550inter6, gate550inter7, gate550inter8, gate550inter9, gate550inter10, gate550inter11, gate550inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate800inter0, gate800inter1, gate800inter2, gate800inter3, gate800inter4, gate800inter5, gate800inter6, gate800inter7, gate800inter8, gate800inter9, gate800inter10, gate800inter11, gate800inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate329inter0, gate329inter1, gate329inter2, gate329inter3, gate329inter4, gate329inter5, gate329inter6, gate329inter7, gate329inter8, gate329inter9, gate329inter10, gate329inter11, gate329inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate841inter0, gate841inter1, gate841inter2, gate841inter3, gate841inter4, gate841inter5, gate841inter6, gate841inter7, gate841inter8, gate841inter9, gate841inter10, gate841inter11, gate841inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate516inter0, gate516inter1, gate516inter2, gate516inter3, gate516inter4, gate516inter5, gate516inter6, gate516inter7, gate516inter8, gate516inter9, gate516inter10, gate516inter11, gate516inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate570inter0, gate570inter1, gate570inter2, gate570inter3, gate570inter4, gate570inter5, gate570inter6, gate570inter7, gate570inter8, gate570inter9, gate570inter10, gate570inter11, gate570inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate665inter0, gate665inter1, gate665inter2, gate665inter3, gate665inter4, gate665inter5, gate665inter6, gate665inter7, gate665inter8, gate665inter9, gate665inter10, gate665inter11, gate665inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate336inter0, gate336inter1, gate336inter2, gate336inter3, gate336inter4, gate336inter5, gate336inter6, gate336inter7, gate336inter8, gate336inter9, gate336inter10, gate336inter11, gate336inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate765inter0, gate765inter1, gate765inter2, gate765inter3, gate765inter4, gate765inter5, gate765inter6, gate765inter7, gate765inter8, gate765inter9, gate765inter10, gate765inter11, gate765inter12, gate380inter0, gate380inter1, gate380inter2, gate380inter3, gate380inter4, gate380inter5, gate380inter6, gate380inter7, gate380inter8, gate380inter9, gate380inter10, gate380inter11, gate380inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate855inter0, gate855inter1, gate855inter2, gate855inter3, gate855inter4, gate855inter5, gate855inter6, gate855inter7, gate855inter8, gate855inter9, gate855inter10, gate855inter11, gate855inter12, gate762inter0, gate762inter1, gate762inter2, gate762inter3, gate762inter4, gate762inter5, gate762inter6, gate762inter7, gate762inter8, gate762inter9, gate762inter10, gate762inter11, gate762inter12, gate319inter0, gate319inter1, gate319inter2, gate319inter3, gate319inter4, gate319inter5, gate319inter6, gate319inter7, gate319inter8, gate319inter9, gate319inter10, gate319inter11, gate319inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate355inter0, gate355inter1, gate355inter2, gate355inter3, gate355inter4, gate355inter5, gate355inter6, gate355inter7, gate355inter8, gate355inter9, gate355inter10, gate355inter11, gate355inter12, gate842inter0, gate842inter1, gate842inter2, gate842inter3, gate842inter4, gate842inter5, gate842inter6, gate842inter7, gate842inter8, gate842inter9, gate842inter10, gate842inter11, gate842inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate816inter0, gate816inter1, gate816inter2, gate816inter3, gate816inter4, gate816inter5, gate816inter6, gate816inter7, gate816inter8, gate816inter9, gate816inter10, gate816inter11, gate816inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate868inter0, gate868inter1, gate868inter2, gate868inter3, gate868inter4, gate868inter5, gate868inter6, gate868inter7, gate868inter8, gate868inter9, gate868inter10, gate868inter11, gate868inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate353inter0, gate353inter1, gate353inter2, gate353inter3, gate353inter4, gate353inter5, gate353inter6, gate353inter7, gate353inter8, gate353inter9, gate353inter10, gate353inter11, gate353inter12, gate837inter0, gate837inter1, gate837inter2, gate837inter3, gate837inter4, gate837inter5, gate837inter6, gate837inter7, gate837inter8, gate837inter9, gate837inter10, gate837inter11, gate837inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate338inter0, gate338inter1, gate338inter2, gate338inter3, gate338inter4, gate338inter5, gate338inter6, gate338inter7, gate338inter8, gate338inter9, gate338inter10, gate338inter11, gate338inter12, gate372inter0, gate372inter1, gate372inter2, gate372inter3, gate372inter4, gate372inter5, gate372inter6, gate372inter7, gate372inter8, gate372inter9, gate372inter10, gate372inter11, gate372inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate361inter0, gate361inter1, gate361inter2, gate361inter3, gate361inter4, gate361inter5, gate361inter6, gate361inter7, gate361inter8, gate361inter9, gate361inter10, gate361inter11, gate361inter12, gate341inter0, gate341inter1, gate341inter2, gate341inter3, gate341inter4, gate341inter5, gate341inter6, gate341inter7, gate341inter8, gate341inter9, gate341inter10, gate341inter11, gate341inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate769inter0, gate769inter1, gate769inter2, gate769inter3, gate769inter4, gate769inter5, gate769inter6, gate769inter7, gate769inter8, gate769inter9, gate769inter10, gate769inter11, gate769inter12, gate851inter0, gate851inter1, gate851inter2, gate851inter3, gate851inter4, gate851inter5, gate851inter6, gate851inter7, gate851inter8, gate851inter9, gate851inter10, gate851inter11, gate851inter12, gate820inter0, gate820inter1, gate820inter2, gate820inter3, gate820inter4, gate820inter5, gate820inter6, gate820inter7, gate820inter8, gate820inter9, gate820inter10, gate820inter11, gate820inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate681inter0, gate681inter1, gate681inter2, gate681inter3, gate681inter4, gate681inter5, gate681inter6, gate681inter7, gate681inter8, gate681inter9, gate681inter10, gate681inter11, gate681inter12, gate357inter0, gate357inter1, gate357inter2, gate357inter3, gate357inter4, gate357inter5, gate357inter6, gate357inter7, gate357inter8, gate357inter9, gate357inter10, gate357inter11, gate357inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate1105(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate1106(.a(gate17inter0), .b(s_32), .O(gate17inter1));
  and2  gate1107(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate1108(.a(s_32), .O(gate17inter3));
  inv1  gate1109(.a(s_33), .O(gate17inter4));
  nand2 gate1110(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1111(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1112(.a(N63), .O(gate17inter7));
  inv1  gate1113(.a(N88), .O(gate17inter8));
  nand2 gate1114(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1115(.a(s_33), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1116(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1117(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1118(.a(gate17inter12), .b(gate17inter1), .O(N251));
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );

  xor2  gate1427(.a(N331), .b(N306), .O(gate75inter0));
  nand2 gate1428(.a(gate75inter0), .b(s_78), .O(gate75inter1));
  and2  gate1429(.a(N331), .b(N306), .O(gate75inter2));
  inv1  gate1430(.a(s_78), .O(gate75inter3));
  inv1  gate1431(.a(s_79), .O(gate75inter4));
  nand2 gate1432(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1433(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1434(.a(N306), .O(gate75inter7));
  inv1  gate1435(.a(N331), .O(gate75inter8));
  nand2 gate1436(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1437(.a(s_79), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1438(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1439(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1440(.a(gate75inter12), .b(gate75inter1), .O(N550));
nand2 gate76( .a(N306), .b(N331), .O(N551) );

  xor2  gate1805(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate1806(.a(gate77inter0), .b(s_132), .O(gate77inter1));
  and2  gate1807(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate1808(.a(s_132), .O(gate77inter3));
  inv1  gate1809(.a(s_133), .O(gate77inter4));
  nand2 gate1810(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1811(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1812(.a(N306), .O(gate77inter7));
  inv1  gate1813(.a(N331), .O(gate77inter8));
  nand2 gate1814(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1815(.a(s_133), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1816(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1817(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1818(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );

  xor2  gate909(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate910(.a(gate79inter0), .b(s_4), .O(gate79inter1));
  and2  gate911(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate912(.a(s_4), .O(gate79inter3));
  inv1  gate913(.a(s_5), .O(gate79inter4));
  nand2 gate914(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate915(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate916(.a(N306), .O(gate79inter7));
  inv1  gate917(.a(N331), .O(gate79inter8));
  nand2 gate918(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate919(.a(s_5), .b(gate79inter3), .O(gate79inter10));
  nor2  gate920(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate921(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate922(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );

  xor2  gate1959(.a(N280), .b(N326), .O(gate97inter0));
  nand2 gate1960(.a(gate97inter0), .b(s_154), .O(gate97inter1));
  and2  gate1961(.a(N280), .b(N326), .O(gate97inter2));
  inv1  gate1962(.a(s_154), .O(gate97inter3));
  inv1  gate1963(.a(s_155), .O(gate97inter4));
  nand2 gate1964(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1965(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1966(.a(N326), .O(gate97inter7));
  inv1  gate1967(.a(N280), .O(gate97inter8));
  nand2 gate1968(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1969(.a(s_155), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1970(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1971(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1972(.a(gate97inter12), .b(gate97inter1), .O(N602));

  xor2  gate1063(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate1064(.a(gate98inter0), .b(s_26), .O(gate98inter1));
  and2  gate1065(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate1066(.a(s_26), .O(gate98inter3));
  inv1  gate1067(.a(s_27), .O(gate98inter4));
  nand2 gate1068(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1069(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1070(.a(N260), .O(gate98inter7));
  inv1  gate1071(.a(N72), .O(gate98inter8));
  nand2 gate1072(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1073(.a(s_27), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1074(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1075(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1076(.a(gate98inter12), .b(gate98inter1), .O(N603));
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );

  xor2  gate1399(.a(N612), .b(N53), .O(gate160inter0));
  nand2 gate1400(.a(gate160inter0), .b(s_74), .O(gate160inter1));
  and2  gate1401(.a(N612), .b(N53), .O(gate160inter2));
  inv1  gate1402(.a(s_74), .O(gate160inter3));
  inv1  gate1403(.a(s_75), .O(gate160inter4));
  nand2 gate1404(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1405(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1406(.a(N53), .O(gate160inter7));
  inv1  gate1407(.a(N612), .O(gate160inter8));
  nand2 gate1408(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1409(.a(s_75), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1410(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1411(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1412(.a(gate160inter12), .b(gate160inter1), .O(N899));

  xor2  gate1077(.a(N608), .b(N60), .O(gate161inter0));
  nand2 gate1078(.a(gate161inter0), .b(s_28), .O(gate161inter1));
  and2  gate1079(.a(N608), .b(N60), .O(gate161inter2));
  inv1  gate1080(.a(s_28), .O(gate161inter3));
  inv1  gate1081(.a(s_29), .O(gate161inter4));
  nand2 gate1082(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1083(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1084(.a(N60), .O(gate161inter7));
  inv1  gate1085(.a(N608), .O(gate161inter8));
  nand2 gate1086(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1087(.a(s_29), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1088(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1089(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1090(.a(gate161inter12), .b(gate161inter1), .O(N903));

  xor2  gate2141(.a(N612), .b(N49), .O(gate162inter0));
  nand2 gate2142(.a(gate162inter0), .b(s_180), .O(gate162inter1));
  and2  gate2143(.a(N612), .b(N49), .O(gate162inter2));
  inv1  gate2144(.a(s_180), .O(gate162inter3));
  inv1  gate2145(.a(s_181), .O(gate162inter4));
  nand2 gate2146(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2147(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2148(.a(N49), .O(gate162inter7));
  inv1  gate2149(.a(N612), .O(gate162inter8));
  nand2 gate2150(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2151(.a(s_181), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2152(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2153(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2154(.a(gate162inter12), .b(gate162inter1), .O(N907));
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );

  xor2  gate1973(.a(N889), .b(N616), .O(gate234inter0));
  nand2 gate1974(.a(gate234inter0), .b(s_156), .O(gate234inter1));
  and2  gate1975(.a(N889), .b(N616), .O(gate234inter2));
  inv1  gate1976(.a(s_156), .O(gate234inter3));
  inv1  gate1977(.a(s_157), .O(gate234inter4));
  nand2 gate1978(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1979(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1980(.a(N616), .O(gate234inter7));
  inv1  gate1981(.a(N889), .O(gate234inter8));
  nand2 gate1982(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1983(.a(s_157), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1984(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1985(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1986(.a(gate234inter12), .b(gate234inter1), .O(N1055));

  xor2  gate993(.a(N890), .b(N625), .O(gate235inter0));
  nand2 gate994(.a(gate235inter0), .b(s_16), .O(gate235inter1));
  and2  gate995(.a(N890), .b(N625), .O(gate235inter2));
  inv1  gate996(.a(s_16), .O(gate235inter3));
  inv1  gate997(.a(s_17), .O(gate235inter4));
  nand2 gate998(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate999(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1000(.a(N625), .O(gate235inter7));
  inv1  gate1001(.a(N890), .O(gate235inter8));
  nand2 gate1002(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1003(.a(s_17), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1004(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1005(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1006(.a(gate235inter12), .b(gate235inter1), .O(N1063));

  xor2  gate1931(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate1932(.a(gate236inter0), .b(s_150), .O(gate236inter1));
  and2  gate1933(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate1934(.a(s_150), .O(gate236inter3));
  inv1  gate1935(.a(s_151), .O(gate236inter4));
  nand2 gate1936(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1937(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1938(.a(N622), .O(gate236inter7));
  inv1  gate1939(.a(N891), .O(gate236inter8));
  nand2 gate1940(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1941(.a(s_151), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1942(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1943(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1944(.a(gate236inter12), .b(gate236inter1), .O(N1064));
nand2 gate237( .a(N655), .b(N895), .O(N1067) );

  xor2  gate1035(.a(N896), .b(N652), .O(gate238inter0));
  nand2 gate1036(.a(gate238inter0), .b(s_22), .O(gate238inter1));
  and2  gate1037(.a(N896), .b(N652), .O(gate238inter2));
  inv1  gate1038(.a(s_22), .O(gate238inter3));
  inv1  gate1039(.a(s_23), .O(gate238inter4));
  nand2 gate1040(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1041(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1042(.a(N652), .O(gate238inter7));
  inv1  gate1043(.a(N896), .O(gate238inter8));
  nand2 gate1044(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1045(.a(s_23), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1046(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1047(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1048(.a(gate238inter12), .b(gate238inter1), .O(N1068));
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );

  xor2  gate1763(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate1764(.a(gate244inter0), .b(s_126), .O(gate244inter1));
  and2  gate1765(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate1766(.a(s_126), .O(gate244inter3));
  inv1  gate1767(.a(s_127), .O(gate244inter4));
  nand2 gate1768(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1769(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1770(.a(N736), .O(gate244inter7));
  inv1  gate1771(.a(N1003), .O(gate244inter8));
  nand2 gate1772(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1773(.a(s_127), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1774(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1775(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1776(.a(gate244inter12), .b(gate244inter1), .O(N1129));
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );

  xor2  gate1553(.a(N1008), .b(N751), .O(gate247inter0));
  nand2 gate1554(.a(gate247inter0), .b(s_96), .O(gate247inter1));
  and2  gate1555(.a(N1008), .b(N751), .O(gate247inter2));
  inv1  gate1556(.a(s_96), .O(gate247inter3));
  inv1  gate1557(.a(s_97), .O(gate247inter4));
  nand2 gate1558(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1559(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1560(.a(N751), .O(gate247inter7));
  inv1  gate1561(.a(N1008), .O(gate247inter8));
  nand2 gate1562(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1563(.a(s_97), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1564(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1565(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1566(.a(gate247inter12), .b(gate247inter1), .O(N1132));
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );

  xor2  gate1749(.a(N1055), .b(N1054), .O(gate251inter0));
  nand2 gate1750(.a(gate251inter0), .b(s_124), .O(gate251inter1));
  and2  gate1751(.a(N1055), .b(N1054), .O(gate251inter2));
  inv1  gate1752(.a(s_124), .O(gate251inter3));
  inv1  gate1753(.a(s_125), .O(gate251inter4));
  nand2 gate1754(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1755(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1756(.a(N1054), .O(gate251inter7));
  inv1  gate1757(.a(N1055), .O(gate251inter8));
  nand2 gate1758(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1759(.a(s_125), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1760(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1761(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1762(.a(gate251inter12), .b(gate251inter1), .O(N1150));
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate951(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate952(.a(gate268inter0), .b(s_10), .O(gate268inter1));
  and2  gate953(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate954(.a(s_10), .O(gate268inter3));
  inv1  gate955(.a(s_11), .O(gate268inter4));
  nand2 gate956(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate957(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate958(.a(N921), .O(gate268inter7));
  inv1  gate959(.a(N923), .O(gate268inter8));
  nand2 gate960(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate961(.a(s_11), .b(gate268inter3), .O(gate268inter10));
  nor2  gate962(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate963(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate964(.a(gate268inter12), .b(gate268inter1), .O(N1171));
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate1119(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate1120(.a(gate273inter0), .b(s_34), .O(gate273inter1));
  and2  gate1121(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate1122(.a(s_34), .O(gate273inter3));
  inv1  gate1123(.a(s_35), .O(gate273inter4));
  nand2 gate1124(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1125(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1126(.a(N1013), .O(gate273inter7));
  inv1  gate1127(.a(N942), .O(gate273inter8));
  nand2 gate1128(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1129(.a(s_35), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1130(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1131(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1132(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate1371(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate1372(.a(gate275inter0), .b(s_70), .O(gate275inter1));
  and2  gate1373(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate1374(.a(s_70), .O(gate275inter3));
  inv1  gate1375(.a(s_71), .O(gate275inter4));
  nand2 gate1376(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1377(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1378(.a(N1016), .O(gate275inter7));
  inv1  gate1379(.a(N946), .O(gate275inter8));
  nand2 gate1380(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1381(.a(s_71), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1382(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1383(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1384(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate1315(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate1316(.a(gate277inter0), .b(s_62), .O(gate277inter1));
  and2  gate1317(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate1318(.a(s_62), .O(gate277inter3));
  inv1  gate1319(.a(s_63), .O(gate277inter4));
  nand2 gate1320(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1321(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1322(.a(N1019), .O(gate277inter7));
  inv1  gate1323(.a(N950), .O(gate277inter8));
  nand2 gate1324(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1325(.a(s_63), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1326(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1327(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1328(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );

  xor2  gate2155(.a(N984), .b(N981), .O(gate296inter0));
  nand2 gate2156(.a(gate296inter0), .b(s_182), .O(gate296inter1));
  and2  gate2157(.a(N984), .b(N981), .O(gate296inter2));
  inv1  gate2158(.a(s_182), .O(gate296inter3));
  inv1  gate2159(.a(s_183), .O(gate296inter4));
  nand2 gate2160(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2161(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2162(.a(N981), .O(gate296inter7));
  inv1  gate2163(.a(N984), .O(gate296inter8));
  nand2 gate2164(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2165(.a(s_183), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2166(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2167(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2168(.a(gate296inter12), .b(gate296inter1), .O(N1231));
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );

  xor2  gate1693(.a(N997), .b(N1046), .O(gate300inter0));
  nand2 gate1694(.a(gate300inter0), .b(s_116), .O(gate300inter1));
  and2  gate1695(.a(N997), .b(N1046), .O(gate300inter2));
  inv1  gate1696(.a(s_116), .O(gate300inter3));
  inv1  gate1697(.a(s_117), .O(gate300inter4));
  nand2 gate1698(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate1699(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate1700(.a(N1046), .O(gate300inter7));
  inv1  gate1701(.a(N997), .O(gate300inter8));
  nand2 gate1702(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate1703(.a(s_117), .b(gate300inter3), .O(gate300inter10));
  nor2  gate1704(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate1705(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate1706(.a(gate300inter12), .b(gate300inter1), .O(N1239));
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate1455(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate1456(.a(gate312inter0), .b(s_82), .O(gate312inter1));
  and2  gate1457(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate1458(.a(s_82), .O(gate312inter3));
  inv1  gate1459(.a(s_83), .O(gate312inter4));
  nand2 gate1460(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate1461(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate1462(.a(N631), .O(gate312inter7));
  inv1  gate1463(.a(N1159), .O(gate312inter8));
  nand2 gate1464(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate1465(.a(s_83), .b(gate312inter3), .O(gate312inter10));
  nor2  gate1466(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate1467(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate1468(.a(gate312inter12), .b(gate312inter1), .O(N1267));
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );

  xor2  gate1903(.a(N1220), .b(N706), .O(gate319inter0));
  nand2 gate1904(.a(gate319inter0), .b(s_146), .O(gate319inter1));
  and2  gate1905(.a(N1220), .b(N706), .O(gate319inter2));
  inv1  gate1906(.a(s_146), .O(gate319inter3));
  inv1  gate1907(.a(s_147), .O(gate319inter4));
  nand2 gate1908(.a(gate319inter4), .b(gate319inter3), .O(gate319inter5));
  nor2  gate1909(.a(gate319inter5), .b(gate319inter2), .O(gate319inter6));
  inv1  gate1910(.a(N706), .O(gate319inter7));
  inv1  gate1911(.a(N1220), .O(gate319inter8));
  nand2 gate1912(.a(gate319inter8), .b(gate319inter7), .O(gate319inter9));
  nand2 gate1913(.a(s_147), .b(gate319inter3), .O(gate319inter10));
  nor2  gate1914(.a(gate319inter10), .b(gate319inter9), .O(gate319inter11));
  nor2  gate1915(.a(gate319inter11), .b(gate319inter6), .O(gate319inter12));
  nand2 gate1916(.a(gate319inter12), .b(gate319inter1), .O(N1315));
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );

  xor2  gate2225(.a(N1228), .b(N715), .O(gate322inter0));
  nand2 gate2226(.a(gate322inter0), .b(s_192), .O(gate322inter1));
  and2  gate2227(.a(N1228), .b(N715), .O(gate322inter2));
  inv1  gate2228(.a(s_192), .O(gate322inter3));
  inv1  gate2229(.a(s_193), .O(gate322inter4));
  nand2 gate2230(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate2231(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate2232(.a(N715), .O(gate322inter7));
  inv1  gate2233(.a(N1228), .O(gate322inter8));
  nand2 gate2234(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate2235(.a(s_193), .b(gate322inter3), .O(gate322inter10));
  nor2  gate2236(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate2237(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate2238(.a(gate322inter12), .b(gate322inter1), .O(N1318));
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );

  xor2  gate1511(.a(N1160), .b(N1267), .O(gate328inter0));
  nand2 gate1512(.a(gate328inter0), .b(s_90), .O(gate328inter1));
  and2  gate1513(.a(N1160), .b(N1267), .O(gate328inter2));
  inv1  gate1514(.a(s_90), .O(gate328inter3));
  inv1  gate1515(.a(s_91), .O(gate328inter4));
  nand2 gate1516(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate1517(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate1518(.a(N1267), .O(gate328inter7));
  inv1  gate1519(.a(N1160), .O(gate328inter8));
  nand2 gate1520(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate1521(.a(s_91), .b(gate328inter3), .O(gate328inter10));
  nor2  gate1522(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate1523(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate1524(.a(gate328inter12), .b(gate328inter1), .O(N1344));

  xor2  gate1539(.a(N894), .b(N1249), .O(gate329inter0));
  nand2 gate1540(.a(gate329inter0), .b(s_94), .O(gate329inter1));
  and2  gate1541(.a(N894), .b(N1249), .O(gate329inter2));
  inv1  gate1542(.a(s_94), .O(gate329inter3));
  inv1  gate1543(.a(s_95), .O(gate329inter4));
  nand2 gate1544(.a(gate329inter4), .b(gate329inter3), .O(gate329inter5));
  nor2  gate1545(.a(gate329inter5), .b(gate329inter2), .O(gate329inter6));
  inv1  gate1546(.a(N1249), .O(gate329inter7));
  inv1  gate1547(.a(N894), .O(gate329inter8));
  nand2 gate1548(.a(gate329inter8), .b(gate329inter7), .O(gate329inter9));
  nand2 gate1549(.a(s_95), .b(gate329inter3), .O(gate329inter10));
  nor2  gate1550(.a(gate329inter10), .b(gate329inter9), .O(gate329inter11));
  nor2  gate1551(.a(gate329inter11), .b(gate329inter6), .O(gate329inter12));
  nand2 gate1552(.a(gate329inter12), .b(gate329inter1), .O(N1345));
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );

  xor2  gate1777(.a(N1208), .b(N1310), .O(gate336inter0));
  nand2 gate1778(.a(gate336inter0), .b(s_128), .O(gate336inter1));
  and2  gate1779(.a(N1208), .b(N1310), .O(gate336inter2));
  inv1  gate1780(.a(s_128), .O(gate336inter3));
  inv1  gate1781(.a(s_129), .O(gate336inter4));
  nand2 gate1782(.a(gate336inter4), .b(gate336inter3), .O(gate336inter5));
  nor2  gate1783(.a(gate336inter5), .b(gate336inter2), .O(gate336inter6));
  inv1  gate1784(.a(N1310), .O(gate336inter7));
  inv1  gate1785(.a(N1208), .O(gate336inter8));
  nand2 gate1786(.a(gate336inter8), .b(gate336inter7), .O(gate336inter9));
  nand2 gate1787(.a(s_129), .b(gate336inter3), .O(gate336inter10));
  nor2  gate1788(.a(gate336inter10), .b(gate336inter9), .O(gate336inter11));
  nor2  gate1789(.a(gate336inter11), .b(gate336inter6), .O(gate336inter12));
  nand2 gate1790(.a(gate336inter12), .b(gate336inter1), .O(N1355));
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );

  xor2  gate2183(.a(N1212), .b(N1312), .O(gate338inter0));
  nand2 gate2184(.a(gate338inter0), .b(s_186), .O(gate338inter1));
  and2  gate2185(.a(N1212), .b(N1312), .O(gate338inter2));
  inv1  gate2186(.a(s_186), .O(gate338inter3));
  inv1  gate2187(.a(s_187), .O(gate338inter4));
  nand2 gate2188(.a(gate338inter4), .b(gate338inter3), .O(gate338inter5));
  nor2  gate2189(.a(gate338inter5), .b(gate338inter2), .O(gate338inter6));
  inv1  gate2190(.a(N1312), .O(gate338inter7));
  inv1  gate2191(.a(N1212), .O(gate338inter8));
  nand2 gate2192(.a(gate338inter8), .b(gate338inter7), .O(gate338inter9));
  nand2 gate2193(.a(s_187), .b(gate338inter3), .O(gate338inter10));
  nor2  gate2194(.a(gate338inter10), .b(gate338inter9), .O(gate338inter11));
  nor2  gate2195(.a(gate338inter11), .b(gate338inter6), .O(gate338inter12));
  nand2 gate2196(.a(gate338inter12), .b(gate338inter1), .O(N1361));
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );

  xor2  gate2253(.a(N1221), .b(N1315), .O(gate341inter0));
  nand2 gate2254(.a(gate341inter0), .b(s_196), .O(gate341inter1));
  and2  gate2255(.a(N1221), .b(N1315), .O(gate341inter2));
  inv1  gate2256(.a(s_196), .O(gate341inter3));
  inv1  gate2257(.a(s_197), .O(gate341inter4));
  nand2 gate2258(.a(gate341inter4), .b(gate341inter3), .O(gate341inter5));
  nor2  gate2259(.a(gate341inter5), .b(gate341inter2), .O(gate341inter6));
  inv1  gate2260(.a(N1315), .O(gate341inter7));
  inv1  gate2261(.a(N1221), .O(gate341inter8));
  nand2 gate2262(.a(gate341inter8), .b(gate341inter7), .O(gate341inter9));
  nand2 gate2263(.a(s_197), .b(gate341inter3), .O(gate341inter10));
  nor2  gate2264(.a(gate341inter10), .b(gate341inter9), .O(gate341inter11));
  nor2  gate2265(.a(gate341inter11), .b(gate341inter6), .O(gate341inter12));
  nand2 gate2266(.a(gate341inter12), .b(gate341inter1), .O(N1370));

  xor2  gate937(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate938(.a(gate342inter0), .b(s_8), .O(gate342inter1));
  and2  gate939(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate940(.a(s_8), .O(gate342inter3));
  inv1  gate941(.a(s_9), .O(gate342inter4));
  nand2 gate942(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate943(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate944(.a(N1316), .O(gate342inter7));
  inv1  gate945(.a(N1224), .O(gate342inter8));
  nand2 gate946(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate947(.a(s_9), .b(gate342inter3), .O(gate342inter10));
  nor2  gate948(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate949(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate950(.a(gate342inter12), .b(gate342inter1), .O(N1373));
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );

  xor2  gate1049(.a(N1229), .b(N1318), .O(gate344inter0));
  nand2 gate1050(.a(gate344inter0), .b(s_24), .O(gate344inter1));
  and2  gate1051(.a(N1229), .b(N1318), .O(gate344inter2));
  inv1  gate1052(.a(s_24), .O(gate344inter3));
  inv1  gate1053(.a(s_25), .O(gate344inter4));
  nand2 gate1054(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate1055(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate1056(.a(N1318), .O(gate344inter7));
  inv1  gate1057(.a(N1229), .O(gate344inter8));
  nand2 gate1058(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate1059(.a(s_25), .b(gate344inter3), .O(gate344inter10));
  nor2  gate1060(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate1061(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate1062(.a(gate344inter12), .b(gate344inter1), .O(N1379));
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );

  xor2  gate2113(.a(N1004), .b(N1243), .O(gate353inter0));
  nand2 gate2114(.a(gate353inter0), .b(s_176), .O(gate353inter1));
  and2  gate2115(.a(N1004), .b(N1243), .O(gate353inter2));
  inv1  gate2116(.a(s_176), .O(gate353inter3));
  inv1  gate2117(.a(s_177), .O(gate353inter4));
  nand2 gate2118(.a(gate353inter4), .b(gate353inter3), .O(gate353inter5));
  nor2  gate2119(.a(gate353inter5), .b(gate353inter2), .O(gate353inter6));
  inv1  gate2120(.a(N1243), .O(gate353inter7));
  inv1  gate2121(.a(N1004), .O(gate353inter8));
  nand2 gate2122(.a(gate353inter8), .b(gate353inter7), .O(gate353inter9));
  nand2 gate2123(.a(s_177), .b(gate353inter3), .O(gate353inter10));
  nor2  gate2124(.a(gate353inter10), .b(gate353inter9), .O(gate353inter11));
  nor2  gate2125(.a(gate353inter11), .b(gate353inter6), .O(gate353inter12));
  nand2 gate2126(.a(gate353inter12), .b(gate353inter1), .O(N1397));
inv1 gate354( .a(N1246), .O(N1398) );

  xor2  gate2001(.a(N1007), .b(N1246), .O(gate355inter0));
  nand2 gate2002(.a(gate355inter0), .b(s_160), .O(gate355inter1));
  and2  gate2003(.a(N1007), .b(N1246), .O(gate355inter2));
  inv1  gate2004(.a(s_160), .O(gate355inter3));
  inv1  gate2005(.a(s_161), .O(gate355inter4));
  nand2 gate2006(.a(gate355inter4), .b(gate355inter3), .O(gate355inter5));
  nor2  gate2007(.a(gate355inter5), .b(gate355inter2), .O(gate355inter6));
  inv1  gate2008(.a(N1246), .O(gate355inter7));
  inv1  gate2009(.a(N1007), .O(gate355inter8));
  nand2 gate2010(.a(gate355inter8), .b(gate355inter7), .O(gate355inter9));
  nand2 gate2011(.a(s_161), .b(gate355inter3), .O(gate355inter10));
  nor2  gate2012(.a(gate355inter10), .b(gate355inter9), .O(gate355inter11));
  nor2  gate2013(.a(gate355inter11), .b(gate355inter6), .O(gate355inter12));
  nand2 gate2014(.a(gate355inter12), .b(gate355inter1), .O(N1399));
inv1 gate356( .a(N1319), .O(N1409) );

  xor2  gate2351(.a(N1346), .b(N649), .O(gate357inter0));
  nand2 gate2352(.a(gate357inter0), .b(s_210), .O(gate357inter1));
  and2  gate2353(.a(N1346), .b(N649), .O(gate357inter2));
  inv1  gate2354(.a(s_210), .O(gate357inter3));
  inv1  gate2355(.a(s_211), .O(gate357inter4));
  nand2 gate2356(.a(gate357inter4), .b(gate357inter3), .O(gate357inter5));
  nor2  gate2357(.a(gate357inter5), .b(gate357inter2), .O(gate357inter6));
  inv1  gate2358(.a(N649), .O(gate357inter7));
  inv1  gate2359(.a(N1346), .O(gate357inter8));
  nand2 gate2360(.a(gate357inter8), .b(gate357inter7), .O(gate357inter9));
  nand2 gate2361(.a(s_211), .b(gate357inter3), .O(gate357inter10));
  nor2  gate2362(.a(gate357inter10), .b(gate357inter9), .O(gate357inter11));
  nor2  gate2363(.a(gate357inter11), .b(gate357inter6), .O(gate357inter12));
  nand2 gate2364(.a(gate357inter12), .b(gate357inter1), .O(N1412));
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );

  xor2  gate2239(.a(N1386), .b(N634), .O(gate361inter0));
  nand2 gate2240(.a(gate361inter0), .b(s_194), .O(gate361inter1));
  and2  gate2241(.a(N1386), .b(N634), .O(gate361inter2));
  inv1  gate2242(.a(s_194), .O(gate361inter3));
  inv1  gate2243(.a(s_195), .O(gate361inter4));
  nand2 gate2244(.a(gate361inter4), .b(gate361inter3), .O(gate361inter5));
  nor2  gate2245(.a(gate361inter5), .b(gate361inter2), .O(gate361inter6));
  inv1  gate2246(.a(N634), .O(gate361inter7));
  inv1  gate2247(.a(N1386), .O(gate361inter8));
  nand2 gate2248(.a(gate361inter8), .b(gate361inter7), .O(gate361inter9));
  nand2 gate2249(.a(s_195), .b(gate361inter3), .O(gate361inter10));
  nor2  gate2250(.a(gate361inter10), .b(gate361inter9), .O(gate361inter11));
  nor2  gate2251(.a(gate361inter11), .b(gate361inter6), .O(gate361inter12));
  nand2 gate2252(.a(gate361inter12), .b(gate361inter1), .O(N1433));
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );

  xor2  gate2197(.a(N1152), .b(N1361), .O(gate372inter0));
  nand2 gate2198(.a(gate372inter0), .b(s_188), .O(gate372inter1));
  and2  gate2199(.a(N1152), .b(N1361), .O(gate372inter2));
  inv1  gate2200(.a(s_188), .O(gate372inter3));
  inv1  gate2201(.a(s_189), .O(gate372inter4));
  nand2 gate2202(.a(gate372inter4), .b(gate372inter3), .O(gate372inter5));
  nor2  gate2203(.a(gate372inter5), .b(gate372inter2), .O(gate372inter6));
  inv1  gate2204(.a(N1361), .O(gate372inter7));
  inv1  gate2205(.a(N1152), .O(gate372inter8));
  nand2 gate2206(.a(gate372inter8), .b(gate372inter7), .O(gate372inter9));
  nand2 gate2207(.a(s_189), .b(gate372inter3), .O(gate372inter10));
  nor2  gate2208(.a(gate372inter10), .b(gate372inter9), .O(gate372inter11));
  nor2  gate2209(.a(gate372inter11), .b(gate372inter6), .O(gate372inter12));
  nand2 gate2210(.a(gate372inter12), .b(gate372inter1), .O(N1451));
inv1 gate373( .a(N1361), .O(N1452) );

  xor2  gate965(.a(N1153), .b(N1367), .O(gate374inter0));
  nand2 gate966(.a(gate374inter0), .b(s_12), .O(gate374inter1));
  and2  gate967(.a(N1153), .b(N1367), .O(gate374inter2));
  inv1  gate968(.a(s_12), .O(gate374inter3));
  inv1  gate969(.a(s_13), .O(gate374inter4));
  nand2 gate970(.a(gate374inter4), .b(gate374inter3), .O(gate374inter5));
  nor2  gate971(.a(gate374inter5), .b(gate374inter2), .O(gate374inter6));
  inv1  gate972(.a(N1367), .O(gate374inter7));
  inv1  gate973(.a(N1153), .O(gate374inter8));
  nand2 gate974(.a(gate374inter8), .b(gate374inter7), .O(gate374inter9));
  nand2 gate975(.a(s_13), .b(gate374inter3), .O(gate374inter10));
  nor2  gate976(.a(gate374inter10), .b(gate374inter9), .O(gate374inter11));
  nor2  gate977(.a(gate374inter11), .b(gate374inter6), .O(gate374inter12));
  nand2 gate978(.a(gate374inter12), .b(gate374inter1), .O(N1453));
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );

  xor2  gate1847(.a(N1157), .b(N1379), .O(gate380inter0));
  nand2 gate1848(.a(gate380inter0), .b(s_138), .O(gate380inter1));
  and2  gate1849(.a(N1157), .b(N1379), .O(gate380inter2));
  inv1  gate1850(.a(s_138), .O(gate380inter3));
  inv1  gate1851(.a(s_139), .O(gate380inter4));
  nand2 gate1852(.a(gate380inter4), .b(gate380inter3), .O(gate380inter5));
  nor2  gate1853(.a(gate380inter5), .b(gate380inter2), .O(gate380inter6));
  inv1  gate1854(.a(N1379), .O(gate380inter7));
  inv1  gate1855(.a(N1157), .O(gate380inter8));
  nand2 gate1856(.a(gate380inter8), .b(gate380inter7), .O(gate380inter9));
  nand2 gate1857(.a(s_139), .b(gate380inter3), .O(gate380inter10));
  nor2  gate1858(.a(gate380inter10), .b(gate380inter9), .O(gate380inter11));
  nor2  gate1859(.a(gate380inter11), .b(gate380inter6), .O(gate380inter12));
  nand2 gate1860(.a(gate380inter12), .b(gate380inter1), .O(N1459));
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );

  xor2  gate1819(.a(N1446), .b(N935), .O(gate397inter0));
  nand2 gate1820(.a(gate397inter0), .b(s_134), .O(gate397inter1));
  and2  gate1821(.a(N1446), .b(N935), .O(gate397inter2));
  inv1  gate1822(.a(s_134), .O(gate397inter3));
  inv1  gate1823(.a(s_135), .O(gate397inter4));
  nand2 gate1824(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1825(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1826(.a(N935), .O(gate397inter7));
  inv1  gate1827(.a(N1446), .O(gate397inter8));
  nand2 gate1828(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1829(.a(s_135), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1830(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1831(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1832(.a(gate397inter12), .b(gate397inter1), .O(N1488));
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );

  xor2  gate881(.a(N1452), .b(N947), .O(gate401inter0));
  nand2 gate882(.a(gate401inter0), .b(s_0), .O(gate401inter1));
  and2  gate883(.a(N1452), .b(N947), .O(gate401inter2));
  inv1  gate884(.a(s_0), .O(gate401inter3));
  inv1  gate885(.a(s_1), .O(gate401inter4));
  nand2 gate886(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate887(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate888(.a(N947), .O(gate401inter7));
  inv1  gate889(.a(N1452), .O(gate401inter8));
  nand2 gate890(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate891(.a(s_1), .b(gate401inter3), .O(gate401inter10));
  nor2  gate892(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate893(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate894(.a(gate401inter12), .b(gate401inter1), .O(N1492));

  xor2  gate1735(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate1736(.a(gate402inter0), .b(s_122), .O(gate402inter1));
  and2  gate1737(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate1738(.a(s_122), .O(gate402inter3));
  inv1  gate1739(.a(s_123), .O(gate402inter4));
  nand2 gate1740(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1741(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1742(.a(N955), .O(gate402inter7));
  inv1  gate1743(.a(N1454), .O(gate402inter8));
  nand2 gate1744(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1745(.a(s_123), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1746(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1747(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1748(.a(gate402inter12), .b(gate402inter1), .O(N1493));
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );

  xor2  gate1231(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate1232(.a(gate406inter0), .b(s_50), .O(gate406inter1));
  and2  gate1233(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate1234(.a(s_50), .O(gate406inter3));
  inv1  gate1235(.a(s_51), .O(gate406inter4));
  nand2 gate1236(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1237(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1238(.a(N998), .O(gate406inter7));
  inv1  gate1239(.a(N1463), .O(gate406inter8));
  nand2 gate1240(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1241(.a(s_51), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1242(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1243(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1244(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );

  xor2  gate1987(.a(N1470), .b(N973), .O(gate409inter0));
  nand2 gate1988(.a(gate409inter0), .b(s_158), .O(gate409inter1));
  and2  gate1989(.a(N1470), .b(N973), .O(gate409inter2));
  inv1  gate1990(.a(s_158), .O(gate409inter3));
  inv1  gate1991(.a(s_159), .O(gate409inter4));
  nand2 gate1992(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1993(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1994(.a(N973), .O(gate409inter7));
  inv1  gate1995(.a(N1470), .O(gate409inter8));
  nand2 gate1996(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1997(.a(s_159), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1998(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1999(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2000(.a(gate409inter12), .b(gate409inter1), .O(N1501));
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );

  xor2  gate1357(.a(N1489), .b(N1447), .O(gate414inter0));
  nand2 gate1358(.a(gate414inter0), .b(s_68), .O(gate414inter1));
  and2  gate1359(.a(N1489), .b(N1447), .O(gate414inter2));
  inv1  gate1360(.a(s_68), .O(gate414inter3));
  inv1  gate1361(.a(s_69), .O(gate414inter4));
  nand2 gate1362(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1363(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1364(.a(N1447), .O(gate414inter7));
  inv1  gate1365(.a(N1489), .O(gate414inter8));
  nand2 gate1366(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1367(.a(s_69), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1368(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1369(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1370(.a(gate414inter12), .b(gate414inter1), .O(N1517));
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );

  xor2  gate1945(.a(N1501), .b(N1471), .O(gate425inter0));
  nand2 gate1946(.a(gate425inter0), .b(s_152), .O(gate425inter1));
  and2  gate1947(.a(N1501), .b(N1471), .O(gate425inter2));
  inv1  gate1948(.a(s_152), .O(gate425inter3));
  inv1  gate1949(.a(s_153), .O(gate425inter4));
  nand2 gate1950(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1951(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1952(.a(N1471), .O(gate425inter7));
  inv1  gate1953(.a(N1501), .O(gate425inter8));
  nand2 gate1954(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1955(.a(s_153), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1956(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1957(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1958(.a(gate425inter12), .b(gate425inter1), .O(N1534));
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );

  xor2  gate1273(.a(N1531), .b(N1484), .O(gate432inter0));
  nand2 gate1274(.a(gate432inter0), .b(s_56), .O(gate432inter1));
  and2  gate1275(.a(N1531), .b(N1484), .O(gate432inter2));
  inv1  gate1276(.a(s_56), .O(gate432inter3));
  inv1  gate1277(.a(s_57), .O(gate432inter4));
  nand2 gate1278(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1279(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1280(.a(N1484), .O(gate432inter7));
  inv1  gate1281(.a(N1531), .O(gate432inter8));
  nand2 gate1282(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1283(.a(s_57), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1284(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1285(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1286(.a(gate432inter12), .b(gate432inter1), .O(N1567));
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );

  xor2  gate2323(.a(N1530), .b(N1540), .O(gate440inter0));
  nand2 gate2324(.a(gate440inter0), .b(s_206), .O(gate440inter1));
  and2  gate2325(.a(N1530), .b(N1540), .O(gate440inter2));
  inv1  gate2326(.a(s_206), .O(gate440inter3));
  inv1  gate2327(.a(s_207), .O(gate440inter4));
  nand2 gate2328(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2329(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2330(.a(N1540), .O(gate440inter7));
  inv1  gate2331(.a(N1530), .O(gate440inter8));
  nand2 gate2332(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2333(.a(s_207), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2334(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2335(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2336(.a(gate440inter12), .b(gate440inter1), .O(N1594));
inv1 gate441( .a(N1540), .O(N1595) );

  xor2  gate1329(.a(N1568), .b(N1567), .O(gate442inter0));
  nand2 gate1330(.a(gate442inter0), .b(s_64), .O(gate442inter1));
  and2  gate1331(.a(N1568), .b(N1567), .O(gate442inter2));
  inv1  gate1332(.a(s_64), .O(gate442inter3));
  inv1  gate1333(.a(s_65), .O(gate442inter4));
  nand2 gate1334(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1335(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1336(.a(N1567), .O(gate442inter7));
  inv1  gate1337(.a(N1568), .O(gate442inter8));
  nand2 gate1338(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1339(.a(s_65), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1340(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1341(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1342(.a(gate442inter12), .b(gate442inter1), .O(N1596));
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );

  xor2  gate1161(.a(N1677), .b(N1651), .O(gate480inter0));
  nand2 gate1162(.a(gate480inter0), .b(s_40), .O(gate480inter1));
  and2  gate1163(.a(N1677), .b(N1651), .O(gate480inter2));
  inv1  gate1164(.a(s_40), .O(gate480inter3));
  inv1  gate1165(.a(s_41), .O(gate480inter4));
  nand2 gate1166(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1167(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1168(.a(N1651), .O(gate480inter7));
  inv1  gate1169(.a(N1677), .O(gate480inter8));
  nand2 gate1170(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1171(.a(s_41), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1172(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1173(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1174(.a(gate480inter12), .b(gate480inter1), .O(N1710));
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );

  xor2  gate2211(.a(N1528), .b(N1685), .O(gate494inter0));
  nand2 gate2212(.a(gate494inter0), .b(s_190), .O(gate494inter1));
  and2  gate2213(.a(N1528), .b(N1685), .O(gate494inter2));
  inv1  gate2214(.a(s_190), .O(gate494inter3));
  inv1  gate2215(.a(s_191), .O(gate494inter4));
  nand2 gate2216(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2217(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2218(.a(N1685), .O(gate494inter7));
  inv1  gate2219(.a(N1528), .O(gate494inter8));
  nand2 gate2220(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2221(.a(s_191), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2222(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2223(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2224(.a(gate494inter12), .b(gate494inter1), .O(N1740));
inv1 gate495( .a(N1685), .O(N1741) );

  xor2  gate2071(.a(N1706), .b(N1671), .O(gate496inter0));
  nand2 gate2072(.a(gate496inter0), .b(s_170), .O(gate496inter1));
  and2  gate2073(.a(N1706), .b(N1671), .O(gate496inter2));
  inv1  gate2074(.a(s_170), .O(gate496inter3));
  inv1  gate2075(.a(s_171), .O(gate496inter4));
  nand2 gate2076(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2077(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2078(.a(N1671), .O(gate496inter7));
  inv1  gate2079(.a(N1706), .O(gate496inter8));
  nand2 gate2080(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2081(.a(s_171), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2082(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2083(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2084(.a(gate496inter12), .b(gate496inter1), .O(N1742));
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );

  xor2  gate2099(.a(N1711), .b(N1603), .O(gate498inter0));
  nand2 gate2100(.a(gate498inter0), .b(s_174), .O(gate498inter1));
  and2  gate2101(.a(N1711), .b(N1603), .O(gate498inter2));
  inv1  gate2102(.a(s_174), .O(gate498inter3));
  inv1  gate2103(.a(s_175), .O(gate498inter4));
  nand2 gate2104(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2105(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2106(.a(N1603), .O(gate498inter7));
  inv1  gate2107(.a(N1711), .O(gate498inter8));
  nand2 gate2108(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2109(.a(s_175), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2110(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2111(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2112(.a(gate498inter12), .b(gate498inter1), .O(N1747));

  xor2  gate1525(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate1526(.a(gate499inter0), .b(s_92), .O(gate499inter1));
  and2  gate1527(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate1528(.a(s_92), .O(gate499inter3));
  inv1  gate1529(.a(s_93), .O(gate499inter4));
  nand2 gate1530(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1531(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1532(.a(N1678), .O(gate499inter7));
  inv1  gate1533(.a(N1712), .O(gate499inter8));
  nand2 gate1534(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1535(.a(s_93), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1536(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1537(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1538(.a(gate499inter12), .b(gate499inter1), .O(N1748));
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );

  xor2  gate1007(.a(N1721), .b(N1537), .O(gate501inter0));
  nand2 gate1008(.a(gate501inter0), .b(s_18), .O(gate501inter1));
  and2  gate1009(.a(N1721), .b(N1537), .O(gate501inter2));
  inv1  gate1010(.a(s_18), .O(gate501inter3));
  inv1  gate1011(.a(s_19), .O(gate501inter4));
  nand2 gate1012(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1013(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1014(.a(N1537), .O(gate501inter7));
  inv1  gate1015(.a(N1721), .O(gate501inter8));
  nand2 gate1016(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1017(.a(s_19), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1018(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1019(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1020(.a(gate501inter12), .b(gate501inter1), .O(N1759));
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );

  xor2  gate1651(.a(N1741), .b(N1472), .O(gate507inter0));
  nand2 gate1652(.a(gate507inter0), .b(s_110), .O(gate507inter1));
  and2  gate1653(.a(N1741), .b(N1472), .O(gate507inter2));
  inv1  gate1654(.a(s_110), .O(gate507inter3));
  inv1  gate1655(.a(s_111), .O(gate507inter4));
  nand2 gate1656(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1657(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1658(.a(N1472), .O(gate507inter7));
  inv1  gate1659(.a(N1741), .O(gate507inter8));
  nand2 gate1660(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1661(.a(s_111), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1662(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1663(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1664(.a(gate507inter12), .b(gate507inter1), .O(N1769));
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );

  xor2  gate2169(.a(N1747), .b(N1710), .O(gate511inter0));
  nand2 gate2170(.a(gate511inter0), .b(s_184), .O(gate511inter1));
  and2  gate2171(.a(N1747), .b(N1710), .O(gate511inter2));
  inv1  gate2172(.a(s_184), .O(gate511inter3));
  inv1  gate2173(.a(s_185), .O(gate511inter4));
  nand2 gate2174(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2175(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2176(.a(N1710), .O(gate511inter7));
  inv1  gate2177(.a(N1747), .O(gate511inter8));
  nand2 gate2178(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2179(.a(s_185), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2180(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2181(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2182(.a(gate511inter12), .b(gate511inter1), .O(N1777));
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1679(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1680(.a(gate513inter0), .b(s_114), .O(gate513inter1));
  and2  gate1681(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1682(.a(s_114), .O(gate513inter3));
  inv1  gate1683(.a(s_115), .O(gate513inter4));
  nand2 gate1684(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1685(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1686(.a(N1731), .O(gate513inter7));
  inv1  gate1687(.a(N1682), .O(gate513inter8));
  nand2 gate1688(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1689(.a(s_115), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1690(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1691(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1692(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );

  xor2  gate1637(.a(N1683), .b(N1734), .O(gate516inter0));
  nand2 gate1638(.a(gate516inter0), .b(s_108), .O(gate516inter1));
  and2  gate1639(.a(N1683), .b(N1734), .O(gate516inter2));
  inv1  gate1640(.a(s_108), .O(gate516inter3));
  inv1  gate1641(.a(s_109), .O(gate516inter4));
  nand2 gate1642(.a(gate516inter4), .b(gate516inter3), .O(gate516inter5));
  nor2  gate1643(.a(gate516inter5), .b(gate516inter2), .O(gate516inter6));
  inv1  gate1644(.a(N1734), .O(gate516inter7));
  inv1  gate1645(.a(N1683), .O(gate516inter8));
  nand2 gate1646(.a(gate516inter8), .b(gate516inter7), .O(gate516inter9));
  nand2 gate1647(.a(s_109), .b(gate516inter3), .O(gate516inter10));
  nor2  gate1648(.a(gate516inter10), .b(gate516inter9), .O(gate516inter11));
  nor2  gate1649(.a(gate516inter11), .b(gate516inter6), .O(gate516inter12));
  nand2 gate1650(.a(gate516inter12), .b(gate516inter1), .O(N1787));
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );

  xor2  gate1917(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate1918(.a(gate520inter0), .b(s_148), .O(gate520inter1));
  and2  gate1919(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate1920(.a(s_148), .O(gate520inter3));
  inv1  gate1921(.a(s_149), .O(gate520inter4));
  nand2 gate1922(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate1923(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate1924(.a(N1751), .O(gate520inter7));
  inv1  gate1925(.a(N1155), .O(gate520inter8));
  nand2 gate1926(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate1927(.a(s_149), .b(gate520inter3), .O(gate520inter10));
  nor2  gate1928(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate1929(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate1930(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate1623(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate1624(.a(gate522inter0), .b(s_106), .O(gate522inter1));
  and2  gate1625(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate1626(.a(s_106), .O(gate522inter3));
  inv1  gate1627(.a(s_107), .O(gate522inter4));
  nand2 gate1628(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate1629(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate1630(.a(N1740), .O(gate522inter7));
  inv1  gate1631(.a(N1769), .O(gate522inter8));
  nand2 gate1632(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate1633(.a(s_107), .b(gate522inter3), .O(gate522inter10));
  nor2  gate1634(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate1635(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate1636(.a(gate522inter12), .b(gate522inter1), .O(N1798));
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );

  xor2  gate1245(.a(N1786), .b(N1615), .O(gate528inter0));
  nand2 gate1246(.a(gate528inter0), .b(s_52), .O(gate528inter1));
  and2  gate1247(.a(N1786), .b(N1615), .O(gate528inter2));
  inv1  gate1248(.a(s_52), .O(gate528inter3));
  inv1  gate1249(.a(s_53), .O(gate528inter4));
  nand2 gate1250(.a(gate528inter4), .b(gate528inter3), .O(gate528inter5));
  nor2  gate1251(.a(gate528inter5), .b(gate528inter2), .O(gate528inter6));
  inv1  gate1252(.a(N1615), .O(gate528inter7));
  inv1  gate1253(.a(N1786), .O(gate528inter8));
  nand2 gate1254(.a(gate528inter8), .b(gate528inter7), .O(gate528inter9));
  nand2 gate1255(.a(s_53), .b(gate528inter3), .O(gate528inter10));
  nor2  gate1256(.a(gate528inter10), .b(gate528inter9), .O(gate528inter11));
  nor2  gate1257(.a(gate528inter11), .b(gate528inter6), .O(gate528inter12));
  nand2 gate1258(.a(gate528inter12), .b(gate528inter1), .O(N1810));

  xor2  gate1203(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate1204(.a(gate529inter0), .b(s_46), .O(gate529inter1));
  and2  gate1205(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate1206(.a(s_46), .O(gate529inter3));
  inv1  gate1207(.a(s_47), .O(gate529inter4));
  nand2 gate1208(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate1209(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate1210(.a(N1791), .O(gate529inter7));
  inv1  gate1211(.a(N1762), .O(gate529inter8));
  nand2 gate1212(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate1213(.a(s_47), .b(gate529inter3), .O(gate529inter10));
  nor2  gate1214(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate1215(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate1216(.a(gate529inter12), .b(gate529inter1), .O(N1812));

  xor2  gate923(.a(N1764), .b(N1792), .O(gate530inter0));
  nand2 gate924(.a(gate530inter0), .b(s_6), .O(gate530inter1));
  and2  gate925(.a(N1764), .b(N1792), .O(gate530inter2));
  inv1  gate926(.a(s_6), .O(gate530inter3));
  inv1  gate927(.a(s_7), .O(gate530inter4));
  nand2 gate928(.a(gate530inter4), .b(gate530inter3), .O(gate530inter5));
  nor2  gate929(.a(gate530inter5), .b(gate530inter2), .O(gate530inter6));
  inv1  gate930(.a(N1792), .O(gate530inter7));
  inv1  gate931(.a(N1764), .O(gate530inter8));
  nand2 gate932(.a(gate530inter8), .b(gate530inter7), .O(gate530inter9));
  nand2 gate933(.a(s_7), .b(gate530inter3), .O(gate530inter10));
  nor2  gate934(.a(gate530inter10), .b(gate530inter9), .O(gate530inter11));
  nor2  gate935(.a(gate530inter11), .b(gate530inter6), .O(gate530inter12));
  nand2 gate936(.a(gate530inter12), .b(gate530inter1), .O(N1815));
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate1609(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate1610(.a(gate532inter0), .b(s_104), .O(gate532inter1));
  and2  gate1611(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate1612(.a(s_104), .O(gate532inter3));
  inv1  gate1613(.a(s_105), .O(gate532inter4));
  nand2 gate1614(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate1615(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate1616(.a(N1777), .O(gate532inter7));
  inv1  gate1617(.a(N1490), .O(gate532inter8));
  nand2 gate1618(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate1619(.a(s_105), .b(gate532inter3), .O(gate532inter10));
  nor2  gate1620(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate1621(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate1622(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );

  xor2  gate1343(.a(N1796), .b(N962), .O(gate536inter0));
  nand2 gate1344(.a(gate536inter0), .b(s_66), .O(gate536inter1));
  and2  gate1345(.a(N1796), .b(N962), .O(gate536inter2));
  inv1  gate1346(.a(s_66), .O(gate536inter3));
  inv1  gate1347(.a(s_67), .O(gate536inter4));
  nand2 gate1348(.a(gate536inter4), .b(gate536inter3), .O(gate536inter5));
  nor2  gate1349(.a(gate536inter5), .b(gate536inter2), .O(gate536inter6));
  inv1  gate1350(.a(N962), .O(gate536inter7));
  inv1  gate1351(.a(N1796), .O(gate536inter8));
  nand2 gate1352(.a(gate536inter8), .b(gate536inter7), .O(gate536inter9));
  nand2 gate1353(.a(s_67), .b(gate536inter3), .O(gate536inter10));
  nor2  gate1354(.a(gate536inter10), .b(gate536inter9), .O(gate536inter11));
  nor2  gate1355(.a(gate536inter11), .b(gate536inter6), .O(gate536inter12));
  nand2 gate1356(.a(gate536inter12), .b(gate536inter1), .O(N1825));
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );

  xor2  gate1301(.a(N1801), .b(N1772), .O(gate539inter0));
  nand2 gate1302(.a(gate539inter0), .b(s_60), .O(gate539inter1));
  and2  gate1303(.a(N1801), .b(N1772), .O(gate539inter2));
  inv1  gate1304(.a(s_60), .O(gate539inter3));
  inv1  gate1305(.a(s_61), .O(gate539inter4));
  nand2 gate1306(.a(gate539inter4), .b(gate539inter3), .O(gate539inter5));
  nor2  gate1307(.a(gate539inter5), .b(gate539inter2), .O(gate539inter6));
  inv1  gate1308(.a(N1772), .O(gate539inter7));
  inv1  gate1309(.a(N1801), .O(gate539inter8));
  nand2 gate1310(.a(gate539inter8), .b(gate539inter7), .O(gate539inter9));
  nand2 gate1311(.a(s_61), .b(gate539inter3), .O(gate539inter10));
  nor2  gate1312(.a(gate539inter10), .b(gate539inter9), .O(gate539inter11));
  nor2  gate1313(.a(gate539inter11), .b(gate539inter6), .O(gate539inter12));
  nand2 gate1314(.a(gate539inter12), .b(gate539inter1), .O(N1830));
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );

  xor2  gate1581(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate1582(.a(gate544inter0), .b(s_100), .O(gate544inter1));
  and2  gate1583(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate1584(.a(s_100), .O(gate544inter3));
  inv1  gate1585(.a(s_101), .O(gate544inter4));
  nand2 gate1586(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate1587(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate1588(.a(N1416), .O(gate544inter7));
  inv1  gate1589(.a(N1824), .O(gate544inter8));
  nand2 gate1590(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate1591(.a(s_101), .b(gate544inter3), .O(gate544inter10));
  nor2  gate1592(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate1593(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate1594(.a(gate544inter12), .b(gate544inter1), .O(N1849));
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );

  xor2  gate1791(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate1792(.a(gate546inter0), .b(s_130), .O(gate546inter1));
  and2  gate1793(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate1794(.a(s_130), .O(gate546inter3));
  inv1  gate1795(.a(s_131), .O(gate546inter4));
  nand2 gate1796(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate1797(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate1798(.a(N1319), .O(gate546inter7));
  inv1  gate1799(.a(N1827), .O(gate546inter8));
  nand2 gate1800(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate1801(.a(s_131), .b(gate546inter3), .O(gate546inter10));
  nor2  gate1802(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate1803(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate1804(.a(gate546inter12), .b(gate546inter1), .O(N1852));
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );

  xor2  gate1413(.a(N290), .b(N1798), .O(gate550inter0));
  nand2 gate1414(.a(gate550inter0), .b(s_76), .O(gate550inter1));
  and2  gate1415(.a(N290), .b(N1798), .O(gate550inter2));
  inv1  gate1416(.a(s_76), .O(gate550inter3));
  inv1  gate1417(.a(s_77), .O(gate550inter4));
  nand2 gate1418(.a(gate550inter4), .b(gate550inter3), .O(gate550inter5));
  nor2  gate1419(.a(gate550inter5), .b(gate550inter2), .O(gate550inter6));
  inv1  gate1420(.a(N1798), .O(gate550inter7));
  inv1  gate1421(.a(N290), .O(gate550inter8));
  nand2 gate1422(.a(gate550inter8), .b(gate550inter7), .O(gate550inter9));
  nand2 gate1423(.a(s_77), .b(gate550inter3), .O(gate550inter10));
  nor2  gate1424(.a(gate550inter10), .b(gate550inter9), .O(gate550inter11));
  nor2  gate1425(.a(gate550inter11), .b(gate550inter6), .O(gate550inter12));
  nand2 gate1426(.a(gate550inter12), .b(gate550inter1), .O(N1858));
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );

  xor2  gate1595(.a(N1848), .b(N1821), .O(gate557inter0));
  nand2 gate1596(.a(gate557inter0), .b(s_102), .O(gate557inter1));
  and2  gate1597(.a(N1848), .b(N1821), .O(gate557inter2));
  inv1  gate1598(.a(s_102), .O(gate557inter3));
  inv1  gate1599(.a(s_103), .O(gate557inter4));
  nand2 gate1600(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate1601(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate1602(.a(N1821), .O(gate557inter7));
  inv1  gate1603(.a(N1848), .O(gate557inter8));
  nand2 gate1604(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate1605(.a(s_103), .b(gate557inter3), .O(gate557inter10));
  nor2  gate1606(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate1607(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate1608(.a(gate557inter12), .b(gate557inter1), .O(N1878));

  xor2  gate1861(.a(N1849), .b(N1823), .O(gate558inter0));
  nand2 gate1862(.a(gate558inter0), .b(s_140), .O(gate558inter1));
  and2  gate1863(.a(N1849), .b(N1823), .O(gate558inter2));
  inv1  gate1864(.a(s_140), .O(gate558inter3));
  inv1  gate1865(.a(s_141), .O(gate558inter4));
  nand2 gate1866(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate1867(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate1868(.a(N1823), .O(gate558inter7));
  inv1  gate1869(.a(N1849), .O(gate558inter8));
  nand2 gate1870(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate1871(.a(s_141), .b(gate558inter3), .O(gate558inter10));
  nor2  gate1872(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate1873(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate1874(.a(gate558inter12), .b(gate558inter1), .O(N1879));
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );

  xor2  gate1665(.a(N1883), .b(N1717), .O(gate570inter0));
  nand2 gate1666(.a(gate570inter0), .b(s_112), .O(gate570inter1));
  and2  gate1667(.a(N1883), .b(N1717), .O(gate570inter2));
  inv1  gate1668(.a(s_112), .O(gate570inter3));
  inv1  gate1669(.a(s_113), .O(gate570inter4));
  nand2 gate1670(.a(gate570inter4), .b(gate570inter3), .O(gate570inter5));
  nor2  gate1671(.a(gate570inter5), .b(gate570inter2), .O(gate570inter6));
  inv1  gate1672(.a(N1717), .O(gate570inter7));
  inv1  gate1673(.a(N1883), .O(gate570inter8));
  nand2 gate1674(.a(gate570inter8), .b(gate570inter7), .O(gate570inter9));
  nand2 gate1675(.a(s_113), .b(gate570inter3), .O(gate570inter10));
  nor2  gate1676(.a(gate570inter10), .b(gate570inter9), .O(gate570inter11));
  nor2  gate1677(.a(gate570inter11), .b(gate570inter6), .O(gate570inter12));
  nand2 gate1678(.a(gate570inter12), .b(gate570inter1), .O(N1911));
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate2029(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate2030(.a(gate579inter0), .b(s_164), .O(gate579inter1));
  and2  gate2031(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate2032(.a(s_164), .O(gate579inter3));
  inv1  gate2033(.a(s_165), .O(gate579inter4));
  nand2 gate2034(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate2035(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate2036(.a(N1714), .O(gate579inter7));
  inv1  gate2037(.a(N1895), .O(gate579inter8));
  nand2 gate2038(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate2039(.a(s_165), .b(gate579inter3), .O(gate579inter10));
  nor2  gate2040(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate2041(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate2042(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );

  xor2  gate1147(.a(N1920), .b(N679), .O(gate586inter0));
  nand2 gate1148(.a(gate586inter0), .b(s_38), .O(gate586inter1));
  and2  gate1149(.a(N1920), .b(N679), .O(gate586inter2));
  inv1  gate1150(.a(s_38), .O(gate586inter3));
  inv1  gate1151(.a(s_39), .O(gate586inter4));
  nand2 gate1152(.a(gate586inter4), .b(gate586inter3), .O(gate586inter5));
  nor2  gate1153(.a(gate586inter5), .b(gate586inter2), .O(gate586inter6));
  inv1  gate1154(.a(N679), .O(gate586inter7));
  inv1  gate1155(.a(N1920), .O(gate586inter8));
  nand2 gate1156(.a(gate586inter8), .b(gate586inter7), .O(gate586inter9));
  nand2 gate1157(.a(s_39), .b(gate586inter3), .O(gate586inter10));
  nor2  gate1158(.a(gate586inter10), .b(gate586inter9), .O(gate586inter11));
  nor2  gate1159(.a(gate586inter11), .b(gate586inter6), .O(gate586inter12));
  nand2 gate1160(.a(gate586inter12), .b(gate586inter1), .O(N1941));
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate1175(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate1176(.a(gate596inter0), .b(s_42), .O(gate596inter1));
  and2  gate1177(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate1178(.a(s_42), .O(gate596inter3));
  inv1  gate1179(.a(s_43), .O(gate596inter4));
  nand2 gate1180(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate1181(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate1182(.a(N1930), .O(gate596inter7));
  inv1  gate1183(.a(N917), .O(gate596inter8));
  nand2 gate1184(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate1185(.a(s_43), .b(gate596inter3), .O(gate596inter10));
  nor2  gate1186(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate1187(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate1188(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );

  xor2  gate1189(.a(N1937), .b(N1944), .O(gate605inter0));
  nand2 gate1190(.a(gate605inter0), .b(s_44), .O(gate605inter1));
  and2  gate1191(.a(N1937), .b(N1944), .O(gate605inter2));
  inv1  gate1192(.a(s_44), .O(gate605inter3));
  inv1  gate1193(.a(s_45), .O(gate605inter4));
  nand2 gate1194(.a(gate605inter4), .b(gate605inter3), .O(gate605inter5));
  nor2  gate1195(.a(gate605inter5), .b(gate605inter2), .O(gate605inter6));
  inv1  gate1196(.a(N1944), .O(gate605inter7));
  inv1  gate1197(.a(N1937), .O(gate605inter8));
  nand2 gate1198(.a(gate605inter8), .b(gate605inter7), .O(gate605inter9));
  nand2 gate1199(.a(s_45), .b(gate605inter3), .O(gate605inter10));
  nor2  gate1200(.a(gate605inter10), .b(gate605inter9), .O(gate605inter11));
  nor2  gate1201(.a(gate605inter11), .b(gate605inter6), .O(gate605inter12));
  nand2 gate1202(.a(gate605inter12), .b(gate605inter1), .O(N2000));
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );

  xor2  gate1217(.a(N1351), .b(N1950), .O(gate610inter0));
  nand2 gate1218(.a(gate610inter0), .b(s_48), .O(gate610inter1));
  and2  gate1219(.a(N1351), .b(N1950), .O(gate610inter2));
  inv1  gate1220(.a(s_48), .O(gate610inter3));
  inv1  gate1221(.a(s_49), .O(gate610inter4));
  nand2 gate1222(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate1223(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate1224(.a(N1950), .O(gate610inter7));
  inv1  gate1225(.a(N1351), .O(gate610inter8));
  nand2 gate1226(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate1227(.a(s_49), .b(gate610inter3), .O(gate610inter10));
  nor2  gate1228(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate1229(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate1230(.a(gate610inter12), .b(gate610inter1), .O(N2006));
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );

  xor2  gate1385(.a(N1635), .b(N1961), .O(gate618inter0));
  nand2 gate1386(.a(gate618inter0), .b(s_72), .O(gate618inter1));
  and2  gate1387(.a(N1635), .b(N1961), .O(gate618inter2));
  inv1  gate1388(.a(s_72), .O(gate618inter3));
  inv1  gate1389(.a(s_73), .O(gate618inter4));
  nand2 gate1390(.a(gate618inter4), .b(gate618inter3), .O(gate618inter5));
  nor2  gate1391(.a(gate618inter5), .b(gate618inter2), .O(gate618inter6));
  inv1  gate1392(.a(N1961), .O(gate618inter7));
  inv1  gate1393(.a(N1635), .O(gate618inter8));
  nand2 gate1394(.a(gate618inter8), .b(gate618inter7), .O(gate618inter9));
  nand2 gate1395(.a(s_73), .b(gate618inter3), .O(gate618inter10));
  nor2  gate1396(.a(gate618inter10), .b(gate618inter9), .O(gate618inter11));
  nor2  gate1397(.a(gate618inter11), .b(gate618inter6), .O(gate618inter12));
  nand2 gate1398(.a(gate618inter12), .b(gate618inter1), .O(N2016));
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );

  xor2  gate1021(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate1022(.a(gate627inter0), .b(s_20), .O(gate627inter1));
  and2  gate1023(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate1024(.a(s_20), .O(gate627inter3));
  inv1  gate1025(.a(s_21), .O(gate627inter4));
  nand2 gate1026(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate1027(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate1028(.a(N1975), .O(gate627inter7));
  inv1  gate1029(.a(N2008), .O(gate627inter8));
  nand2 gate1030(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate1031(.a(s_21), .b(gate627inter3), .O(gate627inter10));
  nor2  gate1032(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate1033(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate1034(.a(gate627inter12), .b(gate627inter1), .O(N2026));
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );

  xor2  gate1091(.a(N2015), .b(N1571), .O(gate632inter0));
  nand2 gate1092(.a(gate632inter0), .b(s_30), .O(gate632inter1));
  and2  gate1093(.a(N2015), .b(N1571), .O(gate632inter2));
  inv1  gate1094(.a(s_30), .O(gate632inter3));
  inv1  gate1095(.a(s_31), .O(gate632inter4));
  nand2 gate1096(.a(gate632inter4), .b(gate632inter3), .O(gate632inter5));
  nor2  gate1097(.a(gate632inter5), .b(gate632inter2), .O(gate632inter6));
  inv1  gate1098(.a(N1571), .O(gate632inter7));
  inv1  gate1099(.a(N2015), .O(gate632inter8));
  nand2 gate1100(.a(gate632inter8), .b(gate632inter7), .O(gate632inter9));
  nand2 gate1101(.a(s_31), .b(gate632inter3), .O(gate632inter10));
  nor2  gate1102(.a(gate632inter10), .b(gate632inter9), .O(gate632inter11));
  nor2  gate1103(.a(gate632inter11), .b(gate632inter6), .O(gate632inter12));
  nand2 gate1104(.a(gate632inter12), .b(gate632inter1), .O(N2037));
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );

  xor2  gate1707(.a(N916), .b(N2148), .O(gate665inter0));
  nand2 gate1708(.a(gate665inter0), .b(s_118), .O(gate665inter1));
  and2  gate1709(.a(N916), .b(N2148), .O(gate665inter2));
  inv1  gate1710(.a(s_118), .O(gate665inter3));
  inv1  gate1711(.a(s_119), .O(gate665inter4));
  nand2 gate1712(.a(gate665inter4), .b(gate665inter3), .O(gate665inter5));
  nor2  gate1713(.a(gate665inter5), .b(gate665inter2), .O(gate665inter6));
  inv1  gate1714(.a(N2148), .O(gate665inter7));
  inv1  gate1715(.a(N916), .O(gate665inter8));
  nand2 gate1716(.a(gate665inter8), .b(gate665inter7), .O(gate665inter9));
  nand2 gate1717(.a(s_119), .b(gate665inter3), .O(gate665inter10));
  nor2  gate1718(.a(gate665inter10), .b(gate665inter9), .O(gate665inter11));
  nor2  gate1719(.a(gate665inter11), .b(gate665inter6), .O(gate665inter12));
  nand2 gate1720(.a(gate665inter12), .b(gate665inter1), .O(N2216));
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );

  xor2  gate1483(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate1484(.a(gate678inter0), .b(s_86), .O(gate678inter1));
  and2  gate1485(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate1486(.a(s_86), .O(gate678inter3));
  inv1  gate1487(.a(s_87), .O(gate678inter4));
  nand2 gate1488(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate1489(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate1490(.a(N1252), .O(gate678inter7));
  inv1  gate1491(.a(N2225), .O(gate678inter8));
  nand2 gate1492(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate1493(.a(s_87), .b(gate678inter3), .O(gate678inter10));
  nor2  gate1494(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate1495(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate1496(.a(gate678inter12), .b(gate678inter1), .O(N2233));
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );

  xor2  gate2337(.a(N2230), .b(N2214), .O(gate681inter0));
  nand2 gate2338(.a(gate681inter0), .b(s_208), .O(gate681inter1));
  and2  gate2339(.a(N2230), .b(N2214), .O(gate681inter2));
  inv1  gate2340(.a(s_208), .O(gate681inter3));
  inv1  gate2341(.a(s_209), .O(gate681inter4));
  nand2 gate2342(.a(gate681inter4), .b(gate681inter3), .O(gate681inter5));
  nor2  gate2343(.a(gate681inter5), .b(gate681inter2), .O(gate681inter6));
  inv1  gate2344(.a(N2214), .O(gate681inter7));
  inv1  gate2345(.a(N2230), .O(gate681inter8));
  nand2 gate2346(.a(gate681inter8), .b(gate681inter7), .O(gate681inter9));
  nand2 gate2347(.a(s_209), .b(gate681inter3), .O(gate681inter10));
  nor2  gate2348(.a(gate681inter10), .b(gate681inter9), .O(gate681inter11));
  nor2  gate2349(.a(gate681inter11), .b(gate681inter6), .O(gate681inter12));
  nand2 gate2350(.a(gate681inter12), .b(gate681inter1), .O(N2236));

  xor2  gate1259(.a(N2231), .b(N2216), .O(gate682inter0));
  nand2 gate1260(.a(gate682inter0), .b(s_54), .O(gate682inter1));
  and2  gate1261(.a(N2231), .b(N2216), .O(gate682inter2));
  inv1  gate1262(.a(s_54), .O(gate682inter3));
  inv1  gate1263(.a(s_55), .O(gate682inter4));
  nand2 gate1264(.a(gate682inter4), .b(gate682inter3), .O(gate682inter5));
  nor2  gate1265(.a(gate682inter5), .b(gate682inter2), .O(gate682inter6));
  inv1  gate1266(.a(N2216), .O(gate682inter7));
  inv1  gate1267(.a(N2231), .O(gate682inter8));
  nand2 gate1268(.a(gate682inter8), .b(gate682inter7), .O(gate682inter9));
  nand2 gate1269(.a(s_55), .b(gate682inter3), .O(gate682inter10));
  nor2  gate1270(.a(gate682inter10), .b(gate682inter9), .O(gate682inter11));
  nor2  gate1271(.a(gate682inter11), .b(gate682inter6), .O(gate682inter12));
  nand2 gate1272(.a(gate682inter12), .b(gate682inter1), .O(N2237));
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );

  xor2  gate1889(.a(N549), .b(N2576), .O(gate762inter0));
  nand2 gate1890(.a(gate762inter0), .b(s_144), .O(gate762inter1));
  and2  gate1891(.a(N549), .b(N2576), .O(gate762inter2));
  inv1  gate1892(.a(s_144), .O(gate762inter3));
  inv1  gate1893(.a(s_145), .O(gate762inter4));
  nand2 gate1894(.a(gate762inter4), .b(gate762inter3), .O(gate762inter5));
  nor2  gate1895(.a(gate762inter5), .b(gate762inter2), .O(gate762inter6));
  inv1  gate1896(.a(N2576), .O(gate762inter7));
  inv1  gate1897(.a(N549), .O(gate762inter8));
  nand2 gate1898(.a(gate762inter8), .b(gate762inter7), .O(gate762inter9));
  nand2 gate1899(.a(s_145), .b(gate762inter3), .O(gate762inter10));
  nor2  gate1900(.a(gate762inter10), .b(gate762inter9), .O(gate762inter11));
  nor2  gate1901(.a(gate762inter11), .b(gate762inter6), .O(gate762inter12));
  nand2 gate1902(.a(gate762inter12), .b(gate762inter1), .O(N2690));
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );

  xor2  gate1833(.a(N2670), .b(N343), .O(gate765inter0));
  nand2 gate1834(.a(gate765inter0), .b(s_136), .O(gate765inter1));
  and2  gate1835(.a(N2670), .b(N343), .O(gate765inter2));
  inv1  gate1836(.a(s_136), .O(gate765inter3));
  inv1  gate1837(.a(s_137), .O(gate765inter4));
  nand2 gate1838(.a(gate765inter4), .b(gate765inter3), .O(gate765inter5));
  nor2  gate1839(.a(gate765inter5), .b(gate765inter2), .O(gate765inter6));
  inv1  gate1840(.a(N343), .O(gate765inter7));
  inv1  gate1841(.a(N2670), .O(gate765inter8));
  nand2 gate1842(.a(gate765inter8), .b(gate765inter7), .O(gate765inter9));
  nand2 gate1843(.a(s_137), .b(gate765inter3), .O(gate765inter10));
  nor2  gate1844(.a(gate765inter10), .b(gate765inter9), .O(gate765inter11));
  nor2  gate1845(.a(gate765inter11), .b(gate765inter6), .O(gate765inter12));
  nand2 gate1846(.a(gate765inter12), .b(gate765inter1), .O(N2720));
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );

  xor2  gate979(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate980(.a(gate768inter0), .b(s_14), .O(gate768inter1));
  and2  gate981(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate982(.a(s_14), .O(gate768inter3));
  inv1  gate983(.a(s_15), .O(gate768inter4));
  nand2 gate984(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate985(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate986(.a(N352), .O(gate768inter7));
  inv1  gate987(.a(N2676), .O(gate768inter8));
  nand2 gate988(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate989(.a(s_15), .b(gate768inter3), .O(gate768inter10));
  nor2  gate990(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate991(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate992(.a(gate768inter12), .b(gate768inter1), .O(N2723));

  xor2  gate2281(.a(N538), .b(N2639), .O(gate769inter0));
  nand2 gate2282(.a(gate769inter0), .b(s_200), .O(gate769inter1));
  and2  gate2283(.a(N538), .b(N2639), .O(gate769inter2));
  inv1  gate2284(.a(s_200), .O(gate769inter3));
  inv1  gate2285(.a(s_201), .O(gate769inter4));
  nand2 gate2286(.a(gate769inter4), .b(gate769inter3), .O(gate769inter5));
  nor2  gate2287(.a(gate769inter5), .b(gate769inter2), .O(gate769inter6));
  inv1  gate2288(.a(N2639), .O(gate769inter7));
  inv1  gate2289(.a(N538), .O(gate769inter8));
  nand2 gate2290(.a(gate769inter8), .b(gate769inter7), .O(gate769inter9));
  nand2 gate2291(.a(s_201), .b(gate769inter3), .O(gate769inter10));
  nor2  gate2292(.a(gate769inter10), .b(gate769inter9), .O(gate769inter11));
  nor2  gate2293(.a(gate769inter11), .b(gate769inter6), .O(gate769inter12));
  nand2 gate2294(.a(gate769inter12), .b(gate769inter1), .O(N2724));
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );

  xor2  gate895(.a(N541), .b(N2648), .O(gate775inter0));
  nand2 gate896(.a(gate775inter0), .b(s_2), .O(gate775inter1));
  and2  gate897(.a(N541), .b(N2648), .O(gate775inter2));
  inv1  gate898(.a(s_2), .O(gate775inter3));
  inv1  gate899(.a(s_3), .O(gate775inter4));
  nand2 gate900(.a(gate775inter4), .b(gate775inter3), .O(gate775inter5));
  nor2  gate901(.a(gate775inter5), .b(gate775inter2), .O(gate775inter6));
  inv1  gate902(.a(N2648), .O(gate775inter7));
  inv1  gate903(.a(N541), .O(gate775inter8));
  nand2 gate904(.a(gate775inter8), .b(gate775inter7), .O(gate775inter9));
  nand2 gate905(.a(s_3), .b(gate775inter3), .O(gate775inter10));
  nor2  gate906(.a(gate775inter10), .b(gate775inter9), .O(gate775inter11));
  nor2  gate907(.a(gate775inter11), .b(gate775inter6), .O(gate775inter12));
  nand2 gate908(.a(gate775inter12), .b(gate775inter1), .O(N2730));
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );

  xor2  gate1287(.a(N547), .b(N2664), .O(gate786inter0));
  nand2 gate1288(.a(gate786inter0), .b(s_58), .O(gate786inter1));
  and2  gate1289(.a(N547), .b(N2664), .O(gate786inter2));
  inv1  gate1290(.a(s_58), .O(gate786inter3));
  inv1  gate1291(.a(s_59), .O(gate786inter4));
  nand2 gate1292(.a(gate786inter4), .b(gate786inter3), .O(gate786inter5));
  nor2  gate1293(.a(gate786inter5), .b(gate786inter2), .O(gate786inter6));
  inv1  gate1294(.a(N2664), .O(gate786inter7));
  inv1  gate1295(.a(N547), .O(gate786inter8));
  nand2 gate1296(.a(gate786inter8), .b(gate786inter7), .O(gate786inter9));
  nand2 gate1297(.a(s_59), .b(gate786inter3), .O(gate786inter10));
  nor2  gate1298(.a(gate786inter10), .b(gate786inter9), .O(gate786inter11));
  nor2  gate1299(.a(gate786inter11), .b(gate786inter6), .O(gate786inter12));
  nand2 gate1300(.a(gate786inter12), .b(gate786inter1), .O(N2741));
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );

  xor2  gate1441(.a(N2729), .b(N361), .O(gate800inter0));
  nand2 gate1442(.a(gate800inter0), .b(s_80), .O(gate800inter1));
  and2  gate1443(.a(N2729), .b(N361), .O(gate800inter2));
  inv1  gate1444(.a(s_80), .O(gate800inter3));
  inv1  gate1445(.a(s_81), .O(gate800inter4));
  nand2 gate1446(.a(gate800inter4), .b(gate800inter3), .O(gate800inter5));
  nor2  gate1447(.a(gate800inter5), .b(gate800inter2), .O(gate800inter6));
  inv1  gate1448(.a(N361), .O(gate800inter7));
  inv1  gate1449(.a(N2729), .O(gate800inter8));
  nand2 gate1450(.a(gate800inter8), .b(gate800inter7), .O(gate800inter9));
  nand2 gate1451(.a(s_81), .b(gate800inter3), .O(gate800inter10));
  nor2  gate1452(.a(gate800inter10), .b(gate800inter9), .O(gate800inter11));
  nor2  gate1453(.a(gate800inter11), .b(gate800inter6), .O(gate800inter12));
  nand2 gate1454(.a(gate800inter12), .b(gate800inter1), .O(N2759));
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );

  xor2  gate2057(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate2058(.a(gate806inter0), .b(s_168), .O(gate806inter1));
  and2  gate2059(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate2060(.a(s_168), .O(gate806inter3));
  inv1  gate2061(.a(s_169), .O(gate806inter4));
  nand2 gate2062(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate2063(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate2064(.a(N379), .O(gate806inter7));
  inv1  gate2065(.a(N2740), .O(gate806inter8));
  nand2 gate2066(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate2067(.a(s_169), .b(gate806inter3), .O(gate806inter10));
  nor2  gate2068(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate2069(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate2070(.a(gate806inter12), .b(gate806inter1), .O(N2765));
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );

  xor2  gate2267(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate2268(.a(gate813inter0), .b(s_198), .O(gate813inter1));
  and2  gate2269(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate2270(.a(s_198), .O(gate813inter3));
  inv1  gate2271(.a(s_199), .O(gate813inter4));
  nand2 gate2272(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate2273(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate2274(.a(N2726), .O(gate813inter7));
  inv1  gate2275(.a(N2758), .O(gate813inter8));
  nand2 gate2276(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate2277(.a(s_199), .b(gate813inter3), .O(gate813inter10));
  nor2  gate2278(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate2279(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate2280(.a(gate813inter12), .b(gate813inter1), .O(N2780));
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );

  xor2  gate2043(.a(N2761), .b(N2732), .O(gate816inter0));
  nand2 gate2044(.a(gate816inter0), .b(s_166), .O(gate816inter1));
  and2  gate2045(.a(N2761), .b(N2732), .O(gate816inter2));
  inv1  gate2046(.a(s_166), .O(gate816inter3));
  inv1  gate2047(.a(s_167), .O(gate816inter4));
  nand2 gate2048(.a(gate816inter4), .b(gate816inter3), .O(gate816inter5));
  nor2  gate2049(.a(gate816inter5), .b(gate816inter2), .O(gate816inter6));
  inv1  gate2050(.a(N2732), .O(gate816inter7));
  inv1  gate2051(.a(N2761), .O(gate816inter8));
  nand2 gate2052(.a(gate816inter8), .b(gate816inter7), .O(gate816inter9));
  nand2 gate2053(.a(s_167), .b(gate816inter3), .O(gate816inter10));
  nor2  gate2054(.a(gate816inter10), .b(gate816inter9), .O(gate816inter11));
  nor2  gate2055(.a(gate816inter11), .b(gate816inter6), .O(gate816inter12));
  nand2 gate2056(.a(gate816inter12), .b(gate816inter1), .O(N2783));
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );

  xor2  gate2309(.a(N2766), .b(N2741), .O(gate820inter0));
  nand2 gate2310(.a(gate820inter0), .b(s_204), .O(gate820inter1));
  and2  gate2311(.a(N2766), .b(N2741), .O(gate820inter2));
  inv1  gate2312(.a(s_204), .O(gate820inter3));
  inv1  gate2313(.a(s_205), .O(gate820inter4));
  nand2 gate2314(.a(gate820inter4), .b(gate820inter3), .O(gate820inter5));
  nor2  gate2315(.a(gate820inter5), .b(gate820inter2), .O(gate820inter6));
  inv1  gate2316(.a(N2741), .O(gate820inter7));
  inv1  gate2317(.a(N2766), .O(gate820inter8));
  nand2 gate2318(.a(gate820inter8), .b(gate820inter7), .O(gate820inter9));
  nand2 gate2319(.a(s_205), .b(gate820inter3), .O(gate820inter10));
  nor2  gate2320(.a(gate820inter10), .b(gate820inter9), .O(gate820inter11));
  nor2  gate2321(.a(gate820inter11), .b(gate820inter6), .O(gate820inter12));
  nand2 gate2322(.a(gate820inter12), .b(gate820inter1), .O(N2787));
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );

  xor2  gate2127(.a(N2827), .b(N2807), .O(gate837inter0));
  nand2 gate2128(.a(gate837inter0), .b(s_178), .O(gate837inter1));
  and2  gate2129(.a(N2827), .b(N2807), .O(gate837inter2));
  inv1  gate2130(.a(s_178), .O(gate837inter3));
  inv1  gate2131(.a(s_179), .O(gate837inter4));
  nand2 gate2132(.a(gate837inter4), .b(gate837inter3), .O(gate837inter5));
  nor2  gate2133(.a(gate837inter5), .b(gate837inter2), .O(gate837inter6));
  inv1  gate2134(.a(N2807), .O(gate837inter7));
  inv1  gate2135(.a(N2827), .O(gate837inter8));
  nand2 gate2136(.a(gate837inter8), .b(gate837inter7), .O(gate837inter9));
  nand2 gate2137(.a(s_179), .b(gate837inter3), .O(gate837inter10));
  nor2  gate2138(.a(gate837inter10), .b(gate837inter9), .O(gate837inter11));
  nor2  gate2139(.a(gate837inter11), .b(gate837inter6), .O(gate837inter12));
  nand2 gate2140(.a(gate837inter12), .b(gate837inter1), .O(N2843));
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );

  xor2  gate1497(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate1498(.a(gate839inter0), .b(s_88), .O(gate839inter1));
  and2  gate1499(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate1500(.a(s_88), .O(gate839inter3));
  inv1  gate1501(.a(s_89), .O(gate839inter4));
  nand2 gate1502(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate1503(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate1504(.a(N2812), .O(gate839inter7));
  inv1  gate1505(.a(N2076), .O(gate839inter8));
  nand2 gate1506(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate1507(.a(s_89), .b(gate839inter3), .O(gate839inter10));
  nor2  gate1508(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate1509(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate1510(.a(gate839inter12), .b(gate839inter1), .O(N2850));
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );

  xor2  gate1567(.a(N1915), .b(N2818), .O(gate841inter0));
  nand2 gate1568(.a(gate841inter0), .b(s_98), .O(gate841inter1));
  and2  gate1569(.a(N1915), .b(N2818), .O(gate841inter2));
  inv1  gate1570(.a(s_98), .O(gate841inter3));
  inv1  gate1571(.a(s_99), .O(gate841inter4));
  nand2 gate1572(.a(gate841inter4), .b(gate841inter3), .O(gate841inter5));
  nor2  gate1573(.a(gate841inter5), .b(gate841inter2), .O(gate841inter6));
  inv1  gate1574(.a(N2818), .O(gate841inter7));
  inv1  gate1575(.a(N1915), .O(gate841inter8));
  nand2 gate1576(.a(gate841inter8), .b(gate841inter7), .O(gate841inter9));
  nand2 gate1577(.a(s_99), .b(gate841inter3), .O(gate841inter10));
  nor2  gate1578(.a(gate841inter10), .b(gate841inter9), .O(gate841inter11));
  nor2  gate1579(.a(gate841inter11), .b(gate841inter6), .O(gate841inter12));
  nand2 gate1580(.a(gate841inter12), .b(gate841inter1), .O(N2852));

  xor2  gate2015(.a(N1857), .b(N2821), .O(gate842inter0));
  nand2 gate2016(.a(gate842inter0), .b(s_162), .O(gate842inter1));
  and2  gate2017(.a(N1857), .b(N2821), .O(gate842inter2));
  inv1  gate2018(.a(s_162), .O(gate842inter3));
  inv1  gate2019(.a(s_163), .O(gate842inter4));
  nand2 gate2020(.a(gate842inter4), .b(gate842inter3), .O(gate842inter5));
  nor2  gate2021(.a(gate842inter5), .b(gate842inter2), .O(gate842inter6));
  inv1  gate2022(.a(N2821), .O(gate842inter7));
  inv1  gate2023(.a(N1857), .O(gate842inter8));
  nand2 gate2024(.a(gate842inter8), .b(gate842inter7), .O(gate842inter9));
  nand2 gate2025(.a(s_163), .b(gate842inter3), .O(gate842inter10));
  nor2  gate2026(.a(gate842inter10), .b(gate842inter9), .O(gate842inter11));
  nor2  gate2027(.a(gate842inter11), .b(gate842inter6), .O(gate842inter12));
  nand2 gate2028(.a(gate842inter12), .b(gate842inter1), .O(N2853));
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );

  xor2  gate2295(.a(N2857), .b(N2052), .O(gate851inter0));
  nand2 gate2296(.a(gate851inter0), .b(s_202), .O(gate851inter1));
  and2  gate2297(.a(N2857), .b(N2052), .O(gate851inter2));
  inv1  gate2298(.a(s_202), .O(gate851inter3));
  inv1  gate2299(.a(s_203), .O(gate851inter4));
  nand2 gate2300(.a(gate851inter4), .b(gate851inter3), .O(gate851inter5));
  nor2  gate2301(.a(gate851inter5), .b(gate851inter2), .O(gate851inter6));
  inv1  gate2302(.a(N2052), .O(gate851inter7));
  inv1  gate2303(.a(N2857), .O(gate851inter8));
  nand2 gate2304(.a(gate851inter8), .b(gate851inter7), .O(gate851inter9));
  nand2 gate2305(.a(s_203), .b(gate851inter3), .O(gate851inter10));
  nor2  gate2306(.a(gate851inter10), .b(gate851inter9), .O(gate851inter11));
  nor2  gate2307(.a(gate851inter11), .b(gate851inter6), .O(gate851inter12));
  nand2 gate2308(.a(gate851inter12), .b(gate851inter1), .O(N2866));
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );

  xor2  gate1875(.a(N2861), .b(N1902), .O(gate855inter0));
  nand2 gate1876(.a(gate855inter0), .b(s_142), .O(gate855inter1));
  and2  gate1877(.a(N2861), .b(N1902), .O(gate855inter2));
  inv1  gate1878(.a(s_142), .O(gate855inter3));
  inv1  gate1879(.a(s_143), .O(gate855inter4));
  nand2 gate1880(.a(gate855inter4), .b(gate855inter3), .O(gate855inter5));
  nor2  gate1881(.a(gate855inter5), .b(gate855inter2), .O(gate855inter6));
  inv1  gate1882(.a(N1902), .O(gate855inter7));
  inv1  gate1883(.a(N2861), .O(gate855inter8));
  nand2 gate1884(.a(gate855inter8), .b(gate855inter7), .O(gate855inter9));
  nand2 gate1885(.a(s_143), .b(gate855inter3), .O(gate855inter10));
  nor2  gate1886(.a(gate855inter10), .b(gate855inter9), .O(gate855inter11));
  nor2  gate1887(.a(gate855inter11), .b(gate855inter6), .O(gate855inter12));
  nand2 gate1888(.a(gate855inter12), .b(gate855inter1), .O(N2870));

  xor2  gate1469(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1470(.a(gate856inter0), .b(s_84), .O(gate856inter1));
  and2  gate1471(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1472(.a(s_84), .O(gate856inter3));
  inv1  gate1473(.a(s_85), .O(gate856inter4));
  nand2 gate1474(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1475(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1476(.a(N2843), .O(gate856inter7));
  inv1  gate1477(.a(N886), .O(gate856inter8));
  nand2 gate1478(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1479(.a(s_85), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1480(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1481(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1482(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );

  xor2  gate1133(.a(N2872), .b(N682), .O(gate866inter0));
  nand2 gate1134(.a(gate866inter0), .b(s_36), .O(gate866inter1));
  and2  gate1135(.a(N2872), .b(N682), .O(gate866inter2));
  inv1  gate1136(.a(s_36), .O(gate866inter3));
  inv1  gate1137(.a(s_37), .O(gate866inter4));
  nand2 gate1138(.a(gate866inter4), .b(gate866inter3), .O(gate866inter5));
  nor2  gate1139(.a(gate866inter5), .b(gate866inter2), .O(gate866inter6));
  inv1  gate1140(.a(N682), .O(gate866inter7));
  inv1  gate1141(.a(N2872), .O(gate866inter8));
  nand2 gate1142(.a(gate866inter8), .b(gate866inter7), .O(gate866inter9));
  nand2 gate1143(.a(s_37), .b(gate866inter3), .O(gate866inter10));
  nor2  gate1144(.a(gate866inter10), .b(gate866inter9), .O(gate866inter11));
  nor2  gate1145(.a(gate866inter11), .b(gate866inter6), .O(gate866inter12));
  nand2 gate1146(.a(gate866inter12), .b(gate866inter1), .O(N2881));
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );

  xor2  gate2085(.a(N2863), .b(N2875), .O(gate868inter0));
  nand2 gate2086(.a(gate868inter0), .b(s_172), .O(gate868inter1));
  and2  gate2087(.a(N2863), .b(N2875), .O(gate868inter2));
  inv1  gate2088(.a(s_172), .O(gate868inter3));
  inv1  gate2089(.a(s_173), .O(gate868inter4));
  nand2 gate2090(.a(gate868inter4), .b(gate868inter3), .O(gate868inter5));
  nor2  gate2091(.a(gate868inter5), .b(gate868inter2), .O(gate868inter6));
  inv1  gate2092(.a(N2875), .O(gate868inter7));
  inv1  gate2093(.a(N2863), .O(gate868inter8));
  nand2 gate2094(.a(gate868inter8), .b(gate868inter7), .O(gate868inter9));
  nand2 gate2095(.a(s_173), .b(gate868inter3), .O(gate868inter10));
  nor2  gate2096(.a(gate868inter10), .b(gate868inter9), .O(gate868inter11));
  nor2  gate2097(.a(gate868inter11), .b(gate868inter6), .O(gate868inter12));
  nand2 gate2098(.a(gate868inter12), .b(gate868inter1), .O(N2883));
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate1721(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate1722(.a(gate874inter0), .b(s_120), .O(gate874inter1));
  and2  gate1723(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate1724(.a(s_120), .O(gate874inter3));
  inv1  gate1725(.a(s_121), .O(gate874inter4));
  nand2 gate1726(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate1727(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate1728(.a(N2871), .O(gate874inter7));
  inv1  gate1729(.a(N2881), .O(gate874inter8));
  nand2 gate1730(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate1731(.a(s_121), .b(gate874inter3), .O(gate874inter10));
  nor2  gate1732(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate1733(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate1734(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule