module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2185(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2186(.a(gate9inter0), .b(s_234), .O(gate9inter1));
  and2  gate2187(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2188(.a(s_234), .O(gate9inter3));
  inv1  gate2189(.a(s_235), .O(gate9inter4));
  nand2 gate2190(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2191(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2192(.a(G1), .O(gate9inter7));
  inv1  gate2193(.a(G2), .O(gate9inter8));
  nand2 gate2194(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2195(.a(s_235), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2196(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2197(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2198(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2577(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2578(.a(gate13inter0), .b(s_290), .O(gate13inter1));
  and2  gate2579(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2580(.a(s_290), .O(gate13inter3));
  inv1  gate2581(.a(s_291), .O(gate13inter4));
  nand2 gate2582(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2583(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2584(.a(G9), .O(gate13inter7));
  inv1  gate2585(.a(G10), .O(gate13inter8));
  nand2 gate2586(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2587(.a(s_291), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2588(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2589(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2590(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate2227(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2228(.a(gate14inter0), .b(s_240), .O(gate14inter1));
  and2  gate2229(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2230(.a(s_240), .O(gate14inter3));
  inv1  gate2231(.a(s_241), .O(gate14inter4));
  nand2 gate2232(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2233(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2234(.a(G11), .O(gate14inter7));
  inv1  gate2235(.a(G12), .O(gate14inter8));
  nand2 gate2236(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2237(.a(s_241), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2238(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2239(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2240(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1541(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1542(.a(gate18inter0), .b(s_142), .O(gate18inter1));
  and2  gate1543(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1544(.a(s_142), .O(gate18inter3));
  inv1  gate1545(.a(s_143), .O(gate18inter4));
  nand2 gate1546(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1547(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1548(.a(G19), .O(gate18inter7));
  inv1  gate1549(.a(G20), .O(gate18inter8));
  nand2 gate1550(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1551(.a(s_143), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1552(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1553(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1554(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate701(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate702(.a(gate20inter0), .b(s_22), .O(gate20inter1));
  and2  gate703(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate704(.a(s_22), .O(gate20inter3));
  inv1  gate705(.a(s_23), .O(gate20inter4));
  nand2 gate706(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate707(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate708(.a(G23), .O(gate20inter7));
  inv1  gate709(.a(G24), .O(gate20inter8));
  nand2 gate710(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate711(.a(s_23), .b(gate20inter3), .O(gate20inter10));
  nor2  gate712(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate713(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate714(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2675(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2676(.a(gate21inter0), .b(s_304), .O(gate21inter1));
  and2  gate2677(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2678(.a(s_304), .O(gate21inter3));
  inv1  gate2679(.a(s_305), .O(gate21inter4));
  nand2 gate2680(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2681(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2682(.a(G25), .O(gate21inter7));
  inv1  gate2683(.a(G26), .O(gate21inter8));
  nand2 gate2684(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2685(.a(s_305), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2686(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2687(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2688(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1345(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1346(.a(gate22inter0), .b(s_114), .O(gate22inter1));
  and2  gate1347(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1348(.a(s_114), .O(gate22inter3));
  inv1  gate1349(.a(s_115), .O(gate22inter4));
  nand2 gate1350(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1351(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1352(.a(G27), .O(gate22inter7));
  inv1  gate1353(.a(G28), .O(gate22inter8));
  nand2 gate1354(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1355(.a(s_115), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1356(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1357(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1358(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1093(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1094(.a(gate25inter0), .b(s_78), .O(gate25inter1));
  and2  gate1095(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1096(.a(s_78), .O(gate25inter3));
  inv1  gate1097(.a(s_79), .O(gate25inter4));
  nand2 gate1098(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1099(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1100(.a(G1), .O(gate25inter7));
  inv1  gate1101(.a(G5), .O(gate25inter8));
  nand2 gate1102(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1103(.a(s_79), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1104(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1105(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1106(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate2871(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2872(.a(gate26inter0), .b(s_332), .O(gate26inter1));
  and2  gate2873(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2874(.a(s_332), .O(gate26inter3));
  inv1  gate2875(.a(s_333), .O(gate26inter4));
  nand2 gate2876(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2877(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2878(.a(G9), .O(gate26inter7));
  inv1  gate2879(.a(G13), .O(gate26inter8));
  nand2 gate2880(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2881(.a(s_333), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2882(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2883(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2884(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2843(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2844(.a(gate33inter0), .b(s_328), .O(gate33inter1));
  and2  gate2845(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2846(.a(s_328), .O(gate33inter3));
  inv1  gate2847(.a(s_329), .O(gate33inter4));
  nand2 gate2848(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2849(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2850(.a(G17), .O(gate33inter7));
  inv1  gate2851(.a(G21), .O(gate33inter8));
  nand2 gate2852(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2853(.a(s_329), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2854(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2855(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2856(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1807(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1808(.a(gate34inter0), .b(s_180), .O(gate34inter1));
  and2  gate1809(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1810(.a(s_180), .O(gate34inter3));
  inv1  gate1811(.a(s_181), .O(gate34inter4));
  nand2 gate1812(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1813(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1814(.a(G25), .O(gate34inter7));
  inv1  gate1815(.a(G29), .O(gate34inter8));
  nand2 gate1816(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1817(.a(s_181), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1818(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1819(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1820(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1387(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1388(.a(gate35inter0), .b(s_120), .O(gate35inter1));
  and2  gate1389(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1390(.a(s_120), .O(gate35inter3));
  inv1  gate1391(.a(s_121), .O(gate35inter4));
  nand2 gate1392(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1393(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1394(.a(G18), .O(gate35inter7));
  inv1  gate1395(.a(G22), .O(gate35inter8));
  nand2 gate1396(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1397(.a(s_121), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1398(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1399(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1400(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate603(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate604(.a(gate37inter0), .b(s_8), .O(gate37inter1));
  and2  gate605(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate606(.a(s_8), .O(gate37inter3));
  inv1  gate607(.a(s_9), .O(gate37inter4));
  nand2 gate608(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate609(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate610(.a(G19), .O(gate37inter7));
  inv1  gate611(.a(G23), .O(gate37inter8));
  nand2 gate612(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate613(.a(s_9), .b(gate37inter3), .O(gate37inter10));
  nor2  gate614(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate615(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate616(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate3081(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate3082(.a(gate39inter0), .b(s_362), .O(gate39inter1));
  and2  gate3083(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate3084(.a(s_362), .O(gate39inter3));
  inv1  gate3085(.a(s_363), .O(gate39inter4));
  nand2 gate3086(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate3087(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate3088(.a(G20), .O(gate39inter7));
  inv1  gate3089(.a(G24), .O(gate39inter8));
  nand2 gate3090(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate3091(.a(s_363), .b(gate39inter3), .O(gate39inter10));
  nor2  gate3092(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate3093(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate3094(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1709(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1710(.a(gate40inter0), .b(s_166), .O(gate40inter1));
  and2  gate1711(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1712(.a(s_166), .O(gate40inter3));
  inv1  gate1713(.a(s_167), .O(gate40inter4));
  nand2 gate1714(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1715(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1716(.a(G28), .O(gate40inter7));
  inv1  gate1717(.a(G32), .O(gate40inter8));
  nand2 gate1718(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1719(.a(s_167), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1720(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1721(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1722(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2591(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2592(.a(gate41inter0), .b(s_292), .O(gate41inter1));
  and2  gate2593(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2594(.a(s_292), .O(gate41inter3));
  inv1  gate2595(.a(s_293), .O(gate41inter4));
  nand2 gate2596(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2597(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2598(.a(G1), .O(gate41inter7));
  inv1  gate2599(.a(G266), .O(gate41inter8));
  nand2 gate2600(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2601(.a(s_293), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2602(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2603(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2604(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate3095(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate3096(.a(gate42inter0), .b(s_364), .O(gate42inter1));
  and2  gate3097(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate3098(.a(s_364), .O(gate42inter3));
  inv1  gate3099(.a(s_365), .O(gate42inter4));
  nand2 gate3100(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate3101(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate3102(.a(G2), .O(gate42inter7));
  inv1  gate3103(.a(G266), .O(gate42inter8));
  nand2 gate3104(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate3105(.a(s_365), .b(gate42inter3), .O(gate42inter10));
  nor2  gate3106(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate3107(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate3108(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1485(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1486(.a(gate43inter0), .b(s_134), .O(gate43inter1));
  and2  gate1487(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1488(.a(s_134), .O(gate43inter3));
  inv1  gate1489(.a(s_135), .O(gate43inter4));
  nand2 gate1490(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1491(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1492(.a(G3), .O(gate43inter7));
  inv1  gate1493(.a(G269), .O(gate43inter8));
  nand2 gate1494(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1495(.a(s_135), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1496(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1497(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1498(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1863(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1864(.a(gate47inter0), .b(s_188), .O(gate47inter1));
  and2  gate1865(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1866(.a(s_188), .O(gate47inter3));
  inv1  gate1867(.a(s_189), .O(gate47inter4));
  nand2 gate1868(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1869(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1870(.a(G7), .O(gate47inter7));
  inv1  gate1871(.a(G275), .O(gate47inter8));
  nand2 gate1872(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1873(.a(s_189), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1874(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1875(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1876(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2983(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2984(.a(gate48inter0), .b(s_348), .O(gate48inter1));
  and2  gate2985(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2986(.a(s_348), .O(gate48inter3));
  inv1  gate2987(.a(s_349), .O(gate48inter4));
  nand2 gate2988(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2989(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2990(.a(G8), .O(gate48inter7));
  inv1  gate2991(.a(G275), .O(gate48inter8));
  nand2 gate2992(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2993(.a(s_349), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2994(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2995(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2996(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1653(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1654(.a(gate50inter0), .b(s_158), .O(gate50inter1));
  and2  gate1655(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1656(.a(s_158), .O(gate50inter3));
  inv1  gate1657(.a(s_159), .O(gate50inter4));
  nand2 gate1658(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1659(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1660(.a(G10), .O(gate50inter7));
  inv1  gate1661(.a(G278), .O(gate50inter8));
  nand2 gate1662(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1663(.a(s_159), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1664(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1665(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1666(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1835(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1836(.a(gate52inter0), .b(s_184), .O(gate52inter1));
  and2  gate1837(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1838(.a(s_184), .O(gate52inter3));
  inv1  gate1839(.a(s_185), .O(gate52inter4));
  nand2 gate1840(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1841(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1842(.a(G12), .O(gate52inter7));
  inv1  gate1843(.a(G281), .O(gate52inter8));
  nand2 gate1844(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1845(.a(s_185), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1846(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1847(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1848(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2437(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2438(.a(gate55inter0), .b(s_270), .O(gate55inter1));
  and2  gate2439(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2440(.a(s_270), .O(gate55inter3));
  inv1  gate2441(.a(s_271), .O(gate55inter4));
  nand2 gate2442(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2443(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2444(.a(G15), .O(gate55inter7));
  inv1  gate2445(.a(G287), .O(gate55inter8));
  nand2 gate2446(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2447(.a(s_271), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2448(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2449(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2450(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2395(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2396(.a(gate56inter0), .b(s_264), .O(gate56inter1));
  and2  gate2397(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2398(.a(s_264), .O(gate56inter3));
  inv1  gate2399(.a(s_265), .O(gate56inter4));
  nand2 gate2400(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2401(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2402(.a(G16), .O(gate56inter7));
  inv1  gate2403(.a(G287), .O(gate56inter8));
  nand2 gate2404(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2405(.a(s_265), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2406(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2407(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2408(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1639(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1640(.a(gate58inter0), .b(s_156), .O(gate58inter1));
  and2  gate1641(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1642(.a(s_156), .O(gate58inter3));
  inv1  gate1643(.a(s_157), .O(gate58inter4));
  nand2 gate1644(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1645(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1646(.a(G18), .O(gate58inter7));
  inv1  gate1647(.a(G290), .O(gate58inter8));
  nand2 gate1648(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1649(.a(s_157), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1650(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1651(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1652(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2129(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2130(.a(gate60inter0), .b(s_226), .O(gate60inter1));
  and2  gate2131(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2132(.a(s_226), .O(gate60inter3));
  inv1  gate2133(.a(s_227), .O(gate60inter4));
  nand2 gate2134(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2135(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2136(.a(G20), .O(gate60inter7));
  inv1  gate2137(.a(G293), .O(gate60inter8));
  nand2 gate2138(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2139(.a(s_227), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2140(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2141(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2142(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2115(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2116(.a(gate62inter0), .b(s_224), .O(gate62inter1));
  and2  gate2117(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2118(.a(s_224), .O(gate62inter3));
  inv1  gate2119(.a(s_225), .O(gate62inter4));
  nand2 gate2120(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2121(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2122(.a(G22), .O(gate62inter7));
  inv1  gate2123(.a(G296), .O(gate62inter8));
  nand2 gate2124(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2125(.a(s_225), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2126(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2127(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2128(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate3025(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate3026(.a(gate64inter0), .b(s_354), .O(gate64inter1));
  and2  gate3027(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate3028(.a(s_354), .O(gate64inter3));
  inv1  gate3029(.a(s_355), .O(gate64inter4));
  nand2 gate3030(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate3031(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate3032(.a(G24), .O(gate64inter7));
  inv1  gate3033(.a(G299), .O(gate64inter8));
  nand2 gate3034(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate3035(.a(s_355), .b(gate64inter3), .O(gate64inter10));
  nor2  gate3036(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate3037(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate3038(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate575(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate576(.a(gate65inter0), .b(s_4), .O(gate65inter1));
  and2  gate577(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate578(.a(s_4), .O(gate65inter3));
  inv1  gate579(.a(s_5), .O(gate65inter4));
  nand2 gate580(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate581(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate582(.a(G25), .O(gate65inter7));
  inv1  gate583(.a(G302), .O(gate65inter8));
  nand2 gate584(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate585(.a(s_5), .b(gate65inter3), .O(gate65inter10));
  nor2  gate586(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate587(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate588(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2927(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2928(.a(gate70inter0), .b(s_340), .O(gate70inter1));
  and2  gate2929(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2930(.a(s_340), .O(gate70inter3));
  inv1  gate2931(.a(s_341), .O(gate70inter4));
  nand2 gate2932(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2933(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2934(.a(G30), .O(gate70inter7));
  inv1  gate2935(.a(G308), .O(gate70inter8));
  nand2 gate2936(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2937(.a(s_341), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2938(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2939(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2940(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate2409(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2410(.a(gate71inter0), .b(s_266), .O(gate71inter1));
  and2  gate2411(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2412(.a(s_266), .O(gate71inter3));
  inv1  gate2413(.a(s_267), .O(gate71inter4));
  nand2 gate2414(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2415(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2416(.a(G31), .O(gate71inter7));
  inv1  gate2417(.a(G311), .O(gate71inter8));
  nand2 gate2418(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2419(.a(s_267), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2420(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2421(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2422(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate561(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate562(.a(gate73inter0), .b(s_2), .O(gate73inter1));
  and2  gate563(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate564(.a(s_2), .O(gate73inter3));
  inv1  gate565(.a(s_3), .O(gate73inter4));
  nand2 gate566(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate567(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate568(.a(G1), .O(gate73inter7));
  inv1  gate569(.a(G314), .O(gate73inter8));
  nand2 gate570(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate571(.a(s_3), .b(gate73inter3), .O(gate73inter10));
  nor2  gate572(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate573(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate574(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2731(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2732(.a(gate77inter0), .b(s_312), .O(gate77inter1));
  and2  gate2733(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2734(.a(s_312), .O(gate77inter3));
  inv1  gate2735(.a(s_313), .O(gate77inter4));
  nand2 gate2736(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2737(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2738(.a(G2), .O(gate77inter7));
  inv1  gate2739(.a(G320), .O(gate77inter8));
  nand2 gate2740(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2741(.a(s_313), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2742(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2743(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2744(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate869(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate870(.a(gate81inter0), .b(s_46), .O(gate81inter1));
  and2  gate871(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate872(.a(s_46), .O(gate81inter3));
  inv1  gate873(.a(s_47), .O(gate81inter4));
  nand2 gate874(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate875(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate876(.a(G3), .O(gate81inter7));
  inv1  gate877(.a(G326), .O(gate81inter8));
  nand2 gate878(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate879(.a(s_47), .b(gate81inter3), .O(gate81inter10));
  nor2  gate880(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate881(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate882(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate925(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate926(.a(gate82inter0), .b(s_54), .O(gate82inter1));
  and2  gate927(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate928(.a(s_54), .O(gate82inter3));
  inv1  gate929(.a(s_55), .O(gate82inter4));
  nand2 gate930(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate931(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate932(.a(G7), .O(gate82inter7));
  inv1  gate933(.a(G326), .O(gate82inter8));
  nand2 gate934(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate935(.a(s_55), .b(gate82inter3), .O(gate82inter10));
  nor2  gate936(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate937(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate938(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate897(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate898(.a(gate87inter0), .b(s_50), .O(gate87inter1));
  and2  gate899(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate900(.a(s_50), .O(gate87inter3));
  inv1  gate901(.a(s_51), .O(gate87inter4));
  nand2 gate902(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate903(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate904(.a(G12), .O(gate87inter7));
  inv1  gate905(.a(G335), .O(gate87inter8));
  nand2 gate906(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate907(.a(s_51), .b(gate87inter3), .O(gate87inter10));
  nor2  gate908(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate909(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate910(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate2913(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2914(.a(gate88inter0), .b(s_338), .O(gate88inter1));
  and2  gate2915(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2916(.a(s_338), .O(gate88inter3));
  inv1  gate2917(.a(s_339), .O(gate88inter4));
  nand2 gate2918(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2919(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2920(.a(G16), .O(gate88inter7));
  inv1  gate2921(.a(G335), .O(gate88inter8));
  nand2 gate2922(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2923(.a(s_339), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2924(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2925(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2926(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2661(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2662(.a(gate89inter0), .b(s_302), .O(gate89inter1));
  and2  gate2663(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2664(.a(s_302), .O(gate89inter3));
  inv1  gate2665(.a(s_303), .O(gate89inter4));
  nand2 gate2666(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2667(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2668(.a(G17), .O(gate89inter7));
  inv1  gate2669(.a(G338), .O(gate89inter8));
  nand2 gate2670(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2671(.a(s_303), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2672(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2673(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2674(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1933(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1934(.a(gate90inter0), .b(s_198), .O(gate90inter1));
  and2  gate1935(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1936(.a(s_198), .O(gate90inter3));
  inv1  gate1937(.a(s_199), .O(gate90inter4));
  nand2 gate1938(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1939(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1940(.a(G21), .O(gate90inter7));
  inv1  gate1941(.a(G338), .O(gate90inter8));
  nand2 gate1942(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1943(.a(s_199), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1944(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1945(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1946(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate547(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate548(.a(gate92inter0), .b(s_0), .O(gate92inter1));
  and2  gate549(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate550(.a(s_0), .O(gate92inter3));
  inv1  gate551(.a(s_1), .O(gate92inter4));
  nand2 gate552(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate553(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate554(.a(G29), .O(gate92inter7));
  inv1  gate555(.a(G341), .O(gate92inter8));
  nand2 gate556(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate557(.a(s_1), .b(gate92inter3), .O(gate92inter10));
  nor2  gate558(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate559(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate560(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate729(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate730(.a(gate93inter0), .b(s_26), .O(gate93inter1));
  and2  gate731(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate732(.a(s_26), .O(gate93inter3));
  inv1  gate733(.a(s_27), .O(gate93inter4));
  nand2 gate734(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate735(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate736(.a(G18), .O(gate93inter7));
  inv1  gate737(.a(G344), .O(gate93inter8));
  nand2 gate738(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate739(.a(s_27), .b(gate93inter3), .O(gate93inter10));
  nor2  gate740(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate741(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate742(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1919(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1920(.a(gate94inter0), .b(s_196), .O(gate94inter1));
  and2  gate1921(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1922(.a(s_196), .O(gate94inter3));
  inv1  gate1923(.a(s_197), .O(gate94inter4));
  nand2 gate1924(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1925(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1926(.a(G22), .O(gate94inter7));
  inv1  gate1927(.a(G344), .O(gate94inter8));
  nand2 gate1928(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1929(.a(s_197), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1930(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1931(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1932(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1471(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1472(.a(gate95inter0), .b(s_132), .O(gate95inter1));
  and2  gate1473(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1474(.a(s_132), .O(gate95inter3));
  inv1  gate1475(.a(s_133), .O(gate95inter4));
  nand2 gate1476(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1477(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1478(.a(G26), .O(gate95inter7));
  inv1  gate1479(.a(G347), .O(gate95inter8));
  nand2 gate1480(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1481(.a(s_133), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1482(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1483(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1484(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate3067(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate3068(.a(gate98inter0), .b(s_360), .O(gate98inter1));
  and2  gate3069(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate3070(.a(s_360), .O(gate98inter3));
  inv1  gate3071(.a(s_361), .O(gate98inter4));
  nand2 gate3072(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate3073(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate3074(.a(G23), .O(gate98inter7));
  inv1  gate3075(.a(G350), .O(gate98inter8));
  nand2 gate3076(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate3077(.a(s_361), .b(gate98inter3), .O(gate98inter10));
  nor2  gate3078(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate3079(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate3080(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1065(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1066(.a(gate99inter0), .b(s_74), .O(gate99inter1));
  and2  gate1067(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1068(.a(s_74), .O(gate99inter3));
  inv1  gate1069(.a(s_75), .O(gate99inter4));
  nand2 gate1070(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1071(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1072(.a(G27), .O(gate99inter7));
  inv1  gate1073(.a(G353), .O(gate99inter8));
  nand2 gate1074(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1075(.a(s_75), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1076(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1077(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1078(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1177(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1178(.a(gate102inter0), .b(s_90), .O(gate102inter1));
  and2  gate1179(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1180(.a(s_90), .O(gate102inter3));
  inv1  gate1181(.a(s_91), .O(gate102inter4));
  nand2 gate1182(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1183(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1184(.a(G24), .O(gate102inter7));
  inv1  gate1185(.a(G356), .O(gate102inter8));
  nand2 gate1186(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1187(.a(s_91), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1188(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1189(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1190(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1359(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1360(.a(gate103inter0), .b(s_116), .O(gate103inter1));
  and2  gate1361(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1362(.a(s_116), .O(gate103inter3));
  inv1  gate1363(.a(s_117), .O(gate103inter4));
  nand2 gate1364(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1365(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1366(.a(G28), .O(gate103inter7));
  inv1  gate1367(.a(G359), .O(gate103inter8));
  nand2 gate1368(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1369(.a(s_117), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1370(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1371(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1372(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate645(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate646(.a(gate108inter0), .b(s_14), .O(gate108inter1));
  and2  gate647(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate648(.a(s_14), .O(gate108inter3));
  inv1  gate649(.a(s_15), .O(gate108inter4));
  nand2 gate650(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate651(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate652(.a(G368), .O(gate108inter7));
  inv1  gate653(.a(G369), .O(gate108inter8));
  nand2 gate654(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate655(.a(s_15), .b(gate108inter3), .O(gate108inter10));
  nor2  gate656(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate657(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate658(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate939(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate940(.a(gate113inter0), .b(s_56), .O(gate113inter1));
  and2  gate941(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate942(.a(s_56), .O(gate113inter3));
  inv1  gate943(.a(s_57), .O(gate113inter4));
  nand2 gate944(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate945(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate946(.a(G378), .O(gate113inter7));
  inv1  gate947(.a(G379), .O(gate113inter8));
  nand2 gate948(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate949(.a(s_57), .b(gate113inter3), .O(gate113inter10));
  nor2  gate950(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate951(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate952(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate2171(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2172(.a(gate114inter0), .b(s_232), .O(gate114inter1));
  and2  gate2173(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2174(.a(s_232), .O(gate114inter3));
  inv1  gate2175(.a(s_233), .O(gate114inter4));
  nand2 gate2176(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2177(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2178(.a(G380), .O(gate114inter7));
  inv1  gate2179(.a(G381), .O(gate114inter8));
  nand2 gate2180(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2181(.a(s_233), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2182(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2183(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2184(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1555(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1556(.a(gate116inter0), .b(s_144), .O(gate116inter1));
  and2  gate1557(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1558(.a(s_144), .O(gate116inter3));
  inv1  gate1559(.a(s_145), .O(gate116inter4));
  nand2 gate1560(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1561(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1562(.a(G384), .O(gate116inter7));
  inv1  gate1563(.a(G385), .O(gate116inter8));
  nand2 gate1564(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1565(.a(s_145), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1566(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1567(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1568(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2899(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2900(.a(gate120inter0), .b(s_336), .O(gate120inter1));
  and2  gate2901(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2902(.a(s_336), .O(gate120inter3));
  inv1  gate2903(.a(s_337), .O(gate120inter4));
  nand2 gate2904(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2905(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2906(.a(G392), .O(gate120inter7));
  inv1  gate2907(.a(G393), .O(gate120inter8));
  nand2 gate2908(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2909(.a(s_337), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2910(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2911(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2912(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1779(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1780(.a(gate124inter0), .b(s_176), .O(gate124inter1));
  and2  gate1781(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1782(.a(s_176), .O(gate124inter3));
  inv1  gate1783(.a(s_177), .O(gate124inter4));
  nand2 gate1784(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1785(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1786(.a(G400), .O(gate124inter7));
  inv1  gate1787(.a(G401), .O(gate124inter8));
  nand2 gate1788(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1789(.a(s_177), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1790(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1791(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1792(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate799(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate800(.a(gate125inter0), .b(s_36), .O(gate125inter1));
  and2  gate801(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate802(.a(s_36), .O(gate125inter3));
  inv1  gate803(.a(s_37), .O(gate125inter4));
  nand2 gate804(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate805(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate806(.a(G402), .O(gate125inter7));
  inv1  gate807(.a(G403), .O(gate125inter8));
  nand2 gate808(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate809(.a(s_37), .b(gate125inter3), .O(gate125inter10));
  nor2  gate810(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate811(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate812(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate2773(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2774(.a(gate126inter0), .b(s_318), .O(gate126inter1));
  and2  gate2775(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2776(.a(s_318), .O(gate126inter3));
  inv1  gate2777(.a(s_319), .O(gate126inter4));
  nand2 gate2778(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2779(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2780(.a(G404), .O(gate126inter7));
  inv1  gate2781(.a(G405), .O(gate126inter8));
  nand2 gate2782(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2783(.a(s_319), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2784(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2785(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2786(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1303(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1304(.a(gate127inter0), .b(s_108), .O(gate127inter1));
  and2  gate1305(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1306(.a(s_108), .O(gate127inter3));
  inv1  gate1307(.a(s_109), .O(gate127inter4));
  nand2 gate1308(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1309(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1310(.a(G406), .O(gate127inter7));
  inv1  gate1311(.a(G407), .O(gate127inter8));
  nand2 gate1312(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1313(.a(s_109), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1314(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1315(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1316(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate2479(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2480(.a(gate128inter0), .b(s_276), .O(gate128inter1));
  and2  gate2481(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2482(.a(s_276), .O(gate128inter3));
  inv1  gate2483(.a(s_277), .O(gate128inter4));
  nand2 gate2484(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2485(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2486(.a(G408), .O(gate128inter7));
  inv1  gate2487(.a(G409), .O(gate128inter8));
  nand2 gate2488(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2489(.a(s_277), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2490(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2491(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2492(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate911(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate912(.a(gate132inter0), .b(s_52), .O(gate132inter1));
  and2  gate913(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate914(.a(s_52), .O(gate132inter3));
  inv1  gate915(.a(s_53), .O(gate132inter4));
  nand2 gate916(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate917(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate918(.a(G416), .O(gate132inter7));
  inv1  gate919(.a(G417), .O(gate132inter8));
  nand2 gate920(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate921(.a(s_53), .b(gate132inter3), .O(gate132inter10));
  nor2  gate922(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate923(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate924(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2535(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2536(.a(gate137inter0), .b(s_284), .O(gate137inter1));
  and2  gate2537(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2538(.a(s_284), .O(gate137inter3));
  inv1  gate2539(.a(s_285), .O(gate137inter4));
  nand2 gate2540(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2541(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2542(.a(G426), .O(gate137inter7));
  inv1  gate2543(.a(G429), .O(gate137inter8));
  nand2 gate2544(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2545(.a(s_285), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2546(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2547(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2548(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1849(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1850(.a(gate139inter0), .b(s_186), .O(gate139inter1));
  and2  gate1851(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1852(.a(s_186), .O(gate139inter3));
  inv1  gate1853(.a(s_187), .O(gate139inter4));
  nand2 gate1854(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1855(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1856(.a(G438), .O(gate139inter7));
  inv1  gate1857(.a(G441), .O(gate139inter8));
  nand2 gate1858(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1859(.a(s_187), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1860(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1861(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1862(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate813(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate814(.a(gate143inter0), .b(s_38), .O(gate143inter1));
  and2  gate815(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate816(.a(s_38), .O(gate143inter3));
  inv1  gate817(.a(s_39), .O(gate143inter4));
  nand2 gate818(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate819(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate820(.a(G462), .O(gate143inter7));
  inv1  gate821(.a(G465), .O(gate143inter8));
  nand2 gate822(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate823(.a(s_39), .b(gate143inter3), .O(gate143inter10));
  nor2  gate824(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate825(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate826(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1527(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1528(.a(gate146inter0), .b(s_140), .O(gate146inter1));
  and2  gate1529(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1530(.a(s_140), .O(gate146inter3));
  inv1  gate1531(.a(s_141), .O(gate146inter4));
  nand2 gate1532(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1533(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1534(.a(G480), .O(gate146inter7));
  inv1  gate1535(.a(G483), .O(gate146inter8));
  nand2 gate1536(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1537(.a(s_141), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1538(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1539(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1540(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2633(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2634(.a(gate147inter0), .b(s_298), .O(gate147inter1));
  and2  gate2635(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2636(.a(s_298), .O(gate147inter3));
  inv1  gate2637(.a(s_299), .O(gate147inter4));
  nand2 gate2638(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2639(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2640(.a(G486), .O(gate147inter7));
  inv1  gate2641(.a(G489), .O(gate147inter8));
  nand2 gate2642(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2643(.a(s_299), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2644(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2645(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2646(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1443(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1444(.a(gate149inter0), .b(s_128), .O(gate149inter1));
  and2  gate1445(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1446(.a(s_128), .O(gate149inter3));
  inv1  gate1447(.a(s_129), .O(gate149inter4));
  nand2 gate1448(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1449(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1450(.a(G498), .O(gate149inter7));
  inv1  gate1451(.a(G501), .O(gate149inter8));
  nand2 gate1452(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1453(.a(s_129), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1454(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1455(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1456(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1905(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1906(.a(gate156inter0), .b(s_194), .O(gate156inter1));
  and2  gate1907(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1908(.a(s_194), .O(gate156inter3));
  inv1  gate1909(.a(s_195), .O(gate156inter4));
  nand2 gate1910(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1911(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1912(.a(G435), .O(gate156inter7));
  inv1  gate1913(.a(G525), .O(gate156inter8));
  nand2 gate1914(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1915(.a(s_195), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1916(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1917(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1918(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate2255(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2256(.a(gate158inter0), .b(s_244), .O(gate158inter1));
  and2  gate2257(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2258(.a(s_244), .O(gate158inter3));
  inv1  gate2259(.a(s_245), .O(gate158inter4));
  nand2 gate2260(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2261(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2262(.a(G441), .O(gate158inter7));
  inv1  gate2263(.a(G528), .O(gate158inter8));
  nand2 gate2264(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2265(.a(s_245), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2266(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2267(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2268(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1247(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1248(.a(gate159inter0), .b(s_100), .O(gate159inter1));
  and2  gate1249(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1250(.a(s_100), .O(gate159inter3));
  inv1  gate1251(.a(s_101), .O(gate159inter4));
  nand2 gate1252(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1253(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1254(.a(G444), .O(gate159inter7));
  inv1  gate1255(.a(G531), .O(gate159inter8));
  nand2 gate1256(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1257(.a(s_101), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1258(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1259(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1260(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2157(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2158(.a(gate162inter0), .b(s_230), .O(gate162inter1));
  and2  gate2159(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2160(.a(s_230), .O(gate162inter3));
  inv1  gate2161(.a(s_231), .O(gate162inter4));
  nand2 gate2162(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2163(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2164(.a(G453), .O(gate162inter7));
  inv1  gate2165(.a(G534), .O(gate162inter8));
  nand2 gate2166(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2167(.a(s_231), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2168(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2169(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2170(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate1947(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1948(.a(gate163inter0), .b(s_200), .O(gate163inter1));
  and2  gate1949(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1950(.a(s_200), .O(gate163inter3));
  inv1  gate1951(.a(s_201), .O(gate163inter4));
  nand2 gate1952(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1953(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1954(.a(G456), .O(gate163inter7));
  inv1  gate1955(.a(G537), .O(gate163inter8));
  nand2 gate1956(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1957(.a(s_201), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1958(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1959(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1960(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate687(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate688(.a(gate164inter0), .b(s_20), .O(gate164inter1));
  and2  gate689(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate690(.a(s_20), .O(gate164inter3));
  inv1  gate691(.a(s_21), .O(gate164inter4));
  nand2 gate692(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate693(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate694(.a(G459), .O(gate164inter7));
  inv1  gate695(.a(G537), .O(gate164inter8));
  nand2 gate696(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate697(.a(s_21), .b(gate164inter3), .O(gate164inter10));
  nor2  gate698(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate699(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate700(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate1023(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1024(.a(gate165inter0), .b(s_68), .O(gate165inter1));
  and2  gate1025(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1026(.a(s_68), .O(gate165inter3));
  inv1  gate1027(.a(s_69), .O(gate165inter4));
  nand2 gate1028(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1029(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1030(.a(G462), .O(gate165inter7));
  inv1  gate1031(.a(G540), .O(gate165inter8));
  nand2 gate1032(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1033(.a(s_69), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1034(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1035(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1036(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2101(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2102(.a(gate168inter0), .b(s_222), .O(gate168inter1));
  and2  gate2103(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2104(.a(s_222), .O(gate168inter3));
  inv1  gate2105(.a(s_223), .O(gate168inter4));
  nand2 gate2106(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2107(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2108(.a(G471), .O(gate168inter7));
  inv1  gate2109(.a(G543), .O(gate168inter8));
  nand2 gate2110(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2111(.a(s_223), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2112(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2113(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2114(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1667(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1668(.a(gate172inter0), .b(s_160), .O(gate172inter1));
  and2  gate1669(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1670(.a(s_160), .O(gate172inter3));
  inv1  gate1671(.a(s_161), .O(gate172inter4));
  nand2 gate1672(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1673(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1674(.a(G483), .O(gate172inter7));
  inv1  gate1675(.a(G549), .O(gate172inter8));
  nand2 gate1676(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1677(.a(s_161), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1678(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1679(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1680(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1723(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1724(.a(gate178inter0), .b(s_168), .O(gate178inter1));
  and2  gate1725(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1726(.a(s_168), .O(gate178inter3));
  inv1  gate1727(.a(s_169), .O(gate178inter4));
  nand2 gate1728(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1729(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1730(.a(G501), .O(gate178inter7));
  inv1  gate1731(.a(G558), .O(gate178inter8));
  nand2 gate1732(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1733(.a(s_169), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1734(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1735(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1736(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2493(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2494(.a(gate181inter0), .b(s_278), .O(gate181inter1));
  and2  gate2495(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2496(.a(s_278), .O(gate181inter3));
  inv1  gate2497(.a(s_279), .O(gate181inter4));
  nand2 gate2498(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2499(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2500(.a(G510), .O(gate181inter7));
  inv1  gate2501(.a(G564), .O(gate181inter8));
  nand2 gate2502(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2503(.a(s_279), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2504(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2505(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2506(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1793(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1794(.a(gate182inter0), .b(s_178), .O(gate182inter1));
  and2  gate1795(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1796(.a(s_178), .O(gate182inter3));
  inv1  gate1797(.a(s_179), .O(gate182inter4));
  nand2 gate1798(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1799(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1800(.a(G513), .O(gate182inter7));
  inv1  gate1801(.a(G564), .O(gate182inter8));
  nand2 gate1802(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1803(.a(s_179), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1804(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1805(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1806(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate2003(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2004(.a(gate183inter0), .b(s_208), .O(gate183inter1));
  and2  gate2005(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2006(.a(s_208), .O(gate183inter3));
  inv1  gate2007(.a(s_209), .O(gate183inter4));
  nand2 gate2008(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2009(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2010(.a(G516), .O(gate183inter7));
  inv1  gate2011(.a(G567), .O(gate183inter8));
  nand2 gate2012(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2013(.a(s_209), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2014(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2015(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2016(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1429(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1430(.a(gate184inter0), .b(s_126), .O(gate184inter1));
  and2  gate1431(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1432(.a(s_126), .O(gate184inter3));
  inv1  gate1433(.a(s_127), .O(gate184inter4));
  nand2 gate1434(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1435(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1436(.a(G519), .O(gate184inter7));
  inv1  gate1437(.a(G567), .O(gate184inter8));
  nand2 gate1438(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1439(.a(s_127), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1440(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1441(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1442(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1457(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1458(.a(gate186inter0), .b(s_130), .O(gate186inter1));
  and2  gate1459(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1460(.a(s_130), .O(gate186inter3));
  inv1  gate1461(.a(s_131), .O(gate186inter4));
  nand2 gate1462(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1463(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1464(.a(G572), .O(gate186inter7));
  inv1  gate1465(.a(G573), .O(gate186inter8));
  nand2 gate1466(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1467(.a(s_131), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1468(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1469(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1470(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate2955(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2956(.a(gate187inter0), .b(s_344), .O(gate187inter1));
  and2  gate2957(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2958(.a(s_344), .O(gate187inter3));
  inv1  gate2959(.a(s_345), .O(gate187inter4));
  nand2 gate2960(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2961(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2962(.a(G574), .O(gate187inter7));
  inv1  gate2963(.a(G575), .O(gate187inter8));
  nand2 gate2964(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2965(.a(s_345), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2966(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2967(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2968(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate673(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate674(.a(gate190inter0), .b(s_18), .O(gate190inter1));
  and2  gate675(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate676(.a(s_18), .O(gate190inter3));
  inv1  gate677(.a(s_19), .O(gate190inter4));
  nand2 gate678(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate679(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate680(.a(G580), .O(gate190inter7));
  inv1  gate681(.a(G581), .O(gate190inter8));
  nand2 gate682(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate683(.a(s_19), .b(gate190inter3), .O(gate190inter10));
  nor2  gate684(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate685(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate686(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1205(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1206(.a(gate191inter0), .b(s_94), .O(gate191inter1));
  and2  gate1207(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1208(.a(s_94), .O(gate191inter3));
  inv1  gate1209(.a(s_95), .O(gate191inter4));
  nand2 gate1210(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1211(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1212(.a(G582), .O(gate191inter7));
  inv1  gate1213(.a(G583), .O(gate191inter8));
  nand2 gate1214(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1215(.a(s_95), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1216(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1217(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1218(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2829(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2830(.a(gate192inter0), .b(s_326), .O(gate192inter1));
  and2  gate2831(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2832(.a(s_326), .O(gate192inter3));
  inv1  gate2833(.a(s_327), .O(gate192inter4));
  nand2 gate2834(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2835(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2836(.a(G584), .O(gate192inter7));
  inv1  gate2837(.a(G585), .O(gate192inter8));
  nand2 gate2838(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2839(.a(s_327), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2840(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2841(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2842(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate841(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate842(.a(gate193inter0), .b(s_42), .O(gate193inter1));
  and2  gate843(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate844(.a(s_42), .O(gate193inter3));
  inv1  gate845(.a(s_43), .O(gate193inter4));
  nand2 gate846(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate847(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate848(.a(G586), .O(gate193inter7));
  inv1  gate849(.a(G587), .O(gate193inter8));
  nand2 gate850(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate851(.a(s_43), .b(gate193inter3), .O(gate193inter10));
  nor2  gate852(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate853(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate854(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2045(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2046(.a(gate195inter0), .b(s_214), .O(gate195inter1));
  and2  gate2047(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2048(.a(s_214), .O(gate195inter3));
  inv1  gate2049(.a(s_215), .O(gate195inter4));
  nand2 gate2050(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2051(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2052(.a(G590), .O(gate195inter7));
  inv1  gate2053(.a(G591), .O(gate195inter8));
  nand2 gate2054(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2055(.a(s_215), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2056(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2057(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2058(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2857(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2858(.a(gate207inter0), .b(s_330), .O(gate207inter1));
  and2  gate2859(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2860(.a(s_330), .O(gate207inter3));
  inv1  gate2861(.a(s_331), .O(gate207inter4));
  nand2 gate2862(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2863(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2864(.a(G622), .O(gate207inter7));
  inv1  gate2865(.a(G632), .O(gate207inter8));
  nand2 gate2866(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2867(.a(s_331), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2868(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2869(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2870(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate743(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate744(.a(gate210inter0), .b(s_28), .O(gate210inter1));
  and2  gate745(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate746(.a(s_28), .O(gate210inter3));
  inv1  gate747(.a(s_29), .O(gate210inter4));
  nand2 gate748(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate749(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate750(.a(G607), .O(gate210inter7));
  inv1  gate751(.a(G666), .O(gate210inter8));
  nand2 gate752(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate753(.a(s_29), .b(gate210inter3), .O(gate210inter10));
  nor2  gate754(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate755(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate756(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate995(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate996(.a(gate211inter0), .b(s_64), .O(gate211inter1));
  and2  gate997(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate998(.a(s_64), .O(gate211inter3));
  inv1  gate999(.a(s_65), .O(gate211inter4));
  nand2 gate1000(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1001(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1002(.a(G612), .O(gate211inter7));
  inv1  gate1003(.a(G669), .O(gate211inter8));
  nand2 gate1004(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1005(.a(s_65), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1006(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1007(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1008(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1121(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1122(.a(gate212inter0), .b(s_82), .O(gate212inter1));
  and2  gate1123(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1124(.a(s_82), .O(gate212inter3));
  inv1  gate1125(.a(s_83), .O(gate212inter4));
  nand2 gate1126(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1127(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1128(.a(G617), .O(gate212inter7));
  inv1  gate1129(.a(G669), .O(gate212inter8));
  nand2 gate1130(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1131(.a(s_83), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1132(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1133(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1134(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate953(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate954(.a(gate214inter0), .b(s_58), .O(gate214inter1));
  and2  gate955(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate956(.a(s_58), .O(gate214inter3));
  inv1  gate957(.a(s_59), .O(gate214inter4));
  nand2 gate958(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate959(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate960(.a(G612), .O(gate214inter7));
  inv1  gate961(.a(G672), .O(gate214inter8));
  nand2 gate962(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate963(.a(s_59), .b(gate214inter3), .O(gate214inter10));
  nor2  gate964(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate965(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate966(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2311(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2312(.a(gate216inter0), .b(s_252), .O(gate216inter1));
  and2  gate2313(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2314(.a(s_252), .O(gate216inter3));
  inv1  gate2315(.a(s_253), .O(gate216inter4));
  nand2 gate2316(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2317(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2318(.a(G617), .O(gate216inter7));
  inv1  gate2319(.a(G675), .O(gate216inter8));
  nand2 gate2320(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2321(.a(s_253), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2322(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2323(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2324(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate771(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate772(.a(gate218inter0), .b(s_32), .O(gate218inter1));
  and2  gate773(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate774(.a(s_32), .O(gate218inter3));
  inv1  gate775(.a(s_33), .O(gate218inter4));
  nand2 gate776(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate777(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate778(.a(G627), .O(gate218inter7));
  inv1  gate779(.a(G678), .O(gate218inter8));
  nand2 gate780(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate781(.a(s_33), .b(gate218inter3), .O(gate218inter10));
  nor2  gate782(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate783(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate784(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1597(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1598(.a(gate224inter0), .b(s_150), .O(gate224inter1));
  and2  gate1599(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1600(.a(s_150), .O(gate224inter3));
  inv1  gate1601(.a(s_151), .O(gate224inter4));
  nand2 gate1602(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1603(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1604(.a(G637), .O(gate224inter7));
  inv1  gate1605(.a(G687), .O(gate224inter8));
  nand2 gate1606(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1607(.a(s_151), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1608(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1609(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1610(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1891(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1892(.a(gate225inter0), .b(s_192), .O(gate225inter1));
  and2  gate1893(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1894(.a(s_192), .O(gate225inter3));
  inv1  gate1895(.a(s_193), .O(gate225inter4));
  nand2 gate1896(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1897(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1898(.a(G690), .O(gate225inter7));
  inv1  gate1899(.a(G691), .O(gate225inter8));
  nand2 gate1900(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1901(.a(s_193), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1902(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1903(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1904(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1289(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1290(.a(gate228inter0), .b(s_106), .O(gate228inter1));
  and2  gate1291(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1292(.a(s_106), .O(gate228inter3));
  inv1  gate1293(.a(s_107), .O(gate228inter4));
  nand2 gate1294(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1295(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1296(.a(G696), .O(gate228inter7));
  inv1  gate1297(.a(G697), .O(gate228inter8));
  nand2 gate1298(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1299(.a(s_107), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1300(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1301(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1302(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2549(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2550(.a(gate234inter0), .b(s_286), .O(gate234inter1));
  and2  gate2551(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2552(.a(s_286), .O(gate234inter3));
  inv1  gate2553(.a(s_287), .O(gate234inter4));
  nand2 gate2554(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2555(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2556(.a(G245), .O(gate234inter7));
  inv1  gate2557(.a(G721), .O(gate234inter8));
  nand2 gate2558(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2559(.a(s_287), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2560(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2561(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2562(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2325(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2326(.a(gate238inter0), .b(s_254), .O(gate238inter1));
  and2  gate2327(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2328(.a(s_254), .O(gate238inter3));
  inv1  gate2329(.a(s_255), .O(gate238inter4));
  nand2 gate2330(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2331(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2332(.a(G257), .O(gate238inter7));
  inv1  gate2333(.a(G709), .O(gate238inter8));
  nand2 gate2334(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2335(.a(s_255), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2336(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2337(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2338(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1009(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1010(.a(gate240inter0), .b(s_66), .O(gate240inter1));
  and2  gate1011(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1012(.a(s_66), .O(gate240inter3));
  inv1  gate1013(.a(s_67), .O(gate240inter4));
  nand2 gate1014(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1015(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1016(.a(G263), .O(gate240inter7));
  inv1  gate1017(.a(G715), .O(gate240inter8));
  nand2 gate1018(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1019(.a(s_67), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1020(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1021(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1022(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1051(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1052(.a(gate245inter0), .b(s_72), .O(gate245inter1));
  and2  gate1053(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1054(.a(s_72), .O(gate245inter3));
  inv1  gate1055(.a(s_73), .O(gate245inter4));
  nand2 gate1056(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1057(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1058(.a(G248), .O(gate245inter7));
  inv1  gate1059(.a(G736), .O(gate245inter8));
  nand2 gate1060(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1061(.a(s_73), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1062(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1063(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1064(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2241(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2242(.a(gate246inter0), .b(s_242), .O(gate246inter1));
  and2  gate2243(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2244(.a(s_242), .O(gate246inter3));
  inv1  gate2245(.a(s_243), .O(gate246inter4));
  nand2 gate2246(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2247(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2248(.a(G724), .O(gate246inter7));
  inv1  gate2249(.a(G736), .O(gate246inter8));
  nand2 gate2250(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2251(.a(s_243), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2252(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2253(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2254(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1233(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1234(.a(gate249inter0), .b(s_98), .O(gate249inter1));
  and2  gate1235(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1236(.a(s_98), .O(gate249inter3));
  inv1  gate1237(.a(s_99), .O(gate249inter4));
  nand2 gate1238(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1239(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1240(.a(G254), .O(gate249inter7));
  inv1  gate1241(.a(G742), .O(gate249inter8));
  nand2 gate1242(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1243(.a(s_99), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1244(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1245(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1246(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2801(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2802(.a(gate250inter0), .b(s_322), .O(gate250inter1));
  and2  gate2803(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2804(.a(s_322), .O(gate250inter3));
  inv1  gate2805(.a(s_323), .O(gate250inter4));
  nand2 gate2806(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2807(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2808(.a(G706), .O(gate250inter7));
  inv1  gate2809(.a(G742), .O(gate250inter8));
  nand2 gate2810(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2811(.a(s_323), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2812(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2813(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2814(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate631(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate632(.a(gate251inter0), .b(s_12), .O(gate251inter1));
  and2  gate633(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate634(.a(s_12), .O(gate251inter3));
  inv1  gate635(.a(s_13), .O(gate251inter4));
  nand2 gate636(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate637(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate638(.a(G257), .O(gate251inter7));
  inv1  gate639(.a(G745), .O(gate251inter8));
  nand2 gate640(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate641(.a(s_13), .b(gate251inter3), .O(gate251inter10));
  nor2  gate642(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate643(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate644(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1569(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1570(.a(gate255inter0), .b(s_146), .O(gate255inter1));
  and2  gate1571(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1572(.a(s_146), .O(gate255inter3));
  inv1  gate1573(.a(s_147), .O(gate255inter4));
  nand2 gate1574(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1575(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1576(.a(G263), .O(gate255inter7));
  inv1  gate1577(.a(G751), .O(gate255inter8));
  nand2 gate1578(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1579(.a(s_147), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1580(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1581(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1582(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2689(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2690(.a(gate257inter0), .b(s_306), .O(gate257inter1));
  and2  gate2691(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2692(.a(s_306), .O(gate257inter3));
  inv1  gate2693(.a(s_307), .O(gate257inter4));
  nand2 gate2694(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2695(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2696(.a(G754), .O(gate257inter7));
  inv1  gate2697(.a(G755), .O(gate257inter8));
  nand2 gate2698(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2699(.a(s_307), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2700(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2701(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2702(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1975(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1976(.a(gate258inter0), .b(s_204), .O(gate258inter1));
  and2  gate1977(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1978(.a(s_204), .O(gate258inter3));
  inv1  gate1979(.a(s_205), .O(gate258inter4));
  nand2 gate1980(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1981(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1982(.a(G756), .O(gate258inter7));
  inv1  gate1983(.a(G757), .O(gate258inter8));
  nand2 gate1984(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1985(.a(s_205), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1986(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1987(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1988(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate855(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate856(.a(gate259inter0), .b(s_44), .O(gate259inter1));
  and2  gate857(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate858(.a(s_44), .O(gate259inter3));
  inv1  gate859(.a(s_45), .O(gate259inter4));
  nand2 gate860(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate861(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate862(.a(G758), .O(gate259inter7));
  inv1  gate863(.a(G759), .O(gate259inter8));
  nand2 gate864(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate865(.a(s_45), .b(gate259inter3), .O(gate259inter10));
  nor2  gate866(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate867(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate868(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1219(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1220(.a(gate260inter0), .b(s_96), .O(gate260inter1));
  and2  gate1221(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1222(.a(s_96), .O(gate260inter3));
  inv1  gate1223(.a(s_97), .O(gate260inter4));
  nand2 gate1224(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1225(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1226(.a(G760), .O(gate260inter7));
  inv1  gate1227(.a(G761), .O(gate260inter8));
  nand2 gate1228(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1229(.a(s_97), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1230(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1231(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1232(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2507(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2508(.a(gate261inter0), .b(s_280), .O(gate261inter1));
  and2  gate2509(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2510(.a(s_280), .O(gate261inter3));
  inv1  gate2511(.a(s_281), .O(gate261inter4));
  nand2 gate2512(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2513(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2514(.a(G762), .O(gate261inter7));
  inv1  gate2515(.a(G763), .O(gate261inter8));
  nand2 gate2516(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2517(.a(s_281), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2518(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2519(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2520(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1401(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1402(.a(gate262inter0), .b(s_122), .O(gate262inter1));
  and2  gate1403(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1404(.a(s_122), .O(gate262inter3));
  inv1  gate1405(.a(s_123), .O(gate262inter4));
  nand2 gate1406(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1407(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1408(.a(G764), .O(gate262inter7));
  inv1  gate1409(.a(G765), .O(gate262inter8));
  nand2 gate1410(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1411(.a(s_123), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1412(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1413(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1414(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2997(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2998(.a(gate263inter0), .b(s_350), .O(gate263inter1));
  and2  gate2999(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate3000(.a(s_350), .O(gate263inter3));
  inv1  gate3001(.a(s_351), .O(gate263inter4));
  nand2 gate3002(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate3003(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate3004(.a(G766), .O(gate263inter7));
  inv1  gate3005(.a(G767), .O(gate263inter8));
  nand2 gate3006(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate3007(.a(s_351), .b(gate263inter3), .O(gate263inter10));
  nor2  gate3008(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate3009(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate3010(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2269(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2270(.a(gate264inter0), .b(s_246), .O(gate264inter1));
  and2  gate2271(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2272(.a(s_246), .O(gate264inter3));
  inv1  gate2273(.a(s_247), .O(gate264inter4));
  nand2 gate2274(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2275(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2276(.a(G768), .O(gate264inter7));
  inv1  gate2277(.a(G769), .O(gate264inter8));
  nand2 gate2278(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2279(.a(s_247), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2280(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2281(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2282(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate967(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate968(.a(gate265inter0), .b(s_60), .O(gate265inter1));
  and2  gate969(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate970(.a(s_60), .O(gate265inter3));
  inv1  gate971(.a(s_61), .O(gate265inter4));
  nand2 gate972(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate973(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate974(.a(G642), .O(gate265inter7));
  inv1  gate975(.a(G770), .O(gate265inter8));
  nand2 gate976(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate977(.a(s_61), .b(gate265inter3), .O(gate265inter10));
  nor2  gate978(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate979(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate980(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1107(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1108(.a(gate268inter0), .b(s_80), .O(gate268inter1));
  and2  gate1109(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1110(.a(s_80), .O(gate268inter3));
  inv1  gate1111(.a(s_81), .O(gate268inter4));
  nand2 gate1112(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1113(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1114(.a(G651), .O(gate268inter7));
  inv1  gate1115(.a(G779), .O(gate268inter8));
  nand2 gate1116(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1117(.a(s_81), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1118(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1119(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1120(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate883(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate884(.a(gate269inter0), .b(s_48), .O(gate269inter1));
  and2  gate885(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate886(.a(s_48), .O(gate269inter3));
  inv1  gate887(.a(s_49), .O(gate269inter4));
  nand2 gate888(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate889(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate890(.a(G654), .O(gate269inter7));
  inv1  gate891(.a(G782), .O(gate269inter8));
  nand2 gate892(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate893(.a(s_49), .b(gate269inter3), .O(gate269inter10));
  nor2  gate894(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate895(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate896(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1163(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1164(.a(gate273inter0), .b(s_88), .O(gate273inter1));
  and2  gate1165(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1166(.a(s_88), .O(gate273inter3));
  inv1  gate1167(.a(s_89), .O(gate273inter4));
  nand2 gate1168(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1169(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1170(.a(G642), .O(gate273inter7));
  inv1  gate1171(.a(G794), .O(gate273inter8));
  nand2 gate1172(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1173(.a(s_89), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1174(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1175(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1176(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2787(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2788(.a(gate276inter0), .b(s_320), .O(gate276inter1));
  and2  gate2789(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2790(.a(s_320), .O(gate276inter3));
  inv1  gate2791(.a(s_321), .O(gate276inter4));
  nand2 gate2792(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2793(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2794(.a(G773), .O(gate276inter7));
  inv1  gate2795(.a(G797), .O(gate276inter8));
  nand2 gate2796(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2797(.a(s_321), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2798(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2799(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2800(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate2381(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2382(.a(gate277inter0), .b(s_262), .O(gate277inter1));
  and2  gate2383(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2384(.a(s_262), .O(gate277inter3));
  inv1  gate2385(.a(s_263), .O(gate277inter4));
  nand2 gate2386(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2387(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2388(.a(G648), .O(gate277inter7));
  inv1  gate2389(.a(G800), .O(gate277inter8));
  nand2 gate2390(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2391(.a(s_263), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2392(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2393(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2394(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2213(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2214(.a(gate279inter0), .b(s_238), .O(gate279inter1));
  and2  gate2215(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2216(.a(s_238), .O(gate279inter3));
  inv1  gate2217(.a(s_239), .O(gate279inter4));
  nand2 gate2218(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2219(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2220(.a(G651), .O(gate279inter7));
  inv1  gate2221(.a(G803), .O(gate279inter8));
  nand2 gate2222(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2223(.a(s_239), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2224(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2225(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2226(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1135(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1136(.a(gate281inter0), .b(s_84), .O(gate281inter1));
  and2  gate1137(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1138(.a(s_84), .O(gate281inter3));
  inv1  gate1139(.a(s_85), .O(gate281inter4));
  nand2 gate1140(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1141(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1142(.a(G654), .O(gate281inter7));
  inv1  gate1143(.a(G806), .O(gate281inter8));
  nand2 gate1144(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1145(.a(s_85), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1146(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1147(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1148(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate2885(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2886(.a(gate284inter0), .b(s_334), .O(gate284inter1));
  and2  gate2887(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2888(.a(s_334), .O(gate284inter3));
  inv1  gate2889(.a(s_335), .O(gate284inter4));
  nand2 gate2890(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2891(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2892(.a(G785), .O(gate284inter7));
  inv1  gate2893(.a(G809), .O(gate284inter8));
  nand2 gate2894(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2895(.a(s_335), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2896(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2897(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2898(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1681(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1682(.a(gate285inter0), .b(s_162), .O(gate285inter1));
  and2  gate1683(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1684(.a(s_162), .O(gate285inter3));
  inv1  gate1685(.a(s_163), .O(gate285inter4));
  nand2 gate1686(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1687(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1688(.a(G660), .O(gate285inter7));
  inv1  gate1689(.a(G812), .O(gate285inter8));
  nand2 gate1690(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1691(.a(s_163), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1692(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1693(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1694(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1513(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1514(.a(gate286inter0), .b(s_138), .O(gate286inter1));
  and2  gate1515(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1516(.a(s_138), .O(gate286inter3));
  inv1  gate1517(.a(s_139), .O(gate286inter4));
  nand2 gate1518(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1519(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1520(.a(G788), .O(gate286inter7));
  inv1  gate1521(.a(G812), .O(gate286inter8));
  nand2 gate1522(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1523(.a(s_139), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1524(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1525(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1526(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate981(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate982(.a(gate290inter0), .b(s_62), .O(gate290inter1));
  and2  gate983(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate984(.a(s_62), .O(gate290inter3));
  inv1  gate985(.a(s_63), .O(gate290inter4));
  nand2 gate986(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate987(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate988(.a(G820), .O(gate290inter7));
  inv1  gate989(.a(G821), .O(gate290inter8));
  nand2 gate990(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate991(.a(s_63), .b(gate290inter3), .O(gate290inter10));
  nor2  gate992(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate993(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate994(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2143(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2144(.a(gate293inter0), .b(s_228), .O(gate293inter1));
  and2  gate2145(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2146(.a(s_228), .O(gate293inter3));
  inv1  gate2147(.a(s_229), .O(gate293inter4));
  nand2 gate2148(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2149(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2150(.a(G828), .O(gate293inter7));
  inv1  gate2151(.a(G829), .O(gate293inter8));
  nand2 gate2152(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2153(.a(s_229), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2154(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2155(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2156(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2059(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2060(.a(gate294inter0), .b(s_216), .O(gate294inter1));
  and2  gate2061(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2062(.a(s_216), .O(gate294inter3));
  inv1  gate2063(.a(s_217), .O(gate294inter4));
  nand2 gate2064(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2065(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2066(.a(G832), .O(gate294inter7));
  inv1  gate2067(.a(G833), .O(gate294inter8));
  nand2 gate2068(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2069(.a(s_217), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2070(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2071(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2072(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2941(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2942(.a(gate388inter0), .b(s_342), .O(gate388inter1));
  and2  gate2943(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2944(.a(s_342), .O(gate388inter3));
  inv1  gate2945(.a(s_343), .O(gate388inter4));
  nand2 gate2946(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2947(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2948(.a(G2), .O(gate388inter7));
  inv1  gate2949(.a(G1039), .O(gate388inter8));
  nand2 gate2950(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2951(.a(s_343), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2952(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2953(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2954(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2353(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2354(.a(gate392inter0), .b(s_258), .O(gate392inter1));
  and2  gate2355(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2356(.a(s_258), .O(gate392inter3));
  inv1  gate2357(.a(s_259), .O(gate392inter4));
  nand2 gate2358(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2359(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2360(.a(G6), .O(gate392inter7));
  inv1  gate2361(.a(G1051), .O(gate392inter8));
  nand2 gate2362(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2363(.a(s_259), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2364(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2365(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2366(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1751(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1752(.a(gate395inter0), .b(s_172), .O(gate395inter1));
  and2  gate1753(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1754(.a(s_172), .O(gate395inter3));
  inv1  gate1755(.a(s_173), .O(gate395inter4));
  nand2 gate1756(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1757(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1758(.a(G9), .O(gate395inter7));
  inv1  gate1759(.a(G1060), .O(gate395inter8));
  nand2 gate1760(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1761(.a(s_173), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1762(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1763(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1764(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2647(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2648(.a(gate397inter0), .b(s_300), .O(gate397inter1));
  and2  gate2649(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2650(.a(s_300), .O(gate397inter3));
  inv1  gate2651(.a(s_301), .O(gate397inter4));
  nand2 gate2652(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2653(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2654(.a(G11), .O(gate397inter7));
  inv1  gate2655(.a(G1066), .O(gate397inter8));
  nand2 gate2656(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2657(.a(s_301), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2658(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2659(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2660(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1737(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1738(.a(gate398inter0), .b(s_170), .O(gate398inter1));
  and2  gate1739(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1740(.a(s_170), .O(gate398inter3));
  inv1  gate1741(.a(s_171), .O(gate398inter4));
  nand2 gate1742(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1743(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1744(.a(G12), .O(gate398inter7));
  inv1  gate1745(.a(G1069), .O(gate398inter8));
  nand2 gate1746(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1747(.a(s_171), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1748(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1749(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1750(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2717(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2718(.a(gate400inter0), .b(s_310), .O(gate400inter1));
  and2  gate2719(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2720(.a(s_310), .O(gate400inter3));
  inv1  gate2721(.a(s_311), .O(gate400inter4));
  nand2 gate2722(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2723(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2724(.a(G14), .O(gate400inter7));
  inv1  gate2725(.a(G1075), .O(gate400inter8));
  nand2 gate2726(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2727(.a(s_311), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2728(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2729(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2730(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1149(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1150(.a(gate401inter0), .b(s_86), .O(gate401inter1));
  and2  gate1151(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1152(.a(s_86), .O(gate401inter3));
  inv1  gate1153(.a(s_87), .O(gate401inter4));
  nand2 gate1154(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1155(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1156(.a(G15), .O(gate401inter7));
  inv1  gate1157(.a(G1078), .O(gate401inter8));
  nand2 gate1158(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1159(.a(s_87), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1160(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1161(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1162(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate617(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate618(.a(gate406inter0), .b(s_10), .O(gate406inter1));
  and2  gate619(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate620(.a(s_10), .O(gate406inter3));
  inv1  gate621(.a(s_11), .O(gate406inter4));
  nand2 gate622(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate623(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate624(.a(G20), .O(gate406inter7));
  inv1  gate625(.a(G1093), .O(gate406inter8));
  nand2 gate626(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate627(.a(s_11), .b(gate406inter3), .O(gate406inter10));
  nor2  gate628(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate629(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate630(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1317(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1318(.a(gate407inter0), .b(s_110), .O(gate407inter1));
  and2  gate1319(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1320(.a(s_110), .O(gate407inter3));
  inv1  gate1321(.a(s_111), .O(gate407inter4));
  nand2 gate1322(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1323(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1324(.a(G21), .O(gate407inter7));
  inv1  gate1325(.a(G1096), .O(gate407inter8));
  nand2 gate1326(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1327(.a(s_111), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1328(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1329(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1330(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2521(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2522(.a(gate409inter0), .b(s_282), .O(gate409inter1));
  and2  gate2523(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2524(.a(s_282), .O(gate409inter3));
  inv1  gate2525(.a(s_283), .O(gate409inter4));
  nand2 gate2526(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2527(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2528(.a(G23), .O(gate409inter7));
  inv1  gate2529(.a(G1102), .O(gate409inter8));
  nand2 gate2530(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2531(.a(s_283), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2532(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2533(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2534(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2563(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2564(.a(gate412inter0), .b(s_288), .O(gate412inter1));
  and2  gate2565(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2566(.a(s_288), .O(gate412inter3));
  inv1  gate2567(.a(s_289), .O(gate412inter4));
  nand2 gate2568(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2569(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2570(.a(G26), .O(gate412inter7));
  inv1  gate2571(.a(G1111), .O(gate412inter8));
  nand2 gate2572(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2573(.a(s_289), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2574(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2575(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2576(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate827(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate828(.a(gate413inter0), .b(s_40), .O(gate413inter1));
  and2  gate829(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate830(.a(s_40), .O(gate413inter3));
  inv1  gate831(.a(s_41), .O(gate413inter4));
  nand2 gate832(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate833(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate834(.a(G27), .O(gate413inter7));
  inv1  gate835(.a(G1114), .O(gate413inter8));
  nand2 gate836(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate837(.a(s_41), .b(gate413inter3), .O(gate413inter10));
  nor2  gate838(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate839(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate840(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2031(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2032(.a(gate414inter0), .b(s_212), .O(gate414inter1));
  and2  gate2033(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2034(.a(s_212), .O(gate414inter3));
  inv1  gate2035(.a(s_213), .O(gate414inter4));
  nand2 gate2036(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2037(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2038(.a(G28), .O(gate414inter7));
  inv1  gate2039(.a(G1117), .O(gate414inter8));
  nand2 gate2040(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2041(.a(s_213), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2042(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2043(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2044(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1989(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1990(.a(gate415inter0), .b(s_206), .O(gate415inter1));
  and2  gate1991(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1992(.a(s_206), .O(gate415inter3));
  inv1  gate1993(.a(s_207), .O(gate415inter4));
  nand2 gate1994(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1995(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1996(.a(G29), .O(gate415inter7));
  inv1  gate1997(.a(G1120), .O(gate415inter8));
  nand2 gate1998(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1999(.a(s_207), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2000(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2001(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2002(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate3053(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate3054(.a(gate416inter0), .b(s_358), .O(gate416inter1));
  and2  gate3055(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate3056(.a(s_358), .O(gate416inter3));
  inv1  gate3057(.a(s_359), .O(gate416inter4));
  nand2 gate3058(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate3059(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate3060(.a(G30), .O(gate416inter7));
  inv1  gate3061(.a(G1123), .O(gate416inter8));
  nand2 gate3062(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate3063(.a(s_359), .b(gate416inter3), .O(gate416inter10));
  nor2  gate3064(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate3065(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate3066(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2087(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2088(.a(gate418inter0), .b(s_220), .O(gate418inter1));
  and2  gate2089(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2090(.a(s_220), .O(gate418inter3));
  inv1  gate2091(.a(s_221), .O(gate418inter4));
  nand2 gate2092(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2093(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2094(.a(G32), .O(gate418inter7));
  inv1  gate2095(.a(G1129), .O(gate418inter8));
  nand2 gate2096(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2097(.a(s_221), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2098(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2099(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2100(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2619(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2620(.a(gate419inter0), .b(s_296), .O(gate419inter1));
  and2  gate2621(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2622(.a(s_296), .O(gate419inter3));
  inv1  gate2623(.a(s_297), .O(gate419inter4));
  nand2 gate2624(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2625(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2626(.a(G1), .O(gate419inter7));
  inv1  gate2627(.a(G1132), .O(gate419inter8));
  nand2 gate2628(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2629(.a(s_297), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2630(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2631(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2632(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2969(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2970(.a(gate420inter0), .b(s_346), .O(gate420inter1));
  and2  gate2971(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2972(.a(s_346), .O(gate420inter3));
  inv1  gate2973(.a(s_347), .O(gate420inter4));
  nand2 gate2974(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2975(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2976(.a(G1036), .O(gate420inter7));
  inv1  gate2977(.a(G1132), .O(gate420inter8));
  nand2 gate2978(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2979(.a(s_347), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2980(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2981(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2982(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2815(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2816(.a(gate422inter0), .b(s_324), .O(gate422inter1));
  and2  gate2817(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2818(.a(s_324), .O(gate422inter3));
  inv1  gate2819(.a(s_325), .O(gate422inter4));
  nand2 gate2820(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2821(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2822(.a(G1039), .O(gate422inter7));
  inv1  gate2823(.a(G1135), .O(gate422inter8));
  nand2 gate2824(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2825(.a(s_325), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2826(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2827(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2828(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1611(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1612(.a(gate423inter0), .b(s_152), .O(gate423inter1));
  and2  gate1613(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1614(.a(s_152), .O(gate423inter3));
  inv1  gate1615(.a(s_153), .O(gate423inter4));
  nand2 gate1616(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1617(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1618(.a(G3), .O(gate423inter7));
  inv1  gate1619(.a(G1138), .O(gate423inter8));
  nand2 gate1620(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1621(.a(s_153), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1622(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1623(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1624(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1275(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1276(.a(gate425inter0), .b(s_104), .O(gate425inter1));
  and2  gate1277(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1278(.a(s_104), .O(gate425inter3));
  inv1  gate1279(.a(s_105), .O(gate425inter4));
  nand2 gate1280(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1281(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1282(.a(G4), .O(gate425inter7));
  inv1  gate1283(.a(G1141), .O(gate425inter8));
  nand2 gate1284(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1285(.a(s_105), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1286(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1287(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1288(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate3109(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate3110(.a(gate427inter0), .b(s_366), .O(gate427inter1));
  and2  gate3111(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate3112(.a(s_366), .O(gate427inter3));
  inv1  gate3113(.a(s_367), .O(gate427inter4));
  nand2 gate3114(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate3115(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate3116(.a(G5), .O(gate427inter7));
  inv1  gate3117(.a(G1144), .O(gate427inter8));
  nand2 gate3118(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate3119(.a(s_367), .b(gate427inter3), .O(gate427inter10));
  nor2  gate3120(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate3121(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate3122(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate3011(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate3012(.a(gate429inter0), .b(s_352), .O(gate429inter1));
  and2  gate3013(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate3014(.a(s_352), .O(gate429inter3));
  inv1  gate3015(.a(s_353), .O(gate429inter4));
  nand2 gate3016(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate3017(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate3018(.a(G6), .O(gate429inter7));
  inv1  gate3019(.a(G1147), .O(gate429inter8));
  nand2 gate3020(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate3021(.a(s_353), .b(gate429inter3), .O(gate429inter10));
  nor2  gate3022(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate3023(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate3024(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2283(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2284(.a(gate432inter0), .b(s_248), .O(gate432inter1));
  and2  gate2285(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2286(.a(s_248), .O(gate432inter3));
  inv1  gate2287(.a(s_249), .O(gate432inter4));
  nand2 gate2288(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2289(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2290(.a(G1054), .O(gate432inter7));
  inv1  gate2291(.a(G1150), .O(gate432inter8));
  nand2 gate2292(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2293(.a(s_249), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2294(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2295(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2296(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1821(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1822(.a(gate433inter0), .b(s_182), .O(gate433inter1));
  and2  gate1823(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1824(.a(s_182), .O(gate433inter3));
  inv1  gate1825(.a(s_183), .O(gate433inter4));
  nand2 gate1826(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1827(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1828(.a(G8), .O(gate433inter7));
  inv1  gate1829(.a(G1153), .O(gate433inter8));
  nand2 gate1830(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1831(.a(s_183), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1832(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1833(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1834(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate715(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate716(.a(gate438inter0), .b(s_24), .O(gate438inter1));
  and2  gate717(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate718(.a(s_24), .O(gate438inter3));
  inv1  gate719(.a(s_25), .O(gate438inter4));
  nand2 gate720(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate721(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate722(.a(G1063), .O(gate438inter7));
  inv1  gate723(.a(G1159), .O(gate438inter8));
  nand2 gate724(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate725(.a(s_25), .b(gate438inter3), .O(gate438inter10));
  nor2  gate726(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate727(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate728(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate3039(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate3040(.a(gate440inter0), .b(s_356), .O(gate440inter1));
  and2  gate3041(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate3042(.a(s_356), .O(gate440inter3));
  inv1  gate3043(.a(s_357), .O(gate440inter4));
  nand2 gate3044(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate3045(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate3046(.a(G1066), .O(gate440inter7));
  inv1  gate3047(.a(G1162), .O(gate440inter8));
  nand2 gate3048(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate3049(.a(s_357), .b(gate440inter3), .O(gate440inter10));
  nor2  gate3050(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate3051(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate3052(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1583(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1584(.a(gate446inter0), .b(s_148), .O(gate446inter1));
  and2  gate1585(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1586(.a(s_148), .O(gate446inter3));
  inv1  gate1587(.a(s_149), .O(gate446inter4));
  nand2 gate1588(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1589(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1590(.a(G1075), .O(gate446inter7));
  inv1  gate1591(.a(G1171), .O(gate446inter8));
  nand2 gate1592(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1593(.a(s_149), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1594(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1595(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1596(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1961(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1962(.a(gate447inter0), .b(s_202), .O(gate447inter1));
  and2  gate1963(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1964(.a(s_202), .O(gate447inter3));
  inv1  gate1965(.a(s_203), .O(gate447inter4));
  nand2 gate1966(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1967(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1968(.a(G15), .O(gate447inter7));
  inv1  gate1969(.a(G1174), .O(gate447inter8));
  nand2 gate1970(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1971(.a(s_203), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1972(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1973(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1974(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate659(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate660(.a(gate449inter0), .b(s_16), .O(gate449inter1));
  and2  gate661(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate662(.a(s_16), .O(gate449inter3));
  inv1  gate663(.a(s_17), .O(gate449inter4));
  nand2 gate664(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate665(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate666(.a(G16), .O(gate449inter7));
  inv1  gate667(.a(G1177), .O(gate449inter8));
  nand2 gate668(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate669(.a(s_17), .b(gate449inter3), .O(gate449inter10));
  nor2  gate670(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate671(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate672(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2605(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2606(.a(gate451inter0), .b(s_294), .O(gate451inter1));
  and2  gate2607(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2608(.a(s_294), .O(gate451inter3));
  inv1  gate2609(.a(s_295), .O(gate451inter4));
  nand2 gate2610(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2611(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2612(.a(G17), .O(gate451inter7));
  inv1  gate2613(.a(G1180), .O(gate451inter8));
  nand2 gate2614(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2615(.a(s_295), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2616(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2617(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2618(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate589(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate590(.a(gate452inter0), .b(s_6), .O(gate452inter1));
  and2  gate591(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate592(.a(s_6), .O(gate452inter3));
  inv1  gate593(.a(s_7), .O(gate452inter4));
  nand2 gate594(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate595(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate596(.a(G1084), .O(gate452inter7));
  inv1  gate597(.a(G1180), .O(gate452inter8));
  nand2 gate598(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate599(.a(s_7), .b(gate452inter3), .O(gate452inter10));
  nor2  gate600(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate601(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate602(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2339(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2340(.a(gate460inter0), .b(s_256), .O(gate460inter1));
  and2  gate2341(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2342(.a(s_256), .O(gate460inter3));
  inv1  gate2343(.a(s_257), .O(gate460inter4));
  nand2 gate2344(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2345(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2346(.a(G1096), .O(gate460inter7));
  inv1  gate2347(.a(G1192), .O(gate460inter8));
  nand2 gate2348(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2349(.a(s_257), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2350(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2351(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2352(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate757(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate758(.a(gate462inter0), .b(s_30), .O(gate462inter1));
  and2  gate759(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate760(.a(s_30), .O(gate462inter3));
  inv1  gate761(.a(s_31), .O(gate462inter4));
  nand2 gate762(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate763(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate764(.a(G1099), .O(gate462inter7));
  inv1  gate765(.a(G1195), .O(gate462inter8));
  nand2 gate766(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate767(.a(s_31), .b(gate462inter3), .O(gate462inter10));
  nor2  gate768(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate769(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate770(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2745(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2746(.a(gate463inter0), .b(s_314), .O(gate463inter1));
  and2  gate2747(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2748(.a(s_314), .O(gate463inter3));
  inv1  gate2749(.a(s_315), .O(gate463inter4));
  nand2 gate2750(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2751(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2752(.a(G23), .O(gate463inter7));
  inv1  gate2753(.a(G1198), .O(gate463inter8));
  nand2 gate2754(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2755(.a(s_315), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2756(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2757(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2758(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2465(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2466(.a(gate469inter0), .b(s_274), .O(gate469inter1));
  and2  gate2467(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2468(.a(s_274), .O(gate469inter3));
  inv1  gate2469(.a(s_275), .O(gate469inter4));
  nand2 gate2470(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2471(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2472(.a(G26), .O(gate469inter7));
  inv1  gate2473(.a(G1207), .O(gate469inter8));
  nand2 gate2474(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2475(.a(s_275), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2476(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2477(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2478(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate1765(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1766(.a(gate470inter0), .b(s_174), .O(gate470inter1));
  and2  gate1767(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1768(.a(s_174), .O(gate470inter3));
  inv1  gate1769(.a(s_175), .O(gate470inter4));
  nand2 gate1770(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1771(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1772(.a(G1111), .O(gate470inter7));
  inv1  gate1773(.a(G1207), .O(gate470inter8));
  nand2 gate1774(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1775(.a(s_175), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1776(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1777(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1778(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1037(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1038(.a(gate471inter0), .b(s_70), .O(gate471inter1));
  and2  gate1039(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1040(.a(s_70), .O(gate471inter3));
  inv1  gate1041(.a(s_71), .O(gate471inter4));
  nand2 gate1042(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1043(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1044(.a(G27), .O(gate471inter7));
  inv1  gate1045(.a(G1210), .O(gate471inter8));
  nand2 gate1046(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1047(.a(s_71), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1048(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1049(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1050(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1373(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1374(.a(gate476inter0), .b(s_118), .O(gate476inter1));
  and2  gate1375(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1376(.a(s_118), .O(gate476inter3));
  inv1  gate1377(.a(s_119), .O(gate476inter4));
  nand2 gate1378(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1379(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1380(.a(G1120), .O(gate476inter7));
  inv1  gate1381(.a(G1216), .O(gate476inter8));
  nand2 gate1382(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1383(.a(s_119), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1384(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1385(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1386(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate2297(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2298(.a(gate477inter0), .b(s_250), .O(gate477inter1));
  and2  gate2299(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2300(.a(s_250), .O(gate477inter3));
  inv1  gate2301(.a(s_251), .O(gate477inter4));
  nand2 gate2302(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2303(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2304(.a(G30), .O(gate477inter7));
  inv1  gate2305(.a(G1219), .O(gate477inter8));
  nand2 gate2306(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2307(.a(s_251), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2308(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2309(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2310(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1695(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1696(.a(gate478inter0), .b(s_164), .O(gate478inter1));
  and2  gate1697(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1698(.a(s_164), .O(gate478inter3));
  inv1  gate1699(.a(s_165), .O(gate478inter4));
  nand2 gate1700(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1701(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1702(.a(G1123), .O(gate478inter7));
  inv1  gate1703(.a(G1219), .O(gate478inter8));
  nand2 gate1704(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1705(.a(s_165), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1706(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1707(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1708(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1415(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1416(.a(gate480inter0), .b(s_124), .O(gate480inter1));
  and2  gate1417(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1418(.a(s_124), .O(gate480inter3));
  inv1  gate1419(.a(s_125), .O(gate480inter4));
  nand2 gate1420(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1421(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1422(.a(G1126), .O(gate480inter7));
  inv1  gate1423(.a(G1222), .O(gate480inter8));
  nand2 gate1424(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1425(.a(s_125), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1426(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1427(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1428(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate3123(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate3124(.a(gate483inter0), .b(s_368), .O(gate483inter1));
  and2  gate3125(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate3126(.a(s_368), .O(gate483inter3));
  inv1  gate3127(.a(s_369), .O(gate483inter4));
  nand2 gate3128(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate3129(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate3130(.a(G1228), .O(gate483inter7));
  inv1  gate3131(.a(G1229), .O(gate483inter8));
  nand2 gate3132(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate3133(.a(s_369), .b(gate483inter3), .O(gate483inter10));
  nor2  gate3134(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate3135(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate3136(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate785(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate786(.a(gate484inter0), .b(s_34), .O(gate484inter1));
  and2  gate787(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate788(.a(s_34), .O(gate484inter3));
  inv1  gate789(.a(s_35), .O(gate484inter4));
  nand2 gate790(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate791(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate792(.a(G1230), .O(gate484inter7));
  inv1  gate793(.a(G1231), .O(gate484inter8));
  nand2 gate794(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate795(.a(s_35), .b(gate484inter3), .O(gate484inter10));
  nor2  gate796(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate797(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate798(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2017(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2018(.a(gate485inter0), .b(s_210), .O(gate485inter1));
  and2  gate2019(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2020(.a(s_210), .O(gate485inter3));
  inv1  gate2021(.a(s_211), .O(gate485inter4));
  nand2 gate2022(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2023(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2024(.a(G1232), .O(gate485inter7));
  inv1  gate2025(.a(G1233), .O(gate485inter8));
  nand2 gate2026(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2027(.a(s_211), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2028(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2029(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2030(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1499(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1500(.a(gate488inter0), .b(s_136), .O(gate488inter1));
  and2  gate1501(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1502(.a(s_136), .O(gate488inter3));
  inv1  gate1503(.a(s_137), .O(gate488inter4));
  nand2 gate1504(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1505(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1506(.a(G1238), .O(gate488inter7));
  inv1  gate1507(.a(G1239), .O(gate488inter8));
  nand2 gate1508(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1509(.a(s_137), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1510(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1511(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1512(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1877(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1878(.a(gate490inter0), .b(s_190), .O(gate490inter1));
  and2  gate1879(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1880(.a(s_190), .O(gate490inter3));
  inv1  gate1881(.a(s_191), .O(gate490inter4));
  nand2 gate1882(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1883(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1884(.a(G1242), .O(gate490inter7));
  inv1  gate1885(.a(G1243), .O(gate490inter8));
  nand2 gate1886(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1887(.a(s_191), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1888(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1889(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1890(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1331(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1332(.a(gate492inter0), .b(s_112), .O(gate492inter1));
  and2  gate1333(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1334(.a(s_112), .O(gate492inter3));
  inv1  gate1335(.a(s_113), .O(gate492inter4));
  nand2 gate1336(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1337(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1338(.a(G1246), .O(gate492inter7));
  inv1  gate1339(.a(G1247), .O(gate492inter8));
  nand2 gate1340(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1341(.a(s_113), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1342(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1343(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1344(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate3137(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate3138(.a(gate495inter0), .b(s_370), .O(gate495inter1));
  and2  gate3139(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate3140(.a(s_370), .O(gate495inter3));
  inv1  gate3141(.a(s_371), .O(gate495inter4));
  nand2 gate3142(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate3143(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate3144(.a(G1252), .O(gate495inter7));
  inv1  gate3145(.a(G1253), .O(gate495inter8));
  nand2 gate3146(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate3147(.a(s_371), .b(gate495inter3), .O(gate495inter10));
  nor2  gate3148(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate3149(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate3150(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2199(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2200(.a(gate497inter0), .b(s_236), .O(gate497inter1));
  and2  gate2201(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2202(.a(s_236), .O(gate497inter3));
  inv1  gate2203(.a(s_237), .O(gate497inter4));
  nand2 gate2204(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2205(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2206(.a(G1256), .O(gate497inter7));
  inv1  gate2207(.a(G1257), .O(gate497inter8));
  nand2 gate2208(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2209(.a(s_237), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2210(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2211(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2212(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1079(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1080(.a(gate498inter0), .b(s_76), .O(gate498inter1));
  and2  gate1081(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1082(.a(s_76), .O(gate498inter3));
  inv1  gate1083(.a(s_77), .O(gate498inter4));
  nand2 gate1084(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1085(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1086(.a(G1258), .O(gate498inter7));
  inv1  gate1087(.a(G1259), .O(gate498inter8));
  nand2 gate1088(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1089(.a(s_77), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1090(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1091(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1092(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2367(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2368(.a(gate502inter0), .b(s_260), .O(gate502inter1));
  and2  gate2369(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2370(.a(s_260), .O(gate502inter3));
  inv1  gate2371(.a(s_261), .O(gate502inter4));
  nand2 gate2372(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2373(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2374(.a(G1266), .O(gate502inter7));
  inv1  gate2375(.a(G1267), .O(gate502inter8));
  nand2 gate2376(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2377(.a(s_261), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2378(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2379(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2380(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1261(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1262(.a(gate503inter0), .b(s_102), .O(gate503inter1));
  and2  gate1263(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1264(.a(s_102), .O(gate503inter3));
  inv1  gate1265(.a(s_103), .O(gate503inter4));
  nand2 gate1266(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1267(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1268(.a(G1268), .O(gate503inter7));
  inv1  gate1269(.a(G1269), .O(gate503inter8));
  nand2 gate1270(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1271(.a(s_103), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1272(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1273(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1274(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2423(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2424(.a(gate505inter0), .b(s_268), .O(gate505inter1));
  and2  gate2425(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2426(.a(s_268), .O(gate505inter3));
  inv1  gate2427(.a(s_269), .O(gate505inter4));
  nand2 gate2428(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2429(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2430(.a(G1272), .O(gate505inter7));
  inv1  gate2431(.a(G1273), .O(gate505inter8));
  nand2 gate2432(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2433(.a(s_269), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2434(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2435(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2436(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1191(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1192(.a(gate506inter0), .b(s_92), .O(gate506inter1));
  and2  gate1193(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1194(.a(s_92), .O(gate506inter3));
  inv1  gate1195(.a(s_93), .O(gate506inter4));
  nand2 gate1196(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1197(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1198(.a(G1274), .O(gate506inter7));
  inv1  gate1199(.a(G1275), .O(gate506inter8));
  nand2 gate1200(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1201(.a(s_93), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1202(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1203(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1204(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2703(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2704(.a(gate508inter0), .b(s_308), .O(gate508inter1));
  and2  gate2705(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2706(.a(s_308), .O(gate508inter3));
  inv1  gate2707(.a(s_309), .O(gate508inter4));
  nand2 gate2708(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2709(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2710(.a(G1278), .O(gate508inter7));
  inv1  gate2711(.a(G1279), .O(gate508inter8));
  nand2 gate2712(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2713(.a(s_309), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2714(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2715(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2716(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2073(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2074(.a(gate509inter0), .b(s_218), .O(gate509inter1));
  and2  gate2075(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2076(.a(s_218), .O(gate509inter3));
  inv1  gate2077(.a(s_219), .O(gate509inter4));
  nand2 gate2078(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2079(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2080(.a(G1280), .O(gate509inter7));
  inv1  gate2081(.a(G1281), .O(gate509inter8));
  nand2 gate2082(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2083(.a(s_219), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2084(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2085(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2086(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate2451(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2452(.a(gate510inter0), .b(s_272), .O(gate510inter1));
  and2  gate2453(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2454(.a(s_272), .O(gate510inter3));
  inv1  gate2455(.a(s_273), .O(gate510inter4));
  nand2 gate2456(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2457(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2458(.a(G1282), .O(gate510inter7));
  inv1  gate2459(.a(G1283), .O(gate510inter8));
  nand2 gate2460(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2461(.a(s_273), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2462(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2463(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2464(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1625(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1626(.a(gate512inter0), .b(s_154), .O(gate512inter1));
  and2  gate1627(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1628(.a(s_154), .O(gate512inter3));
  inv1  gate1629(.a(s_155), .O(gate512inter4));
  nand2 gate1630(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1631(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1632(.a(G1286), .O(gate512inter7));
  inv1  gate1633(.a(G1287), .O(gate512inter8));
  nand2 gate1634(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1635(.a(s_155), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1636(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1637(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1638(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate2759(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2760(.a(gate513inter0), .b(s_316), .O(gate513inter1));
  and2  gate2761(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2762(.a(s_316), .O(gate513inter3));
  inv1  gate2763(.a(s_317), .O(gate513inter4));
  nand2 gate2764(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2765(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2766(.a(G1288), .O(gate513inter7));
  inv1  gate2767(.a(G1289), .O(gate513inter8));
  nand2 gate2768(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2769(.a(s_317), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2770(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2771(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2772(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule