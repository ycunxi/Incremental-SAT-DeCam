module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate883(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate884(.a(gate9inter0), .b(s_48), .O(gate9inter1));
  and2  gate885(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate886(.a(s_48), .O(gate9inter3));
  inv1  gate887(.a(s_49), .O(gate9inter4));
  nand2 gate888(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate889(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate890(.a(G1), .O(gate9inter7));
  inv1  gate891(.a(G2), .O(gate9inter8));
  nand2 gate892(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate893(.a(s_49), .b(gate9inter3), .O(gate9inter10));
  nor2  gate894(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate895(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate896(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1093(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1094(.a(gate11inter0), .b(s_78), .O(gate11inter1));
  and2  gate1095(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1096(.a(s_78), .O(gate11inter3));
  inv1  gate1097(.a(s_79), .O(gate11inter4));
  nand2 gate1098(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1099(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1100(.a(G5), .O(gate11inter7));
  inv1  gate1101(.a(G6), .O(gate11inter8));
  nand2 gate1102(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1103(.a(s_79), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1104(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1105(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1106(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1261(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1262(.a(gate19inter0), .b(s_102), .O(gate19inter1));
  and2  gate1263(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1264(.a(s_102), .O(gate19inter3));
  inv1  gate1265(.a(s_103), .O(gate19inter4));
  nand2 gate1266(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1267(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1268(.a(G21), .O(gate19inter7));
  inv1  gate1269(.a(G22), .O(gate19inter8));
  nand2 gate1270(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1271(.a(s_103), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1272(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1273(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1274(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate575(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate576(.a(gate26inter0), .b(s_4), .O(gate26inter1));
  and2  gate577(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate578(.a(s_4), .O(gate26inter3));
  inv1  gate579(.a(s_5), .O(gate26inter4));
  nand2 gate580(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate581(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate582(.a(G9), .O(gate26inter7));
  inv1  gate583(.a(G13), .O(gate26inter8));
  nand2 gate584(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate585(.a(s_5), .b(gate26inter3), .O(gate26inter10));
  nor2  gate586(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate587(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate588(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1863(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1864(.a(gate29inter0), .b(s_188), .O(gate29inter1));
  and2  gate1865(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1866(.a(s_188), .O(gate29inter3));
  inv1  gate1867(.a(s_189), .O(gate29inter4));
  nand2 gate1868(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1869(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1870(.a(G3), .O(gate29inter7));
  inv1  gate1871(.a(G7), .O(gate29inter8));
  nand2 gate1872(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1873(.a(s_189), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1874(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1875(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1876(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1583(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1584(.a(gate37inter0), .b(s_148), .O(gate37inter1));
  and2  gate1585(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1586(.a(s_148), .O(gate37inter3));
  inv1  gate1587(.a(s_149), .O(gate37inter4));
  nand2 gate1588(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1589(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1590(.a(G19), .O(gate37inter7));
  inv1  gate1591(.a(G23), .O(gate37inter8));
  nand2 gate1592(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1593(.a(s_149), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1594(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1595(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1596(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1233(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1234(.a(gate51inter0), .b(s_98), .O(gate51inter1));
  and2  gate1235(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1236(.a(s_98), .O(gate51inter3));
  inv1  gate1237(.a(s_99), .O(gate51inter4));
  nand2 gate1238(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1239(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1240(.a(G11), .O(gate51inter7));
  inv1  gate1241(.a(G281), .O(gate51inter8));
  nand2 gate1242(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1243(.a(s_99), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1244(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1245(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1246(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1275(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1276(.a(gate60inter0), .b(s_104), .O(gate60inter1));
  and2  gate1277(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1278(.a(s_104), .O(gate60inter3));
  inv1  gate1279(.a(s_105), .O(gate60inter4));
  nand2 gate1280(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1281(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1282(.a(G20), .O(gate60inter7));
  inv1  gate1283(.a(G293), .O(gate60inter8));
  nand2 gate1284(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1285(.a(s_105), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1286(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1287(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1288(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate617(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate618(.a(gate61inter0), .b(s_10), .O(gate61inter1));
  and2  gate619(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate620(.a(s_10), .O(gate61inter3));
  inv1  gate621(.a(s_11), .O(gate61inter4));
  nand2 gate622(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate623(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate624(.a(G21), .O(gate61inter7));
  inv1  gate625(.a(G296), .O(gate61inter8));
  nand2 gate626(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate627(.a(s_11), .b(gate61inter3), .O(gate61inter10));
  nor2  gate628(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate629(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate630(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate799(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate800(.a(gate67inter0), .b(s_36), .O(gate67inter1));
  and2  gate801(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate802(.a(s_36), .O(gate67inter3));
  inv1  gate803(.a(s_37), .O(gate67inter4));
  nand2 gate804(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate805(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate806(.a(G27), .O(gate67inter7));
  inv1  gate807(.a(G305), .O(gate67inter8));
  nand2 gate808(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate809(.a(s_37), .b(gate67inter3), .O(gate67inter10));
  nor2  gate810(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate811(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate812(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate701(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate702(.a(gate68inter0), .b(s_22), .O(gate68inter1));
  and2  gate703(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate704(.a(s_22), .O(gate68inter3));
  inv1  gate705(.a(s_23), .O(gate68inter4));
  nand2 gate706(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate707(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate708(.a(G28), .O(gate68inter7));
  inv1  gate709(.a(G305), .O(gate68inter8));
  nand2 gate710(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate711(.a(s_23), .b(gate68inter3), .O(gate68inter10));
  nor2  gate712(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate713(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate714(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1513(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1514(.a(gate71inter0), .b(s_138), .O(gate71inter1));
  and2  gate1515(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1516(.a(s_138), .O(gate71inter3));
  inv1  gate1517(.a(s_139), .O(gate71inter4));
  nand2 gate1518(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1519(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1520(.a(G31), .O(gate71inter7));
  inv1  gate1521(.a(G311), .O(gate71inter8));
  nand2 gate1522(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1523(.a(s_139), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1524(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1525(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1526(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1163(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1164(.a(gate76inter0), .b(s_88), .O(gate76inter1));
  and2  gate1165(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1166(.a(s_88), .O(gate76inter3));
  inv1  gate1167(.a(s_89), .O(gate76inter4));
  nand2 gate1168(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1169(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1170(.a(G13), .O(gate76inter7));
  inv1  gate1171(.a(G317), .O(gate76inter8));
  nand2 gate1172(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1173(.a(s_89), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1174(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1175(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1176(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate771(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate772(.a(gate80inter0), .b(s_32), .O(gate80inter1));
  and2  gate773(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate774(.a(s_32), .O(gate80inter3));
  inv1  gate775(.a(s_33), .O(gate80inter4));
  nand2 gate776(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate777(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate778(.a(G14), .O(gate80inter7));
  inv1  gate779(.a(G323), .O(gate80inter8));
  nand2 gate780(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate781(.a(s_33), .b(gate80inter3), .O(gate80inter10));
  nor2  gate782(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate783(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate784(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1121(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1122(.a(gate83inter0), .b(s_82), .O(gate83inter1));
  and2  gate1123(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1124(.a(s_82), .O(gate83inter3));
  inv1  gate1125(.a(s_83), .O(gate83inter4));
  nand2 gate1126(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1127(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1128(.a(G11), .O(gate83inter7));
  inv1  gate1129(.a(G329), .O(gate83inter8));
  nand2 gate1130(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1131(.a(s_83), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1132(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1133(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1134(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1639(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1640(.a(gate88inter0), .b(s_156), .O(gate88inter1));
  and2  gate1641(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1642(.a(s_156), .O(gate88inter3));
  inv1  gate1643(.a(s_157), .O(gate88inter4));
  nand2 gate1644(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1645(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1646(.a(G16), .O(gate88inter7));
  inv1  gate1647(.a(G335), .O(gate88inter8));
  nand2 gate1648(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1649(.a(s_157), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1650(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1651(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1652(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1149(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1150(.a(gate98inter0), .b(s_86), .O(gate98inter1));
  and2  gate1151(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1152(.a(s_86), .O(gate98inter3));
  inv1  gate1153(.a(s_87), .O(gate98inter4));
  nand2 gate1154(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1155(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1156(.a(G23), .O(gate98inter7));
  inv1  gate1157(.a(G350), .O(gate98inter8));
  nand2 gate1158(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1159(.a(s_87), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1160(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1161(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1162(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate939(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate940(.a(gate106inter0), .b(s_56), .O(gate106inter1));
  and2  gate941(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate942(.a(s_56), .O(gate106inter3));
  inv1  gate943(.a(s_57), .O(gate106inter4));
  nand2 gate944(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate945(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate946(.a(G364), .O(gate106inter7));
  inv1  gate947(.a(G365), .O(gate106inter8));
  nand2 gate948(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate949(.a(s_57), .b(gate106inter3), .O(gate106inter10));
  nor2  gate950(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate951(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate952(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1023(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1024(.a(gate110inter0), .b(s_68), .O(gate110inter1));
  and2  gate1025(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1026(.a(s_68), .O(gate110inter3));
  inv1  gate1027(.a(s_69), .O(gate110inter4));
  nand2 gate1028(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1029(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1030(.a(G372), .O(gate110inter7));
  inv1  gate1031(.a(G373), .O(gate110inter8));
  nand2 gate1032(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1033(.a(s_69), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1034(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1035(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1036(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1569(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1570(.a(gate114inter0), .b(s_146), .O(gate114inter1));
  and2  gate1571(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1572(.a(s_146), .O(gate114inter3));
  inv1  gate1573(.a(s_147), .O(gate114inter4));
  nand2 gate1574(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1575(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1576(.a(G380), .O(gate114inter7));
  inv1  gate1577(.a(G381), .O(gate114inter8));
  nand2 gate1578(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1579(.a(s_147), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1580(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1581(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1582(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1765(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1766(.a(gate115inter0), .b(s_174), .O(gate115inter1));
  and2  gate1767(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1768(.a(s_174), .O(gate115inter3));
  inv1  gate1769(.a(s_175), .O(gate115inter4));
  nand2 gate1770(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1771(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1772(.a(G382), .O(gate115inter7));
  inv1  gate1773(.a(G383), .O(gate115inter8));
  nand2 gate1774(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1775(.a(s_175), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1776(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1777(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1778(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1345(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1346(.a(gate119inter0), .b(s_114), .O(gate119inter1));
  and2  gate1347(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1348(.a(s_114), .O(gate119inter3));
  inv1  gate1349(.a(s_115), .O(gate119inter4));
  nand2 gate1350(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1351(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1352(.a(G390), .O(gate119inter7));
  inv1  gate1353(.a(G391), .O(gate119inter8));
  nand2 gate1354(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1355(.a(s_115), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1356(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1357(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1358(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1877(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1878(.a(gate135inter0), .b(s_190), .O(gate135inter1));
  and2  gate1879(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1880(.a(s_190), .O(gate135inter3));
  inv1  gate1881(.a(s_191), .O(gate135inter4));
  nand2 gate1882(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1883(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1884(.a(G422), .O(gate135inter7));
  inv1  gate1885(.a(G423), .O(gate135inter8));
  nand2 gate1886(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1887(.a(s_191), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1888(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1889(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1890(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1555(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1556(.a(gate147inter0), .b(s_144), .O(gate147inter1));
  and2  gate1557(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1558(.a(s_144), .O(gate147inter3));
  inv1  gate1559(.a(s_145), .O(gate147inter4));
  nand2 gate1560(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1561(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1562(.a(G486), .O(gate147inter7));
  inv1  gate1563(.a(G489), .O(gate147inter8));
  nand2 gate1564(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1565(.a(s_145), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1566(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1567(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1568(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1359(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1360(.a(gate149inter0), .b(s_116), .O(gate149inter1));
  and2  gate1361(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1362(.a(s_116), .O(gate149inter3));
  inv1  gate1363(.a(s_117), .O(gate149inter4));
  nand2 gate1364(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1365(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1366(.a(G498), .O(gate149inter7));
  inv1  gate1367(.a(G501), .O(gate149inter8));
  nand2 gate1368(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1369(.a(s_117), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1370(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1371(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1372(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1499(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1500(.a(gate153inter0), .b(s_136), .O(gate153inter1));
  and2  gate1501(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1502(.a(s_136), .O(gate153inter3));
  inv1  gate1503(.a(s_137), .O(gate153inter4));
  nand2 gate1504(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1505(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1506(.a(G426), .O(gate153inter7));
  inv1  gate1507(.a(G522), .O(gate153inter8));
  nand2 gate1508(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1509(.a(s_137), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1510(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1511(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1512(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1793(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1794(.a(gate154inter0), .b(s_178), .O(gate154inter1));
  and2  gate1795(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1796(.a(s_178), .O(gate154inter3));
  inv1  gate1797(.a(s_179), .O(gate154inter4));
  nand2 gate1798(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1799(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1800(.a(G429), .O(gate154inter7));
  inv1  gate1801(.a(G522), .O(gate154inter8));
  nand2 gate1802(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1803(.a(s_179), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1804(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1805(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1806(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1331(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1332(.a(gate156inter0), .b(s_112), .O(gate156inter1));
  and2  gate1333(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1334(.a(s_112), .O(gate156inter3));
  inv1  gate1335(.a(s_113), .O(gate156inter4));
  nand2 gate1336(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1337(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1338(.a(G435), .O(gate156inter7));
  inv1  gate1339(.a(G525), .O(gate156inter8));
  nand2 gate1340(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1341(.a(s_113), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1342(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1343(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1344(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1177(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1178(.a(gate162inter0), .b(s_90), .O(gate162inter1));
  and2  gate1179(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1180(.a(s_90), .O(gate162inter3));
  inv1  gate1181(.a(s_91), .O(gate162inter4));
  nand2 gate1182(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1183(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1184(.a(G453), .O(gate162inter7));
  inv1  gate1185(.a(G534), .O(gate162inter8));
  nand2 gate1186(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1187(.a(s_91), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1188(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1189(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1190(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate841(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate842(.a(gate165inter0), .b(s_42), .O(gate165inter1));
  and2  gate843(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate844(.a(s_42), .O(gate165inter3));
  inv1  gate845(.a(s_43), .O(gate165inter4));
  nand2 gate846(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate847(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate848(.a(G462), .O(gate165inter7));
  inv1  gate849(.a(G540), .O(gate165inter8));
  nand2 gate850(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate851(.a(s_43), .b(gate165inter3), .O(gate165inter10));
  nor2  gate852(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate853(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate854(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1611(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1612(.a(gate166inter0), .b(s_152), .O(gate166inter1));
  and2  gate1613(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1614(.a(s_152), .O(gate166inter3));
  inv1  gate1615(.a(s_153), .O(gate166inter4));
  nand2 gate1616(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1617(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1618(.a(G465), .O(gate166inter7));
  inv1  gate1619(.a(G540), .O(gate166inter8));
  nand2 gate1620(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1621(.a(s_153), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1622(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1623(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1624(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate729(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate730(.a(gate167inter0), .b(s_26), .O(gate167inter1));
  and2  gate731(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate732(.a(s_26), .O(gate167inter3));
  inv1  gate733(.a(s_27), .O(gate167inter4));
  nand2 gate734(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate735(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate736(.a(G468), .O(gate167inter7));
  inv1  gate737(.a(G543), .O(gate167inter8));
  nand2 gate738(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate739(.a(s_27), .b(gate167inter3), .O(gate167inter10));
  nor2  gate740(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate741(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate742(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1079(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1080(.a(gate170inter0), .b(s_76), .O(gate170inter1));
  and2  gate1081(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1082(.a(s_76), .O(gate170inter3));
  inv1  gate1083(.a(s_77), .O(gate170inter4));
  nand2 gate1084(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1085(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1086(.a(G477), .O(gate170inter7));
  inv1  gate1087(.a(G546), .O(gate170inter8));
  nand2 gate1088(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1089(.a(s_77), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1090(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1091(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1092(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate981(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate982(.a(gate173inter0), .b(s_62), .O(gate173inter1));
  and2  gate983(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate984(.a(s_62), .O(gate173inter3));
  inv1  gate985(.a(s_63), .O(gate173inter4));
  nand2 gate986(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate987(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate988(.a(G486), .O(gate173inter7));
  inv1  gate989(.a(G552), .O(gate173inter8));
  nand2 gate990(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate991(.a(s_63), .b(gate173inter3), .O(gate173inter10));
  nor2  gate992(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate993(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate994(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate757(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate758(.a(gate174inter0), .b(s_30), .O(gate174inter1));
  and2  gate759(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate760(.a(s_30), .O(gate174inter3));
  inv1  gate761(.a(s_31), .O(gate174inter4));
  nand2 gate762(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate763(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate764(.a(G489), .O(gate174inter7));
  inv1  gate765(.a(G552), .O(gate174inter8));
  nand2 gate766(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate767(.a(s_31), .b(gate174inter3), .O(gate174inter10));
  nor2  gate768(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate769(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate770(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate995(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate996(.a(gate180inter0), .b(s_64), .O(gate180inter1));
  and2  gate997(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate998(.a(s_64), .O(gate180inter3));
  inv1  gate999(.a(s_65), .O(gate180inter4));
  nand2 gate1000(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1001(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1002(.a(G507), .O(gate180inter7));
  inv1  gate1003(.a(G561), .O(gate180inter8));
  nand2 gate1004(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1005(.a(s_65), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1006(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1007(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1008(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1835(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1836(.a(gate186inter0), .b(s_184), .O(gate186inter1));
  and2  gate1837(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1838(.a(s_184), .O(gate186inter3));
  inv1  gate1839(.a(s_185), .O(gate186inter4));
  nand2 gate1840(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1841(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1842(.a(G572), .O(gate186inter7));
  inv1  gate1843(.a(G573), .O(gate186inter8));
  nand2 gate1844(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1845(.a(s_185), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1846(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1847(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1848(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1429(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1430(.a(gate188inter0), .b(s_126), .O(gate188inter1));
  and2  gate1431(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1432(.a(s_126), .O(gate188inter3));
  inv1  gate1433(.a(s_127), .O(gate188inter4));
  nand2 gate1434(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1435(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1436(.a(G576), .O(gate188inter7));
  inv1  gate1437(.a(G577), .O(gate188inter8));
  nand2 gate1438(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1439(.a(s_127), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1440(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1441(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1442(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1457(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1458(.a(gate189inter0), .b(s_130), .O(gate189inter1));
  and2  gate1459(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1460(.a(s_130), .O(gate189inter3));
  inv1  gate1461(.a(s_131), .O(gate189inter4));
  nand2 gate1462(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1463(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1464(.a(G578), .O(gate189inter7));
  inv1  gate1465(.a(G579), .O(gate189inter8));
  nand2 gate1466(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1467(.a(s_131), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1468(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1469(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1470(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1849(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1850(.a(gate193inter0), .b(s_186), .O(gate193inter1));
  and2  gate1851(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1852(.a(s_186), .O(gate193inter3));
  inv1  gate1853(.a(s_187), .O(gate193inter4));
  nand2 gate1854(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1855(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1856(.a(G586), .O(gate193inter7));
  inv1  gate1857(.a(G587), .O(gate193inter8));
  nand2 gate1858(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1859(.a(s_187), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1860(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1861(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1862(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1485(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1486(.a(gate194inter0), .b(s_134), .O(gate194inter1));
  and2  gate1487(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1488(.a(s_134), .O(gate194inter3));
  inv1  gate1489(.a(s_135), .O(gate194inter4));
  nand2 gate1490(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1491(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1492(.a(G588), .O(gate194inter7));
  inv1  gate1493(.a(G589), .O(gate194inter8));
  nand2 gate1494(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1495(.a(s_135), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1496(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1497(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1498(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate827(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate828(.a(gate196inter0), .b(s_40), .O(gate196inter1));
  and2  gate829(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate830(.a(s_40), .O(gate196inter3));
  inv1  gate831(.a(s_41), .O(gate196inter4));
  nand2 gate832(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate833(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate834(.a(G592), .O(gate196inter7));
  inv1  gate835(.a(G593), .O(gate196inter8));
  nand2 gate836(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate837(.a(s_41), .b(gate196inter3), .O(gate196inter10));
  nor2  gate838(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate839(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate840(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate631(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate632(.a(gate197inter0), .b(s_12), .O(gate197inter1));
  and2  gate633(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate634(.a(s_12), .O(gate197inter3));
  inv1  gate635(.a(s_13), .O(gate197inter4));
  nand2 gate636(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate637(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate638(.a(G594), .O(gate197inter7));
  inv1  gate639(.a(G595), .O(gate197inter8));
  nand2 gate640(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate641(.a(s_13), .b(gate197inter3), .O(gate197inter10));
  nor2  gate642(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate643(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate644(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate897(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate898(.a(gate200inter0), .b(s_50), .O(gate200inter1));
  and2  gate899(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate900(.a(s_50), .O(gate200inter3));
  inv1  gate901(.a(s_51), .O(gate200inter4));
  nand2 gate902(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate903(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate904(.a(G600), .O(gate200inter7));
  inv1  gate905(.a(G601), .O(gate200inter8));
  nand2 gate906(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate907(.a(s_51), .b(gate200inter3), .O(gate200inter10));
  nor2  gate908(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate909(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate910(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1205(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1206(.a(gate211inter0), .b(s_94), .O(gate211inter1));
  and2  gate1207(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1208(.a(s_94), .O(gate211inter3));
  inv1  gate1209(.a(s_95), .O(gate211inter4));
  nand2 gate1210(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1211(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1212(.a(G612), .O(gate211inter7));
  inv1  gate1213(.a(G669), .O(gate211inter8));
  nand2 gate1214(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1215(.a(s_95), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1216(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1217(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1218(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1527(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1528(.a(gate215inter0), .b(s_140), .O(gate215inter1));
  and2  gate1529(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1530(.a(s_140), .O(gate215inter3));
  inv1  gate1531(.a(s_141), .O(gate215inter4));
  nand2 gate1532(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1533(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1534(.a(G607), .O(gate215inter7));
  inv1  gate1535(.a(G675), .O(gate215inter8));
  nand2 gate1536(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1537(.a(s_141), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1538(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1539(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1540(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate589(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate590(.a(gate221inter0), .b(s_6), .O(gate221inter1));
  and2  gate591(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate592(.a(s_6), .O(gate221inter3));
  inv1  gate593(.a(s_7), .O(gate221inter4));
  nand2 gate594(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate595(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate596(.a(G622), .O(gate221inter7));
  inv1  gate597(.a(G684), .O(gate221inter8));
  nand2 gate598(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate599(.a(s_7), .b(gate221inter3), .O(gate221inter10));
  nor2  gate600(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate601(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate602(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1779(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1780(.a(gate224inter0), .b(s_176), .O(gate224inter1));
  and2  gate1781(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1782(.a(s_176), .O(gate224inter3));
  inv1  gate1783(.a(s_177), .O(gate224inter4));
  nand2 gate1784(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1785(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1786(.a(G637), .O(gate224inter7));
  inv1  gate1787(.a(G687), .O(gate224inter8));
  nand2 gate1788(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1789(.a(s_177), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1790(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1791(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1792(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1191(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1192(.a(gate225inter0), .b(s_92), .O(gate225inter1));
  and2  gate1193(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1194(.a(s_92), .O(gate225inter3));
  inv1  gate1195(.a(s_93), .O(gate225inter4));
  nand2 gate1196(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1197(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1198(.a(G690), .O(gate225inter7));
  inv1  gate1199(.a(G691), .O(gate225inter8));
  nand2 gate1200(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1201(.a(s_93), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1202(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1203(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1204(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1443(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1444(.a(gate228inter0), .b(s_128), .O(gate228inter1));
  and2  gate1445(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1446(.a(s_128), .O(gate228inter3));
  inv1  gate1447(.a(s_129), .O(gate228inter4));
  nand2 gate1448(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1449(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1450(.a(G696), .O(gate228inter7));
  inv1  gate1451(.a(G697), .O(gate228inter8));
  nand2 gate1452(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1453(.a(s_129), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1454(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1455(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1456(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1065(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1066(.a(gate248inter0), .b(s_74), .O(gate248inter1));
  and2  gate1067(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1068(.a(s_74), .O(gate248inter3));
  inv1  gate1069(.a(s_75), .O(gate248inter4));
  nand2 gate1070(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1071(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1072(.a(G727), .O(gate248inter7));
  inv1  gate1073(.a(G739), .O(gate248inter8));
  nand2 gate1074(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1075(.a(s_75), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1076(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1077(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1078(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate547(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate548(.a(gate249inter0), .b(s_0), .O(gate249inter1));
  and2  gate549(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate550(.a(s_0), .O(gate249inter3));
  inv1  gate551(.a(s_1), .O(gate249inter4));
  nand2 gate552(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate553(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate554(.a(G254), .O(gate249inter7));
  inv1  gate555(.a(G742), .O(gate249inter8));
  nand2 gate556(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate557(.a(s_1), .b(gate249inter3), .O(gate249inter10));
  nor2  gate558(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate559(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate560(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1737(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1738(.a(gate256inter0), .b(s_170), .O(gate256inter1));
  and2  gate1739(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1740(.a(s_170), .O(gate256inter3));
  inv1  gate1741(.a(s_171), .O(gate256inter4));
  nand2 gate1742(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1743(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1744(.a(G715), .O(gate256inter7));
  inv1  gate1745(.a(G751), .O(gate256inter8));
  nand2 gate1746(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1747(.a(s_171), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1748(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1749(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1750(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1373(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1374(.a(gate260inter0), .b(s_118), .O(gate260inter1));
  and2  gate1375(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1376(.a(s_118), .O(gate260inter3));
  inv1  gate1377(.a(s_119), .O(gate260inter4));
  nand2 gate1378(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1379(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1380(.a(G760), .O(gate260inter7));
  inv1  gate1381(.a(G761), .O(gate260inter8));
  nand2 gate1382(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1383(.a(s_119), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1384(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1385(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1386(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1821(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1822(.a(gate261inter0), .b(s_182), .O(gate261inter1));
  and2  gate1823(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1824(.a(s_182), .O(gate261inter3));
  inv1  gate1825(.a(s_183), .O(gate261inter4));
  nand2 gate1826(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1827(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1828(.a(G762), .O(gate261inter7));
  inv1  gate1829(.a(G763), .O(gate261inter8));
  nand2 gate1830(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1831(.a(s_183), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1832(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1833(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1834(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate603(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate604(.a(gate263inter0), .b(s_8), .O(gate263inter1));
  and2  gate605(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate606(.a(s_8), .O(gate263inter3));
  inv1  gate607(.a(s_9), .O(gate263inter4));
  nand2 gate608(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate609(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate610(.a(G766), .O(gate263inter7));
  inv1  gate611(.a(G767), .O(gate263inter8));
  nand2 gate612(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate613(.a(s_9), .b(gate263inter3), .O(gate263inter10));
  nor2  gate614(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate615(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate616(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate785(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate786(.a(gate264inter0), .b(s_34), .O(gate264inter1));
  and2  gate787(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate788(.a(s_34), .O(gate264inter3));
  inv1  gate789(.a(s_35), .O(gate264inter4));
  nand2 gate790(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate791(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate792(.a(G768), .O(gate264inter7));
  inv1  gate793(.a(G769), .O(gate264inter8));
  nand2 gate794(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate795(.a(s_35), .b(gate264inter3), .O(gate264inter10));
  nor2  gate796(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate797(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate798(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate813(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate814(.a(gate271inter0), .b(s_38), .O(gate271inter1));
  and2  gate815(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate816(.a(s_38), .O(gate271inter3));
  inv1  gate817(.a(s_39), .O(gate271inter4));
  nand2 gate818(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate819(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate820(.a(G660), .O(gate271inter7));
  inv1  gate821(.a(G788), .O(gate271inter8));
  nand2 gate822(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate823(.a(s_39), .b(gate271inter3), .O(gate271inter10));
  nor2  gate824(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate825(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate826(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate925(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate926(.a(gate272inter0), .b(s_54), .O(gate272inter1));
  and2  gate927(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate928(.a(s_54), .O(gate272inter3));
  inv1  gate929(.a(s_55), .O(gate272inter4));
  nand2 gate930(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate931(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate932(.a(G663), .O(gate272inter7));
  inv1  gate933(.a(G791), .O(gate272inter8));
  nand2 gate934(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate935(.a(s_55), .b(gate272inter3), .O(gate272inter10));
  nor2  gate936(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate937(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate938(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate645(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate646(.a(gate274inter0), .b(s_14), .O(gate274inter1));
  and2  gate647(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate648(.a(s_14), .O(gate274inter3));
  inv1  gate649(.a(s_15), .O(gate274inter4));
  nand2 gate650(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate651(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate652(.a(G770), .O(gate274inter7));
  inv1  gate653(.a(G794), .O(gate274inter8));
  nand2 gate654(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate655(.a(s_15), .b(gate274inter3), .O(gate274inter10));
  nor2  gate656(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate657(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate658(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate869(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate870(.a(gate279inter0), .b(s_46), .O(gate279inter1));
  and2  gate871(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate872(.a(s_46), .O(gate279inter3));
  inv1  gate873(.a(s_47), .O(gate279inter4));
  nand2 gate874(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate875(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate876(.a(G651), .O(gate279inter7));
  inv1  gate877(.a(G803), .O(gate279inter8));
  nand2 gate878(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate879(.a(s_47), .b(gate279inter3), .O(gate279inter10));
  nor2  gate880(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate881(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate882(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1289(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1290(.a(gate283inter0), .b(s_106), .O(gate283inter1));
  and2  gate1291(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1292(.a(s_106), .O(gate283inter3));
  inv1  gate1293(.a(s_107), .O(gate283inter4));
  nand2 gate1294(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1295(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1296(.a(G657), .O(gate283inter7));
  inv1  gate1297(.a(G809), .O(gate283inter8));
  nand2 gate1298(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1299(.a(s_107), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1300(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1301(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1302(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate911(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate912(.a(gate284inter0), .b(s_52), .O(gate284inter1));
  and2  gate913(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate914(.a(s_52), .O(gate284inter3));
  inv1  gate915(.a(s_53), .O(gate284inter4));
  nand2 gate916(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate917(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate918(.a(G785), .O(gate284inter7));
  inv1  gate919(.a(G809), .O(gate284inter8));
  nand2 gate920(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate921(.a(s_53), .b(gate284inter3), .O(gate284inter10));
  nor2  gate922(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate923(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate924(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1653(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1654(.a(gate286inter0), .b(s_158), .O(gate286inter1));
  and2  gate1655(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1656(.a(s_158), .O(gate286inter3));
  inv1  gate1657(.a(s_159), .O(gate286inter4));
  nand2 gate1658(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1659(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1660(.a(G788), .O(gate286inter7));
  inv1  gate1661(.a(G812), .O(gate286inter8));
  nand2 gate1662(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1663(.a(s_159), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1664(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1665(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1666(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1751(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1752(.a(gate287inter0), .b(s_172), .O(gate287inter1));
  and2  gate1753(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1754(.a(s_172), .O(gate287inter3));
  inv1  gate1755(.a(s_173), .O(gate287inter4));
  nand2 gate1756(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1757(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1758(.a(G663), .O(gate287inter7));
  inv1  gate1759(.a(G815), .O(gate287inter8));
  nand2 gate1760(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1761(.a(s_173), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1762(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1763(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1764(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1009(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1010(.a(gate288inter0), .b(s_66), .O(gate288inter1));
  and2  gate1011(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1012(.a(s_66), .O(gate288inter3));
  inv1  gate1013(.a(s_67), .O(gate288inter4));
  nand2 gate1014(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1015(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1016(.a(G791), .O(gate288inter7));
  inv1  gate1017(.a(G815), .O(gate288inter8));
  nand2 gate1018(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1019(.a(s_67), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1020(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1021(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1022(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate673(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate674(.a(gate289inter0), .b(s_18), .O(gate289inter1));
  and2  gate675(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate676(.a(s_18), .O(gate289inter3));
  inv1  gate677(.a(s_19), .O(gate289inter4));
  nand2 gate678(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate679(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate680(.a(G818), .O(gate289inter7));
  inv1  gate681(.a(G819), .O(gate289inter8));
  nand2 gate682(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate683(.a(s_19), .b(gate289inter3), .O(gate289inter10));
  nor2  gate684(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate685(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate686(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1415(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1416(.a(gate387inter0), .b(s_124), .O(gate387inter1));
  and2  gate1417(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1418(.a(s_124), .O(gate387inter3));
  inv1  gate1419(.a(s_125), .O(gate387inter4));
  nand2 gate1420(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1421(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1422(.a(G1), .O(gate387inter7));
  inv1  gate1423(.a(G1036), .O(gate387inter8));
  nand2 gate1424(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1425(.a(s_125), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1426(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1427(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1428(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1709(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1710(.a(gate395inter0), .b(s_166), .O(gate395inter1));
  and2  gate1711(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1712(.a(s_166), .O(gate395inter3));
  inv1  gate1713(.a(s_167), .O(gate395inter4));
  nand2 gate1714(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1715(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1716(.a(G9), .O(gate395inter7));
  inv1  gate1717(.a(G1060), .O(gate395inter8));
  nand2 gate1718(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1719(.a(s_167), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1720(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1721(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1722(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate687(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate688(.a(gate396inter0), .b(s_20), .O(gate396inter1));
  and2  gate689(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate690(.a(s_20), .O(gate396inter3));
  inv1  gate691(.a(s_21), .O(gate396inter4));
  nand2 gate692(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate693(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate694(.a(G10), .O(gate396inter7));
  inv1  gate695(.a(G1063), .O(gate396inter8));
  nand2 gate696(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate697(.a(s_21), .b(gate396inter3), .O(gate396inter10));
  nor2  gate698(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate699(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate700(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1667(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1668(.a(gate397inter0), .b(s_160), .O(gate397inter1));
  and2  gate1669(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1670(.a(s_160), .O(gate397inter3));
  inv1  gate1671(.a(s_161), .O(gate397inter4));
  nand2 gate1672(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1673(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1674(.a(G11), .O(gate397inter7));
  inv1  gate1675(.a(G1066), .O(gate397inter8));
  nand2 gate1676(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1677(.a(s_161), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1678(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1679(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1680(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1387(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1388(.a(gate402inter0), .b(s_120), .O(gate402inter1));
  and2  gate1389(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1390(.a(s_120), .O(gate402inter3));
  inv1  gate1391(.a(s_121), .O(gate402inter4));
  nand2 gate1392(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1393(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1394(.a(G16), .O(gate402inter7));
  inv1  gate1395(.a(G1081), .O(gate402inter8));
  nand2 gate1396(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1397(.a(s_121), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1398(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1399(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1400(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1695(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1696(.a(gate410inter0), .b(s_164), .O(gate410inter1));
  and2  gate1697(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1698(.a(s_164), .O(gate410inter3));
  inv1  gate1699(.a(s_165), .O(gate410inter4));
  nand2 gate1700(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1701(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1702(.a(G24), .O(gate410inter7));
  inv1  gate1703(.a(G1105), .O(gate410inter8));
  nand2 gate1704(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1705(.a(s_165), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1706(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1707(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1708(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1107(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1108(.a(gate412inter0), .b(s_80), .O(gate412inter1));
  and2  gate1109(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1110(.a(s_80), .O(gate412inter3));
  inv1  gate1111(.a(s_81), .O(gate412inter4));
  nand2 gate1112(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1113(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1114(.a(G26), .O(gate412inter7));
  inv1  gate1115(.a(G1111), .O(gate412inter8));
  nand2 gate1116(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1117(.a(s_81), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1118(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1119(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1120(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate659(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate660(.a(gate419inter0), .b(s_16), .O(gate419inter1));
  and2  gate661(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate662(.a(s_16), .O(gate419inter3));
  inv1  gate663(.a(s_17), .O(gate419inter4));
  nand2 gate664(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate665(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate666(.a(G1), .O(gate419inter7));
  inv1  gate667(.a(G1132), .O(gate419inter8));
  nand2 gate668(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate669(.a(s_17), .b(gate419inter3), .O(gate419inter10));
  nor2  gate670(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate671(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate672(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1723(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1724(.a(gate422inter0), .b(s_168), .O(gate422inter1));
  and2  gate1725(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1726(.a(s_168), .O(gate422inter3));
  inv1  gate1727(.a(s_169), .O(gate422inter4));
  nand2 gate1728(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1729(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1730(.a(G1039), .O(gate422inter7));
  inv1  gate1731(.a(G1135), .O(gate422inter8));
  nand2 gate1732(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1733(.a(s_169), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1734(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1735(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1736(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1303(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1304(.a(gate428inter0), .b(s_108), .O(gate428inter1));
  and2  gate1305(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1306(.a(s_108), .O(gate428inter3));
  inv1  gate1307(.a(s_109), .O(gate428inter4));
  nand2 gate1308(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1309(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1310(.a(G1048), .O(gate428inter7));
  inv1  gate1311(.a(G1144), .O(gate428inter8));
  nand2 gate1312(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1313(.a(s_109), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1314(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1315(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1316(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1051(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1052(.a(gate432inter0), .b(s_72), .O(gate432inter1));
  and2  gate1053(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1054(.a(s_72), .O(gate432inter3));
  inv1  gate1055(.a(s_73), .O(gate432inter4));
  nand2 gate1056(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1057(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1058(.a(G1054), .O(gate432inter7));
  inv1  gate1059(.a(G1150), .O(gate432inter8));
  nand2 gate1060(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1061(.a(s_73), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1062(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1063(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1064(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1135(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1136(.a(gate438inter0), .b(s_84), .O(gate438inter1));
  and2  gate1137(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1138(.a(s_84), .O(gate438inter3));
  inv1  gate1139(.a(s_85), .O(gate438inter4));
  nand2 gate1140(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1141(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1142(.a(G1063), .O(gate438inter7));
  inv1  gate1143(.a(G1159), .O(gate438inter8));
  nand2 gate1144(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1145(.a(s_85), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1146(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1147(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1148(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate953(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate954(.a(gate452inter0), .b(s_58), .O(gate452inter1));
  and2  gate955(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate956(.a(s_58), .O(gate452inter3));
  inv1  gate957(.a(s_59), .O(gate452inter4));
  nand2 gate958(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate959(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate960(.a(G1084), .O(gate452inter7));
  inv1  gate961(.a(G1180), .O(gate452inter8));
  nand2 gate962(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate963(.a(s_59), .b(gate452inter3), .O(gate452inter10));
  nor2  gate964(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate965(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate966(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate715(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate716(.a(gate453inter0), .b(s_24), .O(gate453inter1));
  and2  gate717(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate718(.a(s_24), .O(gate453inter3));
  inv1  gate719(.a(s_25), .O(gate453inter4));
  nand2 gate720(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate721(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate722(.a(G18), .O(gate453inter7));
  inv1  gate723(.a(G1183), .O(gate453inter8));
  nand2 gate724(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate725(.a(s_25), .b(gate453inter3), .O(gate453inter10));
  nor2  gate726(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate727(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate728(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate561(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate562(.a(gate454inter0), .b(s_2), .O(gate454inter1));
  and2  gate563(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate564(.a(s_2), .O(gate454inter3));
  inv1  gate565(.a(s_3), .O(gate454inter4));
  nand2 gate566(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate567(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate568(.a(G1087), .O(gate454inter7));
  inv1  gate569(.a(G1183), .O(gate454inter8));
  nand2 gate570(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate571(.a(s_3), .b(gate454inter3), .O(gate454inter10));
  nor2  gate572(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate573(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate574(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1597(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1598(.a(gate458inter0), .b(s_150), .O(gate458inter1));
  and2  gate1599(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1600(.a(s_150), .O(gate458inter3));
  inv1  gate1601(.a(s_151), .O(gate458inter4));
  nand2 gate1602(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1603(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1604(.a(G1093), .O(gate458inter7));
  inv1  gate1605(.a(G1189), .O(gate458inter8));
  nand2 gate1606(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1607(.a(s_151), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1608(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1609(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1610(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1625(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1626(.a(gate463inter0), .b(s_154), .O(gate463inter1));
  and2  gate1627(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1628(.a(s_154), .O(gate463inter3));
  inv1  gate1629(.a(s_155), .O(gate463inter4));
  nand2 gate1630(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1631(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1632(.a(G23), .O(gate463inter7));
  inv1  gate1633(.a(G1198), .O(gate463inter8));
  nand2 gate1634(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1635(.a(s_155), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1636(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1637(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1638(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1247(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1248(.a(gate466inter0), .b(s_100), .O(gate466inter1));
  and2  gate1249(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1250(.a(s_100), .O(gate466inter3));
  inv1  gate1251(.a(s_101), .O(gate466inter4));
  nand2 gate1252(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1253(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1254(.a(G1105), .O(gate466inter7));
  inv1  gate1255(.a(G1201), .O(gate466inter8));
  nand2 gate1256(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1257(.a(s_101), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1258(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1259(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1260(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1471(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1472(.a(gate467inter0), .b(s_132), .O(gate467inter1));
  and2  gate1473(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1474(.a(s_132), .O(gate467inter3));
  inv1  gate1475(.a(s_133), .O(gate467inter4));
  nand2 gate1476(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1477(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1478(.a(G25), .O(gate467inter7));
  inv1  gate1479(.a(G1204), .O(gate467inter8));
  nand2 gate1480(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1481(.a(s_133), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1482(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1483(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1484(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate967(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate968(.a(gate475inter0), .b(s_60), .O(gate475inter1));
  and2  gate969(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate970(.a(s_60), .O(gate475inter3));
  inv1  gate971(.a(s_61), .O(gate475inter4));
  nand2 gate972(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate973(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate974(.a(G29), .O(gate475inter7));
  inv1  gate975(.a(G1216), .O(gate475inter8));
  nand2 gate976(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate977(.a(s_61), .b(gate475inter3), .O(gate475inter10));
  nor2  gate978(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate979(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate980(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1401(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1402(.a(gate477inter0), .b(s_122), .O(gate477inter1));
  and2  gate1403(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1404(.a(s_122), .O(gate477inter3));
  inv1  gate1405(.a(s_123), .O(gate477inter4));
  nand2 gate1406(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1407(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1408(.a(G30), .O(gate477inter7));
  inv1  gate1409(.a(G1219), .O(gate477inter8));
  nand2 gate1410(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1411(.a(s_123), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1412(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1413(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1414(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate743(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate744(.a(gate484inter0), .b(s_28), .O(gate484inter1));
  and2  gate745(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate746(.a(s_28), .O(gate484inter3));
  inv1  gate747(.a(s_29), .O(gate484inter4));
  nand2 gate748(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate749(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate750(.a(G1230), .O(gate484inter7));
  inv1  gate751(.a(G1231), .O(gate484inter8));
  nand2 gate752(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate753(.a(s_29), .b(gate484inter3), .O(gate484inter10));
  nor2  gate754(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate755(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate756(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1219(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1220(.a(gate491inter0), .b(s_96), .O(gate491inter1));
  and2  gate1221(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1222(.a(s_96), .O(gate491inter3));
  inv1  gate1223(.a(s_97), .O(gate491inter4));
  nand2 gate1224(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1225(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1226(.a(G1244), .O(gate491inter7));
  inv1  gate1227(.a(G1245), .O(gate491inter8));
  nand2 gate1228(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1229(.a(s_97), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1230(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1231(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1232(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1037(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1038(.a(gate493inter0), .b(s_70), .O(gate493inter1));
  and2  gate1039(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1040(.a(s_70), .O(gate493inter3));
  inv1  gate1041(.a(s_71), .O(gate493inter4));
  nand2 gate1042(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1043(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1044(.a(G1248), .O(gate493inter7));
  inv1  gate1045(.a(G1249), .O(gate493inter8));
  nand2 gate1046(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1047(.a(s_71), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1048(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1049(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1050(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1807(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1808(.a(gate496inter0), .b(s_180), .O(gate496inter1));
  and2  gate1809(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1810(.a(s_180), .O(gate496inter3));
  inv1  gate1811(.a(s_181), .O(gate496inter4));
  nand2 gate1812(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1813(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1814(.a(G1254), .O(gate496inter7));
  inv1  gate1815(.a(G1255), .O(gate496inter8));
  nand2 gate1816(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1817(.a(s_181), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1818(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1819(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1820(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate855(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate856(.a(gate501inter0), .b(s_44), .O(gate501inter1));
  and2  gate857(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate858(.a(s_44), .O(gate501inter3));
  inv1  gate859(.a(s_45), .O(gate501inter4));
  nand2 gate860(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate861(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate862(.a(G1264), .O(gate501inter7));
  inv1  gate863(.a(G1265), .O(gate501inter8));
  nand2 gate864(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate865(.a(s_45), .b(gate501inter3), .O(gate501inter10));
  nor2  gate866(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate867(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate868(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1541(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1542(.a(gate502inter0), .b(s_142), .O(gate502inter1));
  and2  gate1543(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1544(.a(s_142), .O(gate502inter3));
  inv1  gate1545(.a(s_143), .O(gate502inter4));
  nand2 gate1546(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1547(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1548(.a(G1266), .O(gate502inter7));
  inv1  gate1549(.a(G1267), .O(gate502inter8));
  nand2 gate1550(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1551(.a(s_143), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1552(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1553(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1554(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1681(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1682(.a(gate505inter0), .b(s_162), .O(gate505inter1));
  and2  gate1683(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1684(.a(s_162), .O(gate505inter3));
  inv1  gate1685(.a(s_163), .O(gate505inter4));
  nand2 gate1686(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1687(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1688(.a(G1272), .O(gate505inter7));
  inv1  gate1689(.a(G1273), .O(gate505inter8));
  nand2 gate1690(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1691(.a(s_163), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1692(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1693(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1694(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1317(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1318(.a(gate512inter0), .b(s_110), .O(gate512inter1));
  and2  gate1319(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1320(.a(s_110), .O(gate512inter3));
  inv1  gate1321(.a(s_111), .O(gate512inter4));
  nand2 gate1322(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1323(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1324(.a(G1286), .O(gate512inter7));
  inv1  gate1325(.a(G1287), .O(gate512inter8));
  nand2 gate1326(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1327(.a(s_111), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1328(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1329(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1330(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule