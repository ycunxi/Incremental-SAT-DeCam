module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate897(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate898(.a(gate9inter0), .b(s_50), .O(gate9inter1));
  and2  gate899(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate900(.a(s_50), .O(gate9inter3));
  inv1  gate901(.a(s_51), .O(gate9inter4));
  nand2 gate902(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate903(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate904(.a(G1), .O(gate9inter7));
  inv1  gate905(.a(G2), .O(gate9inter8));
  nand2 gate906(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate907(.a(s_51), .b(gate9inter3), .O(gate9inter10));
  nor2  gate908(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate909(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate910(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate841(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate842(.a(gate12inter0), .b(s_42), .O(gate12inter1));
  and2  gate843(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate844(.a(s_42), .O(gate12inter3));
  inv1  gate845(.a(s_43), .O(gate12inter4));
  nand2 gate846(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate847(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate848(.a(G7), .O(gate12inter7));
  inv1  gate849(.a(G8), .O(gate12inter8));
  nand2 gate850(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate851(.a(s_43), .b(gate12inter3), .O(gate12inter10));
  nor2  gate852(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate853(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate854(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1079(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1080(.a(gate19inter0), .b(s_76), .O(gate19inter1));
  and2  gate1081(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1082(.a(s_76), .O(gate19inter3));
  inv1  gate1083(.a(s_77), .O(gate19inter4));
  nand2 gate1084(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1085(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1086(.a(G21), .O(gate19inter7));
  inv1  gate1087(.a(G22), .O(gate19inter8));
  nand2 gate1088(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1089(.a(s_77), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1090(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1091(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1092(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate659(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate660(.a(gate24inter0), .b(s_16), .O(gate24inter1));
  and2  gate661(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate662(.a(s_16), .O(gate24inter3));
  inv1  gate663(.a(s_17), .O(gate24inter4));
  nand2 gate664(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate665(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate666(.a(G31), .O(gate24inter7));
  inv1  gate667(.a(G32), .O(gate24inter8));
  nand2 gate668(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate669(.a(s_17), .b(gate24inter3), .O(gate24inter10));
  nor2  gate670(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate671(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate672(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate687(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate688(.a(gate37inter0), .b(s_20), .O(gate37inter1));
  and2  gate689(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate690(.a(s_20), .O(gate37inter3));
  inv1  gate691(.a(s_21), .O(gate37inter4));
  nand2 gate692(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate693(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate694(.a(G19), .O(gate37inter7));
  inv1  gate695(.a(G23), .O(gate37inter8));
  nand2 gate696(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate697(.a(s_21), .b(gate37inter3), .O(gate37inter10));
  nor2  gate698(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate699(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate700(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1317(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1318(.a(gate41inter0), .b(s_110), .O(gate41inter1));
  and2  gate1319(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1320(.a(s_110), .O(gate41inter3));
  inv1  gate1321(.a(s_111), .O(gate41inter4));
  nand2 gate1322(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1323(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1324(.a(G1), .O(gate41inter7));
  inv1  gate1325(.a(G266), .O(gate41inter8));
  nand2 gate1326(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1327(.a(s_111), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1328(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1329(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1330(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate813(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate814(.a(gate42inter0), .b(s_38), .O(gate42inter1));
  and2  gate815(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate816(.a(s_38), .O(gate42inter3));
  inv1  gate817(.a(s_39), .O(gate42inter4));
  nand2 gate818(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate819(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate820(.a(G2), .O(gate42inter7));
  inv1  gate821(.a(G266), .O(gate42inter8));
  nand2 gate822(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate823(.a(s_39), .b(gate42inter3), .O(gate42inter10));
  nor2  gate824(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate825(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate826(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate603(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate604(.a(gate43inter0), .b(s_8), .O(gate43inter1));
  and2  gate605(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate606(.a(s_8), .O(gate43inter3));
  inv1  gate607(.a(s_9), .O(gate43inter4));
  nand2 gate608(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate609(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate610(.a(G3), .O(gate43inter7));
  inv1  gate611(.a(G269), .O(gate43inter8));
  nand2 gate612(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate613(.a(s_9), .b(gate43inter3), .O(gate43inter10));
  nor2  gate614(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate615(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate616(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate995(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate996(.a(gate47inter0), .b(s_64), .O(gate47inter1));
  and2  gate997(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate998(.a(s_64), .O(gate47inter3));
  inv1  gate999(.a(s_65), .O(gate47inter4));
  nand2 gate1000(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1001(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1002(.a(G7), .O(gate47inter7));
  inv1  gate1003(.a(G275), .O(gate47inter8));
  nand2 gate1004(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1005(.a(s_65), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1006(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1007(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1008(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate547(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate548(.a(gate57inter0), .b(s_0), .O(gate57inter1));
  and2  gate549(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate550(.a(s_0), .O(gate57inter3));
  inv1  gate551(.a(s_1), .O(gate57inter4));
  nand2 gate552(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate553(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate554(.a(G17), .O(gate57inter7));
  inv1  gate555(.a(G290), .O(gate57inter8));
  nand2 gate556(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate557(.a(s_1), .b(gate57inter3), .O(gate57inter10));
  nor2  gate558(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate559(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate560(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate645(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate646(.a(gate109inter0), .b(s_14), .O(gate109inter1));
  and2  gate647(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate648(.a(s_14), .O(gate109inter3));
  inv1  gate649(.a(s_15), .O(gate109inter4));
  nand2 gate650(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate651(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate652(.a(G370), .O(gate109inter7));
  inv1  gate653(.a(G371), .O(gate109inter8));
  nand2 gate654(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate655(.a(s_15), .b(gate109inter3), .O(gate109inter10));
  nor2  gate656(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate657(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate658(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1023(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1024(.a(gate117inter0), .b(s_68), .O(gate117inter1));
  and2  gate1025(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1026(.a(s_68), .O(gate117inter3));
  inv1  gate1027(.a(s_69), .O(gate117inter4));
  nand2 gate1028(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1029(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1030(.a(G386), .O(gate117inter7));
  inv1  gate1031(.a(G387), .O(gate117inter8));
  nand2 gate1032(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1033(.a(s_69), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1034(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1035(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1036(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1037(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1038(.a(gate126inter0), .b(s_70), .O(gate126inter1));
  and2  gate1039(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1040(.a(s_70), .O(gate126inter3));
  inv1  gate1041(.a(s_71), .O(gate126inter4));
  nand2 gate1042(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1043(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1044(.a(G404), .O(gate126inter7));
  inv1  gate1045(.a(G405), .O(gate126inter8));
  nand2 gate1046(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1047(.a(s_71), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1048(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1049(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1050(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate617(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate618(.a(gate129inter0), .b(s_10), .O(gate129inter1));
  and2  gate619(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate620(.a(s_10), .O(gate129inter3));
  inv1  gate621(.a(s_11), .O(gate129inter4));
  nand2 gate622(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate623(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate624(.a(G410), .O(gate129inter7));
  inv1  gate625(.a(G411), .O(gate129inter8));
  nand2 gate626(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate627(.a(s_11), .b(gate129inter3), .O(gate129inter10));
  nor2  gate628(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate629(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate630(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1233(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1234(.a(gate141inter0), .b(s_98), .O(gate141inter1));
  and2  gate1235(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1236(.a(s_98), .O(gate141inter3));
  inv1  gate1237(.a(s_99), .O(gate141inter4));
  nand2 gate1238(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1239(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1240(.a(G450), .O(gate141inter7));
  inv1  gate1241(.a(G453), .O(gate141inter8));
  nand2 gate1242(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1243(.a(s_99), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1244(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1245(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1246(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1163(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1164(.a(gate144inter0), .b(s_88), .O(gate144inter1));
  and2  gate1165(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1166(.a(s_88), .O(gate144inter3));
  inv1  gate1167(.a(s_89), .O(gate144inter4));
  nand2 gate1168(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1169(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1170(.a(G468), .O(gate144inter7));
  inv1  gate1171(.a(G471), .O(gate144inter8));
  nand2 gate1172(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1173(.a(s_89), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1174(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1175(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1176(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate673(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate674(.a(gate154inter0), .b(s_18), .O(gate154inter1));
  and2  gate675(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate676(.a(s_18), .O(gate154inter3));
  inv1  gate677(.a(s_19), .O(gate154inter4));
  nand2 gate678(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate679(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate680(.a(G429), .O(gate154inter7));
  inv1  gate681(.a(G522), .O(gate154inter8));
  nand2 gate682(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate683(.a(s_19), .b(gate154inter3), .O(gate154inter10));
  nor2  gate684(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate685(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate686(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1373(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1374(.a(gate156inter0), .b(s_118), .O(gate156inter1));
  and2  gate1375(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1376(.a(s_118), .O(gate156inter3));
  inv1  gate1377(.a(s_119), .O(gate156inter4));
  nand2 gate1378(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1379(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1380(.a(G435), .O(gate156inter7));
  inv1  gate1381(.a(G525), .O(gate156inter8));
  nand2 gate1382(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1383(.a(s_119), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1384(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1385(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1386(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate827(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate828(.a(gate160inter0), .b(s_40), .O(gate160inter1));
  and2  gate829(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate830(.a(s_40), .O(gate160inter3));
  inv1  gate831(.a(s_41), .O(gate160inter4));
  nand2 gate832(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate833(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate834(.a(G447), .O(gate160inter7));
  inv1  gate835(.a(G531), .O(gate160inter8));
  nand2 gate836(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate837(.a(s_41), .b(gate160inter3), .O(gate160inter10));
  nor2  gate838(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate839(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate840(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate561(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate562(.a(gate171inter0), .b(s_2), .O(gate171inter1));
  and2  gate563(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate564(.a(s_2), .O(gate171inter3));
  inv1  gate565(.a(s_3), .O(gate171inter4));
  nand2 gate566(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate567(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate568(.a(G480), .O(gate171inter7));
  inv1  gate569(.a(G549), .O(gate171inter8));
  nand2 gate570(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate571(.a(s_3), .b(gate171inter3), .O(gate171inter10));
  nor2  gate572(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate573(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate574(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1093(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1094(.a(gate182inter0), .b(s_78), .O(gate182inter1));
  and2  gate1095(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1096(.a(s_78), .O(gate182inter3));
  inv1  gate1097(.a(s_79), .O(gate182inter4));
  nand2 gate1098(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1099(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1100(.a(G513), .O(gate182inter7));
  inv1  gate1101(.a(G564), .O(gate182inter8));
  nand2 gate1102(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1103(.a(s_79), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1104(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1105(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1106(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate631(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate632(.a(gate208inter0), .b(s_12), .O(gate208inter1));
  and2  gate633(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate634(.a(s_12), .O(gate208inter3));
  inv1  gate635(.a(s_13), .O(gate208inter4));
  nand2 gate636(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate637(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate638(.a(G627), .O(gate208inter7));
  inv1  gate639(.a(G637), .O(gate208inter8));
  nand2 gate640(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate641(.a(s_13), .b(gate208inter3), .O(gate208inter10));
  nor2  gate642(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate643(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate644(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate715(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate716(.a(gate209inter0), .b(s_24), .O(gate209inter1));
  and2  gate717(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate718(.a(s_24), .O(gate209inter3));
  inv1  gate719(.a(s_25), .O(gate209inter4));
  nand2 gate720(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate721(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate722(.a(G602), .O(gate209inter7));
  inv1  gate723(.a(G666), .O(gate209inter8));
  nand2 gate724(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate725(.a(s_25), .b(gate209inter3), .O(gate209inter10));
  nor2  gate726(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate727(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate728(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1331(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1332(.a(gate216inter0), .b(s_112), .O(gate216inter1));
  and2  gate1333(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1334(.a(s_112), .O(gate216inter3));
  inv1  gate1335(.a(s_113), .O(gate216inter4));
  nand2 gate1336(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1337(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1338(.a(G617), .O(gate216inter7));
  inv1  gate1339(.a(G675), .O(gate216inter8));
  nand2 gate1340(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1341(.a(s_113), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1342(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1343(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1344(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate575(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate576(.a(gate219inter0), .b(s_4), .O(gate219inter1));
  and2  gate577(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate578(.a(s_4), .O(gate219inter3));
  inv1  gate579(.a(s_5), .O(gate219inter4));
  nand2 gate580(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate581(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate582(.a(G632), .O(gate219inter7));
  inv1  gate583(.a(G681), .O(gate219inter8));
  nand2 gate584(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate585(.a(s_5), .b(gate219inter3), .O(gate219inter10));
  nor2  gate586(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate587(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate588(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1065(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1066(.a(gate224inter0), .b(s_74), .O(gate224inter1));
  and2  gate1067(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1068(.a(s_74), .O(gate224inter3));
  inv1  gate1069(.a(s_75), .O(gate224inter4));
  nand2 gate1070(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1071(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1072(.a(G637), .O(gate224inter7));
  inv1  gate1073(.a(G687), .O(gate224inter8));
  nand2 gate1074(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1075(.a(s_75), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1076(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1077(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1078(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1177(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1178(.a(gate228inter0), .b(s_90), .O(gate228inter1));
  and2  gate1179(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1180(.a(s_90), .O(gate228inter3));
  inv1  gate1181(.a(s_91), .O(gate228inter4));
  nand2 gate1182(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1183(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1184(.a(G696), .O(gate228inter7));
  inv1  gate1185(.a(G697), .O(gate228inter8));
  nand2 gate1186(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1187(.a(s_91), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1188(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1189(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1190(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1275(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1276(.a(gate233inter0), .b(s_104), .O(gate233inter1));
  and2  gate1277(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1278(.a(s_104), .O(gate233inter3));
  inv1  gate1279(.a(s_105), .O(gate233inter4));
  nand2 gate1280(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1281(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1282(.a(G242), .O(gate233inter7));
  inv1  gate1283(.a(G718), .O(gate233inter8));
  nand2 gate1284(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1285(.a(s_105), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1286(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1287(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1288(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate785(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate786(.a(gate246inter0), .b(s_34), .O(gate246inter1));
  and2  gate787(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate788(.a(s_34), .O(gate246inter3));
  inv1  gate789(.a(s_35), .O(gate246inter4));
  nand2 gate790(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate791(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate792(.a(G724), .O(gate246inter7));
  inv1  gate793(.a(G736), .O(gate246inter8));
  nand2 gate794(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate795(.a(s_35), .b(gate246inter3), .O(gate246inter10));
  nor2  gate796(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate797(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate798(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1149(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1150(.a(gate250inter0), .b(s_86), .O(gate250inter1));
  and2  gate1151(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1152(.a(s_86), .O(gate250inter3));
  inv1  gate1153(.a(s_87), .O(gate250inter4));
  nand2 gate1154(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1155(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1156(.a(G706), .O(gate250inter7));
  inv1  gate1157(.a(G742), .O(gate250inter8));
  nand2 gate1158(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1159(.a(s_87), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1160(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1161(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1162(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1135(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1136(.a(gate257inter0), .b(s_84), .O(gate257inter1));
  and2  gate1137(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1138(.a(s_84), .O(gate257inter3));
  inv1  gate1139(.a(s_85), .O(gate257inter4));
  nand2 gate1140(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1141(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1142(.a(G754), .O(gate257inter7));
  inv1  gate1143(.a(G755), .O(gate257inter8));
  nand2 gate1144(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1145(.a(s_85), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1146(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1147(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1148(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate911(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate912(.a(gate260inter0), .b(s_52), .O(gate260inter1));
  and2  gate913(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate914(.a(s_52), .O(gate260inter3));
  inv1  gate915(.a(s_53), .O(gate260inter4));
  nand2 gate916(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate917(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate918(.a(G760), .O(gate260inter7));
  inv1  gate919(.a(G761), .O(gate260inter8));
  nand2 gate920(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate921(.a(s_53), .b(gate260inter3), .O(gate260inter10));
  nor2  gate922(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate923(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate924(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate771(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate772(.a(gate270inter0), .b(s_32), .O(gate270inter1));
  and2  gate773(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate774(.a(s_32), .O(gate270inter3));
  inv1  gate775(.a(s_33), .O(gate270inter4));
  nand2 gate776(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate777(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate778(.a(G657), .O(gate270inter7));
  inv1  gate779(.a(G785), .O(gate270inter8));
  nand2 gate780(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate781(.a(s_33), .b(gate270inter3), .O(gate270inter10));
  nor2  gate782(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate783(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate784(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate757(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate758(.a(gate285inter0), .b(s_30), .O(gate285inter1));
  and2  gate759(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate760(.a(s_30), .O(gate285inter3));
  inv1  gate761(.a(s_31), .O(gate285inter4));
  nand2 gate762(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate763(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate764(.a(G660), .O(gate285inter7));
  inv1  gate765(.a(G812), .O(gate285inter8));
  nand2 gate766(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate767(.a(s_31), .b(gate285inter3), .O(gate285inter10));
  nor2  gate768(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate769(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate770(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1051(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1052(.a(gate289inter0), .b(s_72), .O(gate289inter1));
  and2  gate1053(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1054(.a(s_72), .O(gate289inter3));
  inv1  gate1055(.a(s_73), .O(gate289inter4));
  nand2 gate1056(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1057(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1058(.a(G818), .O(gate289inter7));
  inv1  gate1059(.a(G819), .O(gate289inter8));
  nand2 gate1060(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1061(.a(s_73), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1062(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1063(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1064(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate869(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate870(.a(gate387inter0), .b(s_46), .O(gate387inter1));
  and2  gate871(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate872(.a(s_46), .O(gate387inter3));
  inv1  gate873(.a(s_47), .O(gate387inter4));
  nand2 gate874(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate875(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate876(.a(G1), .O(gate387inter7));
  inv1  gate877(.a(G1036), .O(gate387inter8));
  nand2 gate878(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate879(.a(s_47), .b(gate387inter3), .O(gate387inter10));
  nor2  gate880(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate881(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate882(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1121(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1122(.a(gate388inter0), .b(s_82), .O(gate388inter1));
  and2  gate1123(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1124(.a(s_82), .O(gate388inter3));
  inv1  gate1125(.a(s_83), .O(gate388inter4));
  nand2 gate1126(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1127(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1128(.a(G2), .O(gate388inter7));
  inv1  gate1129(.a(G1039), .O(gate388inter8));
  nand2 gate1130(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1131(.a(s_83), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1132(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1133(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1134(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate855(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate856(.a(gate397inter0), .b(s_44), .O(gate397inter1));
  and2  gate857(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate858(.a(s_44), .O(gate397inter3));
  inv1  gate859(.a(s_45), .O(gate397inter4));
  nand2 gate860(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate861(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate862(.a(G11), .O(gate397inter7));
  inv1  gate863(.a(G1066), .O(gate397inter8));
  nand2 gate864(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate865(.a(s_45), .b(gate397inter3), .O(gate397inter10));
  nor2  gate866(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate867(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate868(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1303(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1304(.a(gate405inter0), .b(s_108), .O(gate405inter1));
  and2  gate1305(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1306(.a(s_108), .O(gate405inter3));
  inv1  gate1307(.a(s_109), .O(gate405inter4));
  nand2 gate1308(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1309(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1310(.a(G19), .O(gate405inter7));
  inv1  gate1311(.a(G1090), .O(gate405inter8));
  nand2 gate1312(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1313(.a(s_109), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1314(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1315(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1316(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate939(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate940(.a(gate413inter0), .b(s_56), .O(gate413inter1));
  and2  gate941(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate942(.a(s_56), .O(gate413inter3));
  inv1  gate943(.a(s_57), .O(gate413inter4));
  nand2 gate944(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate945(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate946(.a(G27), .O(gate413inter7));
  inv1  gate947(.a(G1114), .O(gate413inter8));
  nand2 gate948(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate949(.a(s_57), .b(gate413inter3), .O(gate413inter10));
  nor2  gate950(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate951(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate952(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate967(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate968(.a(gate416inter0), .b(s_60), .O(gate416inter1));
  and2  gate969(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate970(.a(s_60), .O(gate416inter3));
  inv1  gate971(.a(s_61), .O(gate416inter4));
  nand2 gate972(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate973(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate974(.a(G30), .O(gate416inter7));
  inv1  gate975(.a(G1123), .O(gate416inter8));
  nand2 gate976(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate977(.a(s_61), .b(gate416inter3), .O(gate416inter10));
  nor2  gate978(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate979(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate980(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1205(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1206(.a(gate419inter0), .b(s_94), .O(gate419inter1));
  and2  gate1207(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1208(.a(s_94), .O(gate419inter3));
  inv1  gate1209(.a(s_95), .O(gate419inter4));
  nand2 gate1210(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1211(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1212(.a(G1), .O(gate419inter7));
  inv1  gate1213(.a(G1132), .O(gate419inter8));
  nand2 gate1214(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1215(.a(s_95), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1216(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1217(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1218(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1345(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1346(.a(gate421inter0), .b(s_114), .O(gate421inter1));
  and2  gate1347(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1348(.a(s_114), .O(gate421inter3));
  inv1  gate1349(.a(s_115), .O(gate421inter4));
  nand2 gate1350(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1351(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1352(.a(G2), .O(gate421inter7));
  inv1  gate1353(.a(G1135), .O(gate421inter8));
  nand2 gate1354(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1355(.a(s_115), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1356(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1357(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1358(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1247(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1248(.a(gate425inter0), .b(s_100), .O(gate425inter1));
  and2  gate1249(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1250(.a(s_100), .O(gate425inter3));
  inv1  gate1251(.a(s_101), .O(gate425inter4));
  nand2 gate1252(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1253(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1254(.a(G4), .O(gate425inter7));
  inv1  gate1255(.a(G1141), .O(gate425inter8));
  nand2 gate1256(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1257(.a(s_101), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1258(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1259(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1260(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate925(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate926(.a(gate428inter0), .b(s_54), .O(gate428inter1));
  and2  gate927(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate928(.a(s_54), .O(gate428inter3));
  inv1  gate929(.a(s_55), .O(gate428inter4));
  nand2 gate930(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate931(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate932(.a(G1048), .O(gate428inter7));
  inv1  gate933(.a(G1144), .O(gate428inter8));
  nand2 gate934(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate935(.a(s_55), .b(gate428inter3), .O(gate428inter10));
  nor2  gate936(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate937(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate938(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1359(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1360(.a(gate429inter0), .b(s_116), .O(gate429inter1));
  and2  gate1361(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1362(.a(s_116), .O(gate429inter3));
  inv1  gate1363(.a(s_117), .O(gate429inter4));
  nand2 gate1364(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1365(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1366(.a(G6), .O(gate429inter7));
  inv1  gate1367(.a(G1147), .O(gate429inter8));
  nand2 gate1368(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1369(.a(s_117), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1370(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1371(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1372(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate589(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate590(.a(gate432inter0), .b(s_6), .O(gate432inter1));
  and2  gate591(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate592(.a(s_6), .O(gate432inter3));
  inv1  gate593(.a(s_7), .O(gate432inter4));
  nand2 gate594(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate595(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate596(.a(G1054), .O(gate432inter7));
  inv1  gate597(.a(G1150), .O(gate432inter8));
  nand2 gate598(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate599(.a(s_7), .b(gate432inter3), .O(gate432inter10));
  nor2  gate600(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate601(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate602(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate953(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate954(.a(gate444inter0), .b(s_58), .O(gate444inter1));
  and2  gate955(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate956(.a(s_58), .O(gate444inter3));
  inv1  gate957(.a(s_59), .O(gate444inter4));
  nand2 gate958(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate959(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate960(.a(G1072), .O(gate444inter7));
  inv1  gate961(.a(G1168), .O(gate444inter8));
  nand2 gate962(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate963(.a(s_59), .b(gate444inter3), .O(gate444inter10));
  nor2  gate964(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate965(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate966(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1107(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1108(.a(gate454inter0), .b(s_80), .O(gate454inter1));
  and2  gate1109(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1110(.a(s_80), .O(gate454inter3));
  inv1  gate1111(.a(s_81), .O(gate454inter4));
  nand2 gate1112(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1113(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1114(.a(G1087), .O(gate454inter7));
  inv1  gate1115(.a(G1183), .O(gate454inter8));
  nand2 gate1116(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1117(.a(s_81), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1118(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1119(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1120(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate701(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate702(.a(gate456inter0), .b(s_22), .O(gate456inter1));
  and2  gate703(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate704(.a(s_22), .O(gate456inter3));
  inv1  gate705(.a(s_23), .O(gate456inter4));
  nand2 gate706(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate707(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate708(.a(G1090), .O(gate456inter7));
  inv1  gate709(.a(G1186), .O(gate456inter8));
  nand2 gate710(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate711(.a(s_23), .b(gate456inter3), .O(gate456inter10));
  nor2  gate712(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate713(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate714(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate743(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate744(.a(gate464inter0), .b(s_28), .O(gate464inter1));
  and2  gate745(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate746(.a(s_28), .O(gate464inter3));
  inv1  gate747(.a(s_29), .O(gate464inter4));
  nand2 gate748(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate749(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate750(.a(G1102), .O(gate464inter7));
  inv1  gate751(.a(G1198), .O(gate464inter8));
  nand2 gate752(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate753(.a(s_29), .b(gate464inter3), .O(gate464inter10));
  nor2  gate754(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate755(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate756(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate981(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate982(.a(gate467inter0), .b(s_62), .O(gate467inter1));
  and2  gate983(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate984(.a(s_62), .O(gate467inter3));
  inv1  gate985(.a(s_63), .O(gate467inter4));
  nand2 gate986(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate987(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate988(.a(G25), .O(gate467inter7));
  inv1  gate989(.a(G1204), .O(gate467inter8));
  nand2 gate990(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate991(.a(s_63), .b(gate467inter3), .O(gate467inter10));
  nor2  gate992(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate993(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate994(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate883(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate884(.a(gate474inter0), .b(s_48), .O(gate474inter1));
  and2  gate885(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate886(.a(s_48), .O(gate474inter3));
  inv1  gate887(.a(s_49), .O(gate474inter4));
  nand2 gate888(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate889(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate890(.a(G1117), .O(gate474inter7));
  inv1  gate891(.a(G1213), .O(gate474inter8));
  nand2 gate892(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate893(.a(s_49), .b(gate474inter3), .O(gate474inter10));
  nor2  gate894(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate895(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate896(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1219(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1220(.a(gate480inter0), .b(s_96), .O(gate480inter1));
  and2  gate1221(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1222(.a(s_96), .O(gate480inter3));
  inv1  gate1223(.a(s_97), .O(gate480inter4));
  nand2 gate1224(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1225(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1226(.a(G1126), .O(gate480inter7));
  inv1  gate1227(.a(G1222), .O(gate480inter8));
  nand2 gate1228(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1229(.a(s_97), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1230(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1231(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1232(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1191(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1192(.a(gate482inter0), .b(s_92), .O(gate482inter1));
  and2  gate1193(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1194(.a(s_92), .O(gate482inter3));
  inv1  gate1195(.a(s_93), .O(gate482inter4));
  nand2 gate1196(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1197(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1198(.a(G1129), .O(gate482inter7));
  inv1  gate1199(.a(G1225), .O(gate482inter8));
  nand2 gate1200(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1201(.a(s_93), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1202(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1203(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1204(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1387(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1388(.a(gate483inter0), .b(s_120), .O(gate483inter1));
  and2  gate1389(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1390(.a(s_120), .O(gate483inter3));
  inv1  gate1391(.a(s_121), .O(gate483inter4));
  nand2 gate1392(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1393(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1394(.a(G1228), .O(gate483inter7));
  inv1  gate1395(.a(G1229), .O(gate483inter8));
  nand2 gate1396(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1397(.a(s_121), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1398(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1399(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1400(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate729(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate730(.a(gate487inter0), .b(s_26), .O(gate487inter1));
  and2  gate731(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate732(.a(s_26), .O(gate487inter3));
  inv1  gate733(.a(s_27), .O(gate487inter4));
  nand2 gate734(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate735(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate736(.a(G1236), .O(gate487inter7));
  inv1  gate737(.a(G1237), .O(gate487inter8));
  nand2 gate738(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate739(.a(s_27), .b(gate487inter3), .O(gate487inter10));
  nor2  gate740(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate741(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate742(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1009(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1010(.a(gate489inter0), .b(s_66), .O(gate489inter1));
  and2  gate1011(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1012(.a(s_66), .O(gate489inter3));
  inv1  gate1013(.a(s_67), .O(gate489inter4));
  nand2 gate1014(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1015(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1016(.a(G1240), .O(gate489inter7));
  inv1  gate1017(.a(G1241), .O(gate489inter8));
  nand2 gate1018(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1019(.a(s_67), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1020(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1021(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1022(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate799(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate800(.a(gate495inter0), .b(s_36), .O(gate495inter1));
  and2  gate801(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate802(.a(s_36), .O(gate495inter3));
  inv1  gate803(.a(s_37), .O(gate495inter4));
  nand2 gate804(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate805(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate806(.a(G1252), .O(gate495inter7));
  inv1  gate807(.a(G1253), .O(gate495inter8));
  nand2 gate808(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate809(.a(s_37), .b(gate495inter3), .O(gate495inter10));
  nor2  gate810(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate811(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate812(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1289(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1290(.a(gate502inter0), .b(s_106), .O(gate502inter1));
  and2  gate1291(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1292(.a(s_106), .O(gate502inter3));
  inv1  gate1293(.a(s_107), .O(gate502inter4));
  nand2 gate1294(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1295(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1296(.a(G1266), .O(gate502inter7));
  inv1  gate1297(.a(G1267), .O(gate502inter8));
  nand2 gate1298(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1299(.a(s_107), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1300(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1301(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1302(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1261(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1262(.a(gate511inter0), .b(s_102), .O(gate511inter1));
  and2  gate1263(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1264(.a(s_102), .O(gate511inter3));
  inv1  gate1265(.a(s_103), .O(gate511inter4));
  nand2 gate1266(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1267(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1268(.a(G1284), .O(gate511inter7));
  inv1  gate1269(.a(G1285), .O(gate511inter8));
  nand2 gate1270(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1271(.a(s_103), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1272(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1273(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1274(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule