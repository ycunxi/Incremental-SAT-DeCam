module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate561(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate562(.a(gate11inter0), .b(s_2), .O(gate11inter1));
  and2  gate563(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate564(.a(s_2), .O(gate11inter3));
  inv1  gate565(.a(s_3), .O(gate11inter4));
  nand2 gate566(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate567(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate568(.a(G5), .O(gate11inter7));
  inv1  gate569(.a(G6), .O(gate11inter8));
  nand2 gate570(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate571(.a(s_3), .b(gate11inter3), .O(gate11inter10));
  nor2  gate572(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate573(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate574(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1093(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1094(.a(gate12inter0), .b(s_78), .O(gate12inter1));
  and2  gate1095(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1096(.a(s_78), .O(gate12inter3));
  inv1  gate1097(.a(s_79), .O(gate12inter4));
  nand2 gate1098(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1099(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1100(.a(G7), .O(gate12inter7));
  inv1  gate1101(.a(G8), .O(gate12inter8));
  nand2 gate1102(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1103(.a(s_79), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1104(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1105(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1106(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1849(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1850(.a(gate14inter0), .b(s_186), .O(gate14inter1));
  and2  gate1851(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1852(.a(s_186), .O(gate14inter3));
  inv1  gate1853(.a(s_187), .O(gate14inter4));
  nand2 gate1854(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1855(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1856(.a(G11), .O(gate14inter7));
  inv1  gate1857(.a(G12), .O(gate14inter8));
  nand2 gate1858(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1859(.a(s_187), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1860(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1861(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1862(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1667(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1668(.a(gate22inter0), .b(s_160), .O(gate22inter1));
  and2  gate1669(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1670(.a(s_160), .O(gate22inter3));
  inv1  gate1671(.a(s_161), .O(gate22inter4));
  nand2 gate1672(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1673(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1674(.a(G27), .O(gate22inter7));
  inv1  gate1675(.a(G28), .O(gate22inter8));
  nand2 gate1676(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1677(.a(s_161), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1678(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1679(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1680(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1471(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1472(.a(gate26inter0), .b(s_132), .O(gate26inter1));
  and2  gate1473(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1474(.a(s_132), .O(gate26inter3));
  inv1  gate1475(.a(s_133), .O(gate26inter4));
  nand2 gate1476(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1477(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1478(.a(G9), .O(gate26inter7));
  inv1  gate1479(.a(G13), .O(gate26inter8));
  nand2 gate1480(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1481(.a(s_133), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1482(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1483(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1484(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1051(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1052(.a(gate29inter0), .b(s_72), .O(gate29inter1));
  and2  gate1053(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1054(.a(s_72), .O(gate29inter3));
  inv1  gate1055(.a(s_73), .O(gate29inter4));
  nand2 gate1056(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1057(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1058(.a(G3), .O(gate29inter7));
  inv1  gate1059(.a(G7), .O(gate29inter8));
  nand2 gate1060(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1061(.a(s_73), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1062(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1063(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1064(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1261(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1262(.a(gate35inter0), .b(s_102), .O(gate35inter1));
  and2  gate1263(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1264(.a(s_102), .O(gate35inter3));
  inv1  gate1265(.a(s_103), .O(gate35inter4));
  nand2 gate1266(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1267(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1268(.a(G18), .O(gate35inter7));
  inv1  gate1269(.a(G22), .O(gate35inter8));
  nand2 gate1270(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1271(.a(s_103), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1272(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1273(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1274(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1121(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1122(.a(gate37inter0), .b(s_82), .O(gate37inter1));
  and2  gate1123(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1124(.a(s_82), .O(gate37inter3));
  inv1  gate1125(.a(s_83), .O(gate37inter4));
  nand2 gate1126(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1127(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1128(.a(G19), .O(gate37inter7));
  inv1  gate1129(.a(G23), .O(gate37inter8));
  nand2 gate1130(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1131(.a(s_83), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1132(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1133(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1134(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1513(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1514(.a(gate40inter0), .b(s_138), .O(gate40inter1));
  and2  gate1515(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1516(.a(s_138), .O(gate40inter3));
  inv1  gate1517(.a(s_139), .O(gate40inter4));
  nand2 gate1518(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1519(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1520(.a(G28), .O(gate40inter7));
  inv1  gate1521(.a(G32), .O(gate40inter8));
  nand2 gate1522(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1523(.a(s_139), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1524(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1525(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1526(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate645(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate646(.a(gate43inter0), .b(s_14), .O(gate43inter1));
  and2  gate647(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate648(.a(s_14), .O(gate43inter3));
  inv1  gate649(.a(s_15), .O(gate43inter4));
  nand2 gate650(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate651(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate652(.a(G3), .O(gate43inter7));
  inv1  gate653(.a(G269), .O(gate43inter8));
  nand2 gate654(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate655(.a(s_15), .b(gate43inter3), .O(gate43inter10));
  nor2  gate656(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate657(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate658(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate939(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate940(.a(gate44inter0), .b(s_56), .O(gate44inter1));
  and2  gate941(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate942(.a(s_56), .O(gate44inter3));
  inv1  gate943(.a(s_57), .O(gate44inter4));
  nand2 gate944(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate945(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate946(.a(G4), .O(gate44inter7));
  inv1  gate947(.a(G269), .O(gate44inter8));
  nand2 gate948(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate949(.a(s_57), .b(gate44inter3), .O(gate44inter10));
  nor2  gate950(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate951(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate952(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1079(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1080(.a(gate46inter0), .b(s_76), .O(gate46inter1));
  and2  gate1081(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1082(.a(s_76), .O(gate46inter3));
  inv1  gate1083(.a(s_77), .O(gate46inter4));
  nand2 gate1084(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1085(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1086(.a(G6), .O(gate46inter7));
  inv1  gate1087(.a(G272), .O(gate46inter8));
  nand2 gate1088(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1089(.a(s_77), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1090(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1091(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1092(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1779(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1780(.a(gate51inter0), .b(s_176), .O(gate51inter1));
  and2  gate1781(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1782(.a(s_176), .O(gate51inter3));
  inv1  gate1783(.a(s_177), .O(gate51inter4));
  nand2 gate1784(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1785(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1786(.a(G11), .O(gate51inter7));
  inv1  gate1787(.a(G281), .O(gate51inter8));
  nand2 gate1788(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1789(.a(s_177), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1790(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1791(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1792(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1135(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1136(.a(gate53inter0), .b(s_84), .O(gate53inter1));
  and2  gate1137(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1138(.a(s_84), .O(gate53inter3));
  inv1  gate1139(.a(s_85), .O(gate53inter4));
  nand2 gate1140(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1141(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1142(.a(G13), .O(gate53inter7));
  inv1  gate1143(.a(G284), .O(gate53inter8));
  nand2 gate1144(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1145(.a(s_85), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1146(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1147(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1148(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1583(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1584(.a(gate54inter0), .b(s_148), .O(gate54inter1));
  and2  gate1585(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1586(.a(s_148), .O(gate54inter3));
  inv1  gate1587(.a(s_149), .O(gate54inter4));
  nand2 gate1588(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1589(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1590(.a(G14), .O(gate54inter7));
  inv1  gate1591(.a(G284), .O(gate54inter8));
  nand2 gate1592(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1593(.a(s_149), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1594(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1595(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1596(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1863(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1864(.a(gate58inter0), .b(s_188), .O(gate58inter1));
  and2  gate1865(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1866(.a(s_188), .O(gate58inter3));
  inv1  gate1867(.a(s_189), .O(gate58inter4));
  nand2 gate1868(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1869(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1870(.a(G18), .O(gate58inter7));
  inv1  gate1871(.a(G290), .O(gate58inter8));
  nand2 gate1872(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1873(.a(s_189), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1874(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1875(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1876(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1289(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1290(.a(gate59inter0), .b(s_106), .O(gate59inter1));
  and2  gate1291(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1292(.a(s_106), .O(gate59inter3));
  inv1  gate1293(.a(s_107), .O(gate59inter4));
  nand2 gate1294(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1295(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1296(.a(G19), .O(gate59inter7));
  inv1  gate1297(.a(G293), .O(gate59inter8));
  nand2 gate1298(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1299(.a(s_107), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1300(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1301(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1302(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1723(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1724(.a(gate63inter0), .b(s_168), .O(gate63inter1));
  and2  gate1725(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1726(.a(s_168), .O(gate63inter3));
  inv1  gate1727(.a(s_169), .O(gate63inter4));
  nand2 gate1728(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1729(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1730(.a(G23), .O(gate63inter7));
  inv1  gate1731(.a(G299), .O(gate63inter8));
  nand2 gate1732(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1733(.a(s_169), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1734(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1735(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1736(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1709(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1710(.a(gate65inter0), .b(s_166), .O(gate65inter1));
  and2  gate1711(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1712(.a(s_166), .O(gate65inter3));
  inv1  gate1713(.a(s_167), .O(gate65inter4));
  nand2 gate1714(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1715(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1716(.a(G25), .O(gate65inter7));
  inv1  gate1717(.a(G302), .O(gate65inter8));
  nand2 gate1718(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1719(.a(s_167), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1720(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1721(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1722(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1387(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1388(.a(gate70inter0), .b(s_120), .O(gate70inter1));
  and2  gate1389(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1390(.a(s_120), .O(gate70inter3));
  inv1  gate1391(.a(s_121), .O(gate70inter4));
  nand2 gate1392(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1393(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1394(.a(G30), .O(gate70inter7));
  inv1  gate1395(.a(G308), .O(gate70inter8));
  nand2 gate1396(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1397(.a(s_121), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1398(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1399(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1400(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1037(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1038(.a(gate77inter0), .b(s_70), .O(gate77inter1));
  and2  gate1039(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1040(.a(s_70), .O(gate77inter3));
  inv1  gate1041(.a(s_71), .O(gate77inter4));
  nand2 gate1042(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1043(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1044(.a(G2), .O(gate77inter7));
  inv1  gate1045(.a(G320), .O(gate77inter8));
  nand2 gate1046(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1047(.a(s_71), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1048(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1049(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1050(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1625(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1626(.a(gate78inter0), .b(s_154), .O(gate78inter1));
  and2  gate1627(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1628(.a(s_154), .O(gate78inter3));
  inv1  gate1629(.a(s_155), .O(gate78inter4));
  nand2 gate1630(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1631(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1632(.a(G6), .O(gate78inter7));
  inv1  gate1633(.a(G320), .O(gate78inter8));
  nand2 gate1634(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1635(.a(s_155), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1636(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1637(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1638(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate799(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate800(.a(gate82inter0), .b(s_36), .O(gate82inter1));
  and2  gate801(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate802(.a(s_36), .O(gate82inter3));
  inv1  gate803(.a(s_37), .O(gate82inter4));
  nand2 gate804(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate805(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate806(.a(G7), .O(gate82inter7));
  inv1  gate807(.a(G326), .O(gate82inter8));
  nand2 gate808(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate809(.a(s_37), .b(gate82inter3), .O(gate82inter10));
  nor2  gate810(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate811(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate812(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1765(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1766(.a(gate90inter0), .b(s_174), .O(gate90inter1));
  and2  gate1767(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1768(.a(s_174), .O(gate90inter3));
  inv1  gate1769(.a(s_175), .O(gate90inter4));
  nand2 gate1770(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1771(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1772(.a(G21), .O(gate90inter7));
  inv1  gate1773(.a(G338), .O(gate90inter8));
  nand2 gate1774(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1775(.a(s_175), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1776(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1777(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1778(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1149(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1150(.a(gate91inter0), .b(s_86), .O(gate91inter1));
  and2  gate1151(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1152(.a(s_86), .O(gate91inter3));
  inv1  gate1153(.a(s_87), .O(gate91inter4));
  nand2 gate1154(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1155(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1156(.a(G25), .O(gate91inter7));
  inv1  gate1157(.a(G341), .O(gate91inter8));
  nand2 gate1158(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1159(.a(s_87), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1160(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1161(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1162(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1065(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1066(.a(gate96inter0), .b(s_74), .O(gate96inter1));
  and2  gate1067(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1068(.a(s_74), .O(gate96inter3));
  inv1  gate1069(.a(s_75), .O(gate96inter4));
  nand2 gate1070(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1071(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1072(.a(G30), .O(gate96inter7));
  inv1  gate1073(.a(G347), .O(gate96inter8));
  nand2 gate1074(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1075(.a(s_75), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1076(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1077(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1078(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate603(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate604(.a(gate97inter0), .b(s_8), .O(gate97inter1));
  and2  gate605(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate606(.a(s_8), .O(gate97inter3));
  inv1  gate607(.a(s_9), .O(gate97inter4));
  nand2 gate608(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate609(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate610(.a(G19), .O(gate97inter7));
  inv1  gate611(.a(G350), .O(gate97inter8));
  nand2 gate612(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate613(.a(s_9), .b(gate97inter3), .O(gate97inter10));
  nor2  gate614(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate615(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate616(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate897(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate898(.a(gate102inter0), .b(s_50), .O(gate102inter1));
  and2  gate899(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate900(.a(s_50), .O(gate102inter3));
  inv1  gate901(.a(s_51), .O(gate102inter4));
  nand2 gate902(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate903(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate904(.a(G24), .O(gate102inter7));
  inv1  gate905(.a(G356), .O(gate102inter8));
  nand2 gate906(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate907(.a(s_51), .b(gate102inter3), .O(gate102inter10));
  nor2  gate908(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate909(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate910(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1611(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1612(.a(gate106inter0), .b(s_152), .O(gate106inter1));
  and2  gate1613(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1614(.a(s_152), .O(gate106inter3));
  inv1  gate1615(.a(s_153), .O(gate106inter4));
  nand2 gate1616(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1617(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1618(.a(G364), .O(gate106inter7));
  inv1  gate1619(.a(G365), .O(gate106inter8));
  nand2 gate1620(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1621(.a(s_153), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1622(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1623(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1624(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate589(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate590(.a(gate107inter0), .b(s_6), .O(gate107inter1));
  and2  gate591(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate592(.a(s_6), .O(gate107inter3));
  inv1  gate593(.a(s_7), .O(gate107inter4));
  nand2 gate594(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate595(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate596(.a(G366), .O(gate107inter7));
  inv1  gate597(.a(G367), .O(gate107inter8));
  nand2 gate598(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate599(.a(s_7), .b(gate107inter3), .O(gate107inter10));
  nor2  gate600(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate601(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate602(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate771(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate772(.a(gate108inter0), .b(s_32), .O(gate108inter1));
  and2  gate773(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate774(.a(s_32), .O(gate108inter3));
  inv1  gate775(.a(s_33), .O(gate108inter4));
  nand2 gate776(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate777(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate778(.a(G368), .O(gate108inter7));
  inv1  gate779(.a(G369), .O(gate108inter8));
  nand2 gate780(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate781(.a(s_33), .b(gate108inter3), .O(gate108inter10));
  nor2  gate782(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate783(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate784(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate813(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate814(.a(gate115inter0), .b(s_38), .O(gate115inter1));
  and2  gate815(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate816(.a(s_38), .O(gate115inter3));
  inv1  gate817(.a(s_39), .O(gate115inter4));
  nand2 gate818(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate819(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate820(.a(G382), .O(gate115inter7));
  inv1  gate821(.a(G383), .O(gate115inter8));
  nand2 gate822(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate823(.a(s_39), .b(gate115inter3), .O(gate115inter10));
  nor2  gate824(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate825(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate826(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate715(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate716(.a(gate117inter0), .b(s_24), .O(gate117inter1));
  and2  gate717(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate718(.a(s_24), .O(gate117inter3));
  inv1  gate719(.a(s_25), .O(gate117inter4));
  nand2 gate720(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate721(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate722(.a(G386), .O(gate117inter7));
  inv1  gate723(.a(G387), .O(gate117inter8));
  nand2 gate724(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate725(.a(s_25), .b(gate117inter3), .O(gate117inter10));
  nor2  gate726(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate727(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate728(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1107(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1108(.a(gate119inter0), .b(s_80), .O(gate119inter1));
  and2  gate1109(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1110(.a(s_80), .O(gate119inter3));
  inv1  gate1111(.a(s_81), .O(gate119inter4));
  nand2 gate1112(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1113(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1114(.a(G390), .O(gate119inter7));
  inv1  gate1115(.a(G391), .O(gate119inter8));
  nand2 gate1116(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1117(.a(s_81), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1118(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1119(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1120(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate757(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate758(.a(gate122inter0), .b(s_30), .O(gate122inter1));
  and2  gate759(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate760(.a(s_30), .O(gate122inter3));
  inv1  gate761(.a(s_31), .O(gate122inter4));
  nand2 gate762(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate763(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate764(.a(G396), .O(gate122inter7));
  inv1  gate765(.a(G397), .O(gate122inter8));
  nand2 gate766(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate767(.a(s_31), .b(gate122inter3), .O(gate122inter10));
  nor2  gate768(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate769(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate770(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate827(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate828(.a(gate124inter0), .b(s_40), .O(gate124inter1));
  and2  gate829(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate830(.a(s_40), .O(gate124inter3));
  inv1  gate831(.a(s_41), .O(gate124inter4));
  nand2 gate832(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate833(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate834(.a(G400), .O(gate124inter7));
  inv1  gate835(.a(G401), .O(gate124inter8));
  nand2 gate836(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate837(.a(s_41), .b(gate124inter3), .O(gate124inter10));
  nor2  gate838(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate839(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate840(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate547(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate548(.a(gate126inter0), .b(s_0), .O(gate126inter1));
  and2  gate549(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate550(.a(s_0), .O(gate126inter3));
  inv1  gate551(.a(s_1), .O(gate126inter4));
  nand2 gate552(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate553(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate554(.a(G404), .O(gate126inter7));
  inv1  gate555(.a(G405), .O(gate126inter8));
  nand2 gate556(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate557(.a(s_1), .b(gate126inter3), .O(gate126inter10));
  nor2  gate558(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate559(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate560(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate729(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate730(.a(gate128inter0), .b(s_26), .O(gate128inter1));
  and2  gate731(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate732(.a(s_26), .O(gate128inter3));
  inv1  gate733(.a(s_27), .O(gate128inter4));
  nand2 gate734(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate735(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate736(.a(G408), .O(gate128inter7));
  inv1  gate737(.a(G409), .O(gate128inter8));
  nand2 gate738(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate739(.a(s_27), .b(gate128inter3), .O(gate128inter10));
  nor2  gate740(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate741(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate742(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1457(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1458(.a(gate131inter0), .b(s_130), .O(gate131inter1));
  and2  gate1459(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1460(.a(s_130), .O(gate131inter3));
  inv1  gate1461(.a(s_131), .O(gate131inter4));
  nand2 gate1462(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1463(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1464(.a(G414), .O(gate131inter7));
  inv1  gate1465(.a(G415), .O(gate131inter8));
  nand2 gate1466(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1467(.a(s_131), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1468(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1469(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1470(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate855(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate856(.a(gate134inter0), .b(s_44), .O(gate134inter1));
  and2  gate857(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate858(.a(s_44), .O(gate134inter3));
  inv1  gate859(.a(s_45), .O(gate134inter4));
  nand2 gate860(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate861(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate862(.a(G420), .O(gate134inter7));
  inv1  gate863(.a(G421), .O(gate134inter8));
  nand2 gate864(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate865(.a(s_45), .b(gate134inter3), .O(gate134inter10));
  nor2  gate866(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate867(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate868(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate911(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate912(.a(gate144inter0), .b(s_52), .O(gate144inter1));
  and2  gate913(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate914(.a(s_52), .O(gate144inter3));
  inv1  gate915(.a(s_53), .O(gate144inter4));
  nand2 gate916(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate917(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate918(.a(G468), .O(gate144inter7));
  inv1  gate919(.a(G471), .O(gate144inter8));
  nand2 gate920(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate921(.a(s_53), .b(gate144inter3), .O(gate144inter10));
  nor2  gate922(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate923(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate924(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1555(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1556(.a(gate145inter0), .b(s_144), .O(gate145inter1));
  and2  gate1557(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1558(.a(s_144), .O(gate145inter3));
  inv1  gate1559(.a(s_145), .O(gate145inter4));
  nand2 gate1560(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1561(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1562(.a(G474), .O(gate145inter7));
  inv1  gate1563(.a(G477), .O(gate145inter8));
  nand2 gate1564(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1565(.a(s_145), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1566(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1567(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1568(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate659(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate660(.a(gate153inter0), .b(s_16), .O(gate153inter1));
  and2  gate661(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate662(.a(s_16), .O(gate153inter3));
  inv1  gate663(.a(s_17), .O(gate153inter4));
  nand2 gate664(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate665(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate666(.a(G426), .O(gate153inter7));
  inv1  gate667(.a(G522), .O(gate153inter8));
  nand2 gate668(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate669(.a(s_17), .b(gate153inter3), .O(gate153inter10));
  nor2  gate670(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate671(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate672(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1359(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1360(.a(gate156inter0), .b(s_116), .O(gate156inter1));
  and2  gate1361(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1362(.a(s_116), .O(gate156inter3));
  inv1  gate1363(.a(s_117), .O(gate156inter4));
  nand2 gate1364(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1365(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1366(.a(G435), .O(gate156inter7));
  inv1  gate1367(.a(G525), .O(gate156inter8));
  nand2 gate1368(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1369(.a(s_117), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1370(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1371(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1372(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1303(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1304(.a(gate158inter0), .b(s_108), .O(gate158inter1));
  and2  gate1305(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1306(.a(s_108), .O(gate158inter3));
  inv1  gate1307(.a(s_109), .O(gate158inter4));
  nand2 gate1308(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1309(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1310(.a(G441), .O(gate158inter7));
  inv1  gate1311(.a(G528), .O(gate158inter8));
  nand2 gate1312(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1313(.a(s_109), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1314(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1315(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1316(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate673(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate674(.a(gate172inter0), .b(s_18), .O(gate172inter1));
  and2  gate675(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate676(.a(s_18), .O(gate172inter3));
  inv1  gate677(.a(s_19), .O(gate172inter4));
  nand2 gate678(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate679(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate680(.a(G483), .O(gate172inter7));
  inv1  gate681(.a(G549), .O(gate172inter8));
  nand2 gate682(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate683(.a(s_19), .b(gate172inter3), .O(gate172inter10));
  nor2  gate684(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate685(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate686(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1345(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1346(.a(gate175inter0), .b(s_114), .O(gate175inter1));
  and2  gate1347(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1348(.a(s_114), .O(gate175inter3));
  inv1  gate1349(.a(s_115), .O(gate175inter4));
  nand2 gate1350(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1351(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1352(.a(G492), .O(gate175inter7));
  inv1  gate1353(.a(G555), .O(gate175inter8));
  nand2 gate1354(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1355(.a(s_115), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1356(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1357(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1358(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1835(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1836(.a(gate176inter0), .b(s_184), .O(gate176inter1));
  and2  gate1837(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1838(.a(s_184), .O(gate176inter3));
  inv1  gate1839(.a(s_185), .O(gate176inter4));
  nand2 gate1840(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1841(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1842(.a(G495), .O(gate176inter7));
  inv1  gate1843(.a(G555), .O(gate176inter8));
  nand2 gate1844(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1845(.a(s_185), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1846(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1847(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1848(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate743(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate744(.a(gate182inter0), .b(s_28), .O(gate182inter1));
  and2  gate745(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate746(.a(s_28), .O(gate182inter3));
  inv1  gate747(.a(s_29), .O(gate182inter4));
  nand2 gate748(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate749(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate750(.a(G513), .O(gate182inter7));
  inv1  gate751(.a(G564), .O(gate182inter8));
  nand2 gate752(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate753(.a(s_29), .b(gate182inter3), .O(gate182inter10));
  nor2  gate754(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate755(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate756(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1317(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1318(.a(gate190inter0), .b(s_110), .O(gate190inter1));
  and2  gate1319(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1320(.a(s_110), .O(gate190inter3));
  inv1  gate1321(.a(s_111), .O(gate190inter4));
  nand2 gate1322(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1323(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1324(.a(G580), .O(gate190inter7));
  inv1  gate1325(.a(G581), .O(gate190inter8));
  nand2 gate1326(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1327(.a(s_111), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1328(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1329(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1330(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1247(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1248(.a(gate197inter0), .b(s_100), .O(gate197inter1));
  and2  gate1249(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1250(.a(s_100), .O(gate197inter3));
  inv1  gate1251(.a(s_101), .O(gate197inter4));
  nand2 gate1252(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1253(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1254(.a(G594), .O(gate197inter7));
  inv1  gate1255(.a(G595), .O(gate197inter8));
  nand2 gate1256(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1257(.a(s_101), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1258(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1259(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1260(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate631(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate632(.a(gate198inter0), .b(s_12), .O(gate198inter1));
  and2  gate633(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate634(.a(s_12), .O(gate198inter3));
  inv1  gate635(.a(s_13), .O(gate198inter4));
  nand2 gate636(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate637(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate638(.a(G596), .O(gate198inter7));
  inv1  gate639(.a(G597), .O(gate198inter8));
  nand2 gate640(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate641(.a(s_13), .b(gate198inter3), .O(gate198inter10));
  nor2  gate642(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate643(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate644(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1191(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1192(.a(gate199inter0), .b(s_92), .O(gate199inter1));
  and2  gate1193(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1194(.a(s_92), .O(gate199inter3));
  inv1  gate1195(.a(s_93), .O(gate199inter4));
  nand2 gate1196(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1197(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1198(.a(G598), .O(gate199inter7));
  inv1  gate1199(.a(G599), .O(gate199inter8));
  nand2 gate1200(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1201(.a(s_93), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1202(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1203(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1204(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1205(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1206(.a(gate209inter0), .b(s_94), .O(gate209inter1));
  and2  gate1207(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1208(.a(s_94), .O(gate209inter3));
  inv1  gate1209(.a(s_95), .O(gate209inter4));
  nand2 gate1210(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1211(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1212(.a(G602), .O(gate209inter7));
  inv1  gate1213(.a(G666), .O(gate209inter8));
  nand2 gate1214(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1215(.a(s_95), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1216(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1217(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1218(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1541(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1542(.a(gate236inter0), .b(s_142), .O(gate236inter1));
  and2  gate1543(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1544(.a(s_142), .O(gate236inter3));
  inv1  gate1545(.a(s_143), .O(gate236inter4));
  nand2 gate1546(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1547(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1548(.a(G251), .O(gate236inter7));
  inv1  gate1549(.a(G727), .O(gate236inter8));
  nand2 gate1550(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1551(.a(s_143), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1552(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1553(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1554(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1275(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1276(.a(gate249inter0), .b(s_104), .O(gate249inter1));
  and2  gate1277(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1278(.a(s_104), .O(gate249inter3));
  inv1  gate1279(.a(s_105), .O(gate249inter4));
  nand2 gate1280(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1281(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1282(.a(G254), .O(gate249inter7));
  inv1  gate1283(.a(G742), .O(gate249inter8));
  nand2 gate1284(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1285(.a(s_105), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1286(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1287(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1288(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1653(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1654(.a(gate250inter0), .b(s_158), .O(gate250inter1));
  and2  gate1655(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1656(.a(s_158), .O(gate250inter3));
  inv1  gate1657(.a(s_159), .O(gate250inter4));
  nand2 gate1658(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1659(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1660(.a(G706), .O(gate250inter7));
  inv1  gate1661(.a(G742), .O(gate250inter8));
  nand2 gate1662(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1663(.a(s_159), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1664(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1665(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1666(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1373(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1374(.a(gate255inter0), .b(s_118), .O(gate255inter1));
  and2  gate1375(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1376(.a(s_118), .O(gate255inter3));
  inv1  gate1377(.a(s_119), .O(gate255inter4));
  nand2 gate1378(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1379(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1380(.a(G263), .O(gate255inter7));
  inv1  gate1381(.a(G751), .O(gate255inter8));
  nand2 gate1382(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1383(.a(s_119), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1384(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1385(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1386(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1681(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1682(.a(gate257inter0), .b(s_162), .O(gate257inter1));
  and2  gate1683(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1684(.a(s_162), .O(gate257inter3));
  inv1  gate1685(.a(s_163), .O(gate257inter4));
  nand2 gate1686(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1687(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1688(.a(G754), .O(gate257inter7));
  inv1  gate1689(.a(G755), .O(gate257inter8));
  nand2 gate1690(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1691(.a(s_163), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1692(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1693(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1694(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1415(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1416(.a(gate268inter0), .b(s_124), .O(gate268inter1));
  and2  gate1417(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1418(.a(s_124), .O(gate268inter3));
  inv1  gate1419(.a(s_125), .O(gate268inter4));
  nand2 gate1420(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1421(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1422(.a(G651), .O(gate268inter7));
  inv1  gate1423(.a(G779), .O(gate268inter8));
  nand2 gate1424(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1425(.a(s_125), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1426(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1427(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1428(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1695(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1696(.a(gate272inter0), .b(s_164), .O(gate272inter1));
  and2  gate1697(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1698(.a(s_164), .O(gate272inter3));
  inv1  gate1699(.a(s_165), .O(gate272inter4));
  nand2 gate1700(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1701(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1702(.a(G663), .O(gate272inter7));
  inv1  gate1703(.a(G791), .O(gate272inter8));
  nand2 gate1704(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1705(.a(s_165), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1706(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1707(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1708(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1429(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1430(.a(gate275inter0), .b(s_126), .O(gate275inter1));
  and2  gate1431(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1432(.a(s_126), .O(gate275inter3));
  inv1  gate1433(.a(s_127), .O(gate275inter4));
  nand2 gate1434(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1435(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1436(.a(G645), .O(gate275inter7));
  inv1  gate1437(.a(G797), .O(gate275inter8));
  nand2 gate1438(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1439(.a(s_127), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1440(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1441(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1442(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate785(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate786(.a(gate279inter0), .b(s_34), .O(gate279inter1));
  and2  gate787(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate788(.a(s_34), .O(gate279inter3));
  inv1  gate789(.a(s_35), .O(gate279inter4));
  nand2 gate790(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate791(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate792(.a(G651), .O(gate279inter7));
  inv1  gate793(.a(G803), .O(gate279inter8));
  nand2 gate794(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate795(.a(s_35), .b(gate279inter3), .O(gate279inter10));
  nor2  gate796(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate797(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate798(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1639(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1640(.a(gate283inter0), .b(s_156), .O(gate283inter1));
  and2  gate1641(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1642(.a(s_156), .O(gate283inter3));
  inv1  gate1643(.a(s_157), .O(gate283inter4));
  nand2 gate1644(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1645(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1646(.a(G657), .O(gate283inter7));
  inv1  gate1647(.a(G809), .O(gate283inter8));
  nand2 gate1648(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1649(.a(s_157), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1650(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1651(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1652(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1751(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1752(.a(gate284inter0), .b(s_172), .O(gate284inter1));
  and2  gate1753(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1754(.a(s_172), .O(gate284inter3));
  inv1  gate1755(.a(s_173), .O(gate284inter4));
  nand2 gate1756(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1757(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1758(.a(G785), .O(gate284inter7));
  inv1  gate1759(.a(G809), .O(gate284inter8));
  nand2 gate1760(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1761(.a(s_173), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1762(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1763(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1764(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate617(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate618(.a(gate285inter0), .b(s_10), .O(gate285inter1));
  and2  gate619(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate620(.a(s_10), .O(gate285inter3));
  inv1  gate621(.a(s_11), .O(gate285inter4));
  nand2 gate622(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate623(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate624(.a(G660), .O(gate285inter7));
  inv1  gate625(.a(G812), .O(gate285inter8));
  nand2 gate626(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate627(.a(s_11), .b(gate285inter3), .O(gate285inter10));
  nor2  gate628(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate629(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate630(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate953(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate954(.a(gate288inter0), .b(s_58), .O(gate288inter1));
  and2  gate955(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate956(.a(s_58), .O(gate288inter3));
  inv1  gate957(.a(s_59), .O(gate288inter4));
  nand2 gate958(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate959(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate960(.a(G791), .O(gate288inter7));
  inv1  gate961(.a(G815), .O(gate288inter8));
  nand2 gate962(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate963(.a(s_59), .b(gate288inter3), .O(gate288inter10));
  nor2  gate964(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate965(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate966(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate925(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate926(.a(gate391inter0), .b(s_54), .O(gate391inter1));
  and2  gate927(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate928(.a(s_54), .O(gate391inter3));
  inv1  gate929(.a(s_55), .O(gate391inter4));
  nand2 gate930(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate931(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate932(.a(G5), .O(gate391inter7));
  inv1  gate933(.a(G1048), .O(gate391inter8));
  nand2 gate934(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate935(.a(s_55), .b(gate391inter3), .O(gate391inter10));
  nor2  gate936(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate937(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate938(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1821(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1822(.a(gate395inter0), .b(s_182), .O(gate395inter1));
  and2  gate1823(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1824(.a(s_182), .O(gate395inter3));
  inv1  gate1825(.a(s_183), .O(gate395inter4));
  nand2 gate1826(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1827(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1828(.a(G9), .O(gate395inter7));
  inv1  gate1829(.a(G1060), .O(gate395inter8));
  nand2 gate1830(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1831(.a(s_183), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1832(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1833(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1834(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1569(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1570(.a(gate397inter0), .b(s_146), .O(gate397inter1));
  and2  gate1571(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1572(.a(s_146), .O(gate397inter3));
  inv1  gate1573(.a(s_147), .O(gate397inter4));
  nand2 gate1574(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1575(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1576(.a(G11), .O(gate397inter7));
  inv1  gate1577(.a(G1066), .O(gate397inter8));
  nand2 gate1578(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1579(.a(s_147), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1580(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1581(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1582(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1009(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1010(.a(gate403inter0), .b(s_66), .O(gate403inter1));
  and2  gate1011(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1012(.a(s_66), .O(gate403inter3));
  inv1  gate1013(.a(s_67), .O(gate403inter4));
  nand2 gate1014(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1015(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1016(.a(G17), .O(gate403inter7));
  inv1  gate1017(.a(G1084), .O(gate403inter8));
  nand2 gate1018(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1019(.a(s_67), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1020(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1021(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1022(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1737(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1738(.a(gate406inter0), .b(s_170), .O(gate406inter1));
  and2  gate1739(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1740(.a(s_170), .O(gate406inter3));
  inv1  gate1741(.a(s_171), .O(gate406inter4));
  nand2 gate1742(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1743(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1744(.a(G20), .O(gate406inter7));
  inv1  gate1745(.a(G1093), .O(gate406inter8));
  nand2 gate1746(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1747(.a(s_171), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1748(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1749(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1750(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate981(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate982(.a(gate410inter0), .b(s_62), .O(gate410inter1));
  and2  gate983(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate984(.a(s_62), .O(gate410inter3));
  inv1  gate985(.a(s_63), .O(gate410inter4));
  nand2 gate986(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate987(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate988(.a(G24), .O(gate410inter7));
  inv1  gate989(.a(G1105), .O(gate410inter8));
  nand2 gate990(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate991(.a(s_63), .b(gate410inter3), .O(gate410inter10));
  nor2  gate992(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate993(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate994(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate967(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate968(.a(gate414inter0), .b(s_60), .O(gate414inter1));
  and2  gate969(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate970(.a(s_60), .O(gate414inter3));
  inv1  gate971(.a(s_61), .O(gate414inter4));
  nand2 gate972(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate973(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate974(.a(G28), .O(gate414inter7));
  inv1  gate975(.a(G1117), .O(gate414inter8));
  nand2 gate976(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate977(.a(s_61), .b(gate414inter3), .O(gate414inter10));
  nor2  gate978(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate979(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate980(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1331(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1332(.a(gate416inter0), .b(s_112), .O(gate416inter1));
  and2  gate1333(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1334(.a(s_112), .O(gate416inter3));
  inv1  gate1335(.a(s_113), .O(gate416inter4));
  nand2 gate1336(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1337(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1338(.a(G30), .O(gate416inter7));
  inv1  gate1339(.a(G1123), .O(gate416inter8));
  nand2 gate1340(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1341(.a(s_113), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1342(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1343(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1344(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1485(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1486(.a(gate417inter0), .b(s_134), .O(gate417inter1));
  and2  gate1487(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1488(.a(s_134), .O(gate417inter3));
  inv1  gate1489(.a(s_135), .O(gate417inter4));
  nand2 gate1490(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1491(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1492(.a(G31), .O(gate417inter7));
  inv1  gate1493(.a(G1126), .O(gate417inter8));
  nand2 gate1494(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1495(.a(s_135), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1496(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1497(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1498(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate841(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate842(.a(gate419inter0), .b(s_42), .O(gate419inter1));
  and2  gate843(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate844(.a(s_42), .O(gate419inter3));
  inv1  gate845(.a(s_43), .O(gate419inter4));
  nand2 gate846(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate847(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate848(.a(G1), .O(gate419inter7));
  inv1  gate849(.a(G1132), .O(gate419inter8));
  nand2 gate850(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate851(.a(s_43), .b(gate419inter3), .O(gate419inter10));
  nor2  gate852(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate853(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate854(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1233(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1234(.a(gate424inter0), .b(s_98), .O(gate424inter1));
  and2  gate1235(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1236(.a(s_98), .O(gate424inter3));
  inv1  gate1237(.a(s_99), .O(gate424inter4));
  nand2 gate1238(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1239(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1240(.a(G1042), .O(gate424inter7));
  inv1  gate1241(.a(G1138), .O(gate424inter8));
  nand2 gate1242(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1243(.a(s_99), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1244(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1245(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1246(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate869(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate870(.a(gate426inter0), .b(s_46), .O(gate426inter1));
  and2  gate871(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate872(.a(s_46), .O(gate426inter3));
  inv1  gate873(.a(s_47), .O(gate426inter4));
  nand2 gate874(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate875(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate876(.a(G1045), .O(gate426inter7));
  inv1  gate877(.a(G1141), .O(gate426inter8));
  nand2 gate878(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate879(.a(s_47), .b(gate426inter3), .O(gate426inter10));
  nor2  gate880(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate881(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate882(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1793(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1794(.a(gate432inter0), .b(s_178), .O(gate432inter1));
  and2  gate1795(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1796(.a(s_178), .O(gate432inter3));
  inv1  gate1797(.a(s_179), .O(gate432inter4));
  nand2 gate1798(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1799(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1800(.a(G1054), .O(gate432inter7));
  inv1  gate1801(.a(G1150), .O(gate432inter8));
  nand2 gate1802(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1803(.a(s_179), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1804(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1805(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1806(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate701(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate702(.a(gate438inter0), .b(s_22), .O(gate438inter1));
  and2  gate703(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate704(.a(s_22), .O(gate438inter3));
  inv1  gate705(.a(s_23), .O(gate438inter4));
  nand2 gate706(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate707(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate708(.a(G1063), .O(gate438inter7));
  inv1  gate709(.a(G1159), .O(gate438inter8));
  nand2 gate710(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate711(.a(s_23), .b(gate438inter3), .O(gate438inter10));
  nor2  gate712(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate713(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate714(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate883(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate884(.a(gate441inter0), .b(s_48), .O(gate441inter1));
  and2  gate885(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate886(.a(s_48), .O(gate441inter3));
  inv1  gate887(.a(s_49), .O(gate441inter4));
  nand2 gate888(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate889(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate890(.a(G12), .O(gate441inter7));
  inv1  gate891(.a(G1165), .O(gate441inter8));
  nand2 gate892(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate893(.a(s_49), .b(gate441inter3), .O(gate441inter10));
  nor2  gate894(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate895(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate896(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1219(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1220(.a(gate442inter0), .b(s_96), .O(gate442inter1));
  and2  gate1221(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1222(.a(s_96), .O(gate442inter3));
  inv1  gate1223(.a(s_97), .O(gate442inter4));
  nand2 gate1224(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1225(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1226(.a(G1069), .O(gate442inter7));
  inv1  gate1227(.a(G1165), .O(gate442inter8));
  nand2 gate1228(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1229(.a(s_97), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1230(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1231(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1232(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1877(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1878(.a(gate446inter0), .b(s_190), .O(gate446inter1));
  and2  gate1879(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1880(.a(s_190), .O(gate446inter3));
  inv1  gate1881(.a(s_191), .O(gate446inter4));
  nand2 gate1882(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1883(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1884(.a(G1075), .O(gate446inter7));
  inv1  gate1885(.a(G1171), .O(gate446inter8));
  nand2 gate1886(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1887(.a(s_191), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1888(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1889(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1890(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1443(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1444(.a(gate447inter0), .b(s_128), .O(gate447inter1));
  and2  gate1445(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1446(.a(s_128), .O(gate447inter3));
  inv1  gate1447(.a(s_129), .O(gate447inter4));
  nand2 gate1448(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1449(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1450(.a(G15), .O(gate447inter7));
  inv1  gate1451(.a(G1174), .O(gate447inter8));
  nand2 gate1452(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1453(.a(s_129), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1454(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1455(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1456(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate995(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate996(.a(gate455inter0), .b(s_64), .O(gate455inter1));
  and2  gate997(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate998(.a(s_64), .O(gate455inter3));
  inv1  gate999(.a(s_65), .O(gate455inter4));
  nand2 gate1000(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1001(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1002(.a(G19), .O(gate455inter7));
  inv1  gate1003(.a(G1186), .O(gate455inter8));
  nand2 gate1004(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1005(.a(s_65), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1006(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1007(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1008(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate687(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate688(.a(gate460inter0), .b(s_20), .O(gate460inter1));
  and2  gate689(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate690(.a(s_20), .O(gate460inter3));
  inv1  gate691(.a(s_21), .O(gate460inter4));
  nand2 gate692(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate693(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate694(.a(G1096), .O(gate460inter7));
  inv1  gate695(.a(G1192), .O(gate460inter8));
  nand2 gate696(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate697(.a(s_21), .b(gate460inter3), .O(gate460inter10));
  nor2  gate698(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate699(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate700(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate1807(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1808(.a(gate461inter0), .b(s_180), .O(gate461inter1));
  and2  gate1809(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1810(.a(s_180), .O(gate461inter3));
  inv1  gate1811(.a(s_181), .O(gate461inter4));
  nand2 gate1812(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1813(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1814(.a(G22), .O(gate461inter7));
  inv1  gate1815(.a(G1195), .O(gate461inter8));
  nand2 gate1816(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1817(.a(s_181), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1818(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1819(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1820(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1401(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1402(.a(gate472inter0), .b(s_122), .O(gate472inter1));
  and2  gate1403(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1404(.a(s_122), .O(gate472inter3));
  inv1  gate1405(.a(s_123), .O(gate472inter4));
  nand2 gate1406(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1407(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1408(.a(G1114), .O(gate472inter7));
  inv1  gate1409(.a(G1210), .O(gate472inter8));
  nand2 gate1410(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1411(.a(s_123), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1412(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1413(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1414(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1597(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1598(.a(gate480inter0), .b(s_150), .O(gate480inter1));
  and2  gate1599(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1600(.a(s_150), .O(gate480inter3));
  inv1  gate1601(.a(s_151), .O(gate480inter4));
  nand2 gate1602(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1603(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1604(.a(G1126), .O(gate480inter7));
  inv1  gate1605(.a(G1222), .O(gate480inter8));
  nand2 gate1606(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1607(.a(s_151), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1608(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1609(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1610(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1023(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1024(.a(gate483inter0), .b(s_68), .O(gate483inter1));
  and2  gate1025(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1026(.a(s_68), .O(gate483inter3));
  inv1  gate1027(.a(s_69), .O(gate483inter4));
  nand2 gate1028(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1029(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1030(.a(G1228), .O(gate483inter7));
  inv1  gate1031(.a(G1229), .O(gate483inter8));
  nand2 gate1032(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1033(.a(s_69), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1034(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1035(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1036(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate575(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate576(.a(gate497inter0), .b(s_4), .O(gate497inter1));
  and2  gate577(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate578(.a(s_4), .O(gate497inter3));
  inv1  gate579(.a(s_5), .O(gate497inter4));
  nand2 gate580(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate581(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate582(.a(G1256), .O(gate497inter7));
  inv1  gate583(.a(G1257), .O(gate497inter8));
  nand2 gate584(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate585(.a(s_5), .b(gate497inter3), .O(gate497inter10));
  nor2  gate586(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate587(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate588(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1177(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1178(.a(gate504inter0), .b(s_90), .O(gate504inter1));
  and2  gate1179(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1180(.a(s_90), .O(gate504inter3));
  inv1  gate1181(.a(s_91), .O(gate504inter4));
  nand2 gate1182(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1183(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1184(.a(G1270), .O(gate504inter7));
  inv1  gate1185(.a(G1271), .O(gate504inter8));
  nand2 gate1186(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1187(.a(s_91), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1188(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1189(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1190(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1163(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1164(.a(gate507inter0), .b(s_88), .O(gate507inter1));
  and2  gate1165(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1166(.a(s_88), .O(gate507inter3));
  inv1  gate1167(.a(s_89), .O(gate507inter4));
  nand2 gate1168(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1169(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1170(.a(G1276), .O(gate507inter7));
  inv1  gate1171(.a(G1277), .O(gate507inter8));
  nand2 gate1172(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1173(.a(s_89), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1174(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1175(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1176(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1527(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1528(.a(gate508inter0), .b(s_140), .O(gate508inter1));
  and2  gate1529(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1530(.a(s_140), .O(gate508inter3));
  inv1  gate1531(.a(s_141), .O(gate508inter4));
  nand2 gate1532(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1533(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1534(.a(G1278), .O(gate508inter7));
  inv1  gate1535(.a(G1279), .O(gate508inter8));
  nand2 gate1536(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1537(.a(s_141), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1538(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1539(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1540(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1499(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1500(.a(gate512inter0), .b(s_136), .O(gate512inter1));
  and2  gate1501(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1502(.a(s_136), .O(gate512inter3));
  inv1  gate1503(.a(s_137), .O(gate512inter4));
  nand2 gate1504(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1505(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1506(.a(G1286), .O(gate512inter7));
  inv1  gate1507(.a(G1287), .O(gate512inter8));
  nand2 gate1508(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1509(.a(s_137), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1510(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1511(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1512(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule