module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate385inter0, gate385inter1, gate385inter2, gate385inter3, gate385inter4, gate385inter5, gate385inter6, gate385inter7, gate385inter8, gate385inter9, gate385inter10, gate385inter11, gate385inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate851inter0, gate851inter1, gate851inter2, gate851inter3, gate851inter4, gate851inter5, gate851inter6, gate851inter7, gate851inter8, gate851inter9, gate851inter10, gate851inter11, gate851inter12, gate760inter0, gate760inter1, gate760inter2, gate760inter3, gate760inter4, gate760inter5, gate760inter6, gate760inter7, gate760inter8, gate760inter9, gate760inter10, gate760inter11, gate760inter12, gate618inter0, gate618inter1, gate618inter2, gate618inter3, gate618inter4, gate618inter5, gate618inter6, gate618inter7, gate618inter8, gate618inter9, gate618inter10, gate618inter11, gate618inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate679inter0, gate679inter1, gate679inter2, gate679inter3, gate679inter4, gate679inter5, gate679inter6, gate679inter7, gate679inter8, gate679inter9, gate679inter10, gate679inter11, gate679inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate762inter0, gate762inter1, gate762inter2, gate762inter3, gate762inter4, gate762inter5, gate762inter6, gate762inter7, gate762inter8, gate762inter9, gate762inter10, gate762inter11, gate762inter12, gate824inter0, gate824inter1, gate824inter2, gate824inter3, gate824inter4, gate824inter5, gate824inter6, gate824inter7, gate824inter8, gate824inter9, gate824inter10, gate824inter11, gate824inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate363inter0, gate363inter1, gate363inter2, gate363inter3, gate363inter4, gate363inter5, gate363inter6, gate363inter7, gate363inter8, gate363inter9, gate363inter10, gate363inter11, gate363inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate780inter0, gate780inter1, gate780inter2, gate780inter3, gate780inter4, gate780inter5, gate780inter6, gate780inter7, gate780inter8, gate780inter9, gate780inter10, gate780inter11, gate780inter12, gate752inter0, gate752inter1, gate752inter2, gate752inter3, gate752inter4, gate752inter5, gate752inter6, gate752inter7, gate752inter8, gate752inter9, gate752inter10, gate752inter11, gate752inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate624inter0, gate624inter1, gate624inter2, gate624inter3, gate624inter4, gate624inter5, gate624inter6, gate624inter7, gate624inter8, gate624inter9, gate624inter10, gate624inter11, gate624inter12, gate834inter0, gate834inter1, gate834inter2, gate834inter3, gate834inter4, gate834inter5, gate834inter6, gate834inter7, gate834inter8, gate834inter9, gate834inter10, gate834inter11, gate834inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate626inter0, gate626inter1, gate626inter2, gate626inter3, gate626inter4, gate626inter5, gate626inter6, gate626inter7, gate626inter8, gate626inter9, gate626inter10, gate626inter11, gate626inter12, gate366inter0, gate366inter1, gate366inter2, gate366inter3, gate366inter4, gate366inter5, gate366inter6, gate366inter7, gate366inter8, gate366inter9, gate366inter10, gate366inter11, gate366inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate804inter0, gate804inter1, gate804inter2, gate804inter3, gate804inter4, gate804inter5, gate804inter6, gate804inter7, gate804inter8, gate804inter9, gate804inter10, gate804inter11, gate804inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate797inter0, gate797inter1, gate797inter2, gate797inter3, gate797inter4, gate797inter5, gate797inter6, gate797inter7, gate797inter8, gate797inter9, gate797inter10, gate797inter11, gate797inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate805inter0, gate805inter1, gate805inter2, gate805inter3, gate805inter4, gate805inter5, gate805inter6, gate805inter7, gate805inter8, gate805inter9, gate805inter10, gate805inter11, gate805inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate812inter0, gate812inter1, gate812inter2, gate812inter3, gate812inter4, gate812inter5, gate812inter6, gate812inter7, gate812inter8, gate812inter9, gate812inter10, gate812inter11, gate812inter12, gate608inter0, gate608inter1, gate608inter2, gate608inter3, gate608inter4, gate608inter5, gate608inter6, gate608inter7, gate608inter8, gate608inter9, gate608inter10, gate608inter11, gate608inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate545inter0, gate545inter1, gate545inter2, gate545inter3, gate545inter4, gate545inter5, gate545inter6, gate545inter7, gate545inter8, gate545inter9, gate545inter10, gate545inter11, gate545inter12, gate876inter0, gate876inter1, gate876inter2, gate876inter3, gate876inter4, gate876inter5, gate876inter6, gate876inter7, gate876inter8, gate876inter9, gate876inter10, gate876inter11, gate876inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate878inter0, gate878inter1, gate878inter2, gate878inter3, gate878inter4, gate878inter5, gate878inter6, gate878inter7, gate878inter8, gate878inter9, gate878inter10, gate878inter11, gate878inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate556inter0, gate556inter1, gate556inter2, gate556inter3, gate556inter4, gate556inter5, gate556inter6, gate556inter7, gate556inter8, gate556inter9, gate556inter10, gate556inter11, gate556inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate345inter0, gate345inter1, gate345inter2, gate345inter3, gate345inter4, gate345inter5, gate345inter6, gate345inter7, gate345inter8, gate345inter9, gate345inter10, gate345inter11, gate345inter12, gate632inter0, gate632inter1, gate632inter2, gate632inter3, gate632inter4, gate632inter5, gate632inter6, gate632inter7, gate632inter8, gate632inter9, gate632inter10, gate632inter11, gate632inter12, gate616inter0, gate616inter1, gate616inter2, gate616inter3, gate616inter4, gate616inter5, gate616inter6, gate616inter7, gate616inter8, gate616inter9, gate616inter10, gate616inter11, gate616inter12, gate686inter0, gate686inter1, gate686inter2, gate686inter3, gate686inter4, gate686inter5, gate686inter6, gate686inter7, gate686inter8, gate686inter9, gate686inter10, gate686inter11, gate686inter12, gate818inter0, gate818inter1, gate818inter2, gate818inter3, gate818inter4, gate818inter5, gate818inter6, gate818inter7, gate818inter8, gate818inter9, gate818inter10, gate818inter11, gate818inter12, gate835inter0, gate835inter1, gate835inter2, gate835inter3, gate835inter4, gate835inter5, gate835inter6, gate835inter7, gate835inter8, gate835inter9, gate835inter10, gate835inter11, gate835inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate561inter0, gate561inter1, gate561inter2, gate561inter3, gate561inter4, gate561inter5, gate561inter6, gate561inter7, gate561inter8, gate561inter9, gate561inter10, gate561inter11, gate561inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate380inter0, gate380inter1, gate380inter2, gate380inter3, gate380inter4, gate380inter5, gate380inter6, gate380inter7, gate380inter8, gate380inter9, gate380inter10, gate380inter11, gate380inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate613inter0, gate613inter1, gate613inter2, gate613inter3, gate613inter4, gate613inter5, gate613inter6, gate613inter7, gate613inter8, gate613inter9, gate613inter10, gate613inter11, gate613inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate771inter0, gate771inter1, gate771inter2, gate771inter3, gate771inter4, gate771inter5, gate771inter6, gate771inter7, gate771inter8, gate771inter9, gate771inter10, gate771inter11, gate771inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate682inter0, gate682inter1, gate682inter2, gate682inter3, gate682inter4, gate682inter5, gate682inter6, gate682inter7, gate682inter8, gate682inter9, gate682inter10, gate682inter11, gate682inter12, gate572inter0, gate572inter1, gate572inter2, gate572inter3, gate572inter4, gate572inter5, gate572inter6, gate572inter7, gate572inter8, gate572inter9, gate572inter10, gate572inter11, gate572inter12, gate843inter0, gate843inter1, gate843inter2, gate843inter3, gate843inter4, gate843inter5, gate843inter6, gate843inter7, gate843inter8, gate843inter9, gate843inter10, gate843inter11, gate843inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate837inter0, gate837inter1, gate837inter2, gate837inter3, gate837inter4, gate837inter5, gate837inter6, gate837inter7, gate837inter8, gate837inter9, gate837inter10, gate837inter11, gate837inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate640inter0, gate640inter1, gate640inter2, gate640inter3, gate640inter4, gate640inter5, gate640inter6, gate640inter7, gate640inter8, gate640inter9, gate640inter10, gate640inter11, gate640inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate766inter0, gate766inter1, gate766inter2, gate766inter3, gate766inter4, gate766inter5, gate766inter6, gate766inter7, gate766inter8, gate766inter9, gate766inter10, gate766inter11, gate766inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate306inter0, gate306inter1, gate306inter2, gate306inter3, gate306inter4, gate306inter5, gate306inter6, gate306inter7, gate306inter8, gate306inter9, gate306inter10, gate306inter11, gate306inter12, gate303inter0, gate303inter1, gate303inter2, gate303inter3, gate303inter4, gate303inter5, gate303inter6, gate303inter7, gate303inter8, gate303inter9, gate303inter10, gate303inter11, gate303inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate838inter0, gate838inter1, gate838inter2, gate838inter3, gate838inter4, gate838inter5, gate838inter6, gate838inter7, gate838inter8, gate838inter9, gate838inter10, gate838inter11, gate838inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate541inter0, gate541inter1, gate541inter2, gate541inter3, gate541inter4, gate541inter5, gate541inter6, gate541inter7, gate541inter8, gate541inter9, gate541inter10, gate541inter11, gate541inter12, gate374inter0, gate374inter1, gate374inter2, gate374inter3, gate374inter4, gate374inter5, gate374inter6, gate374inter7, gate374inter8, gate374inter9, gate374inter10, gate374inter11, gate374inter12, gate802inter0, gate802inter1, gate802inter2, gate802inter3, gate802inter4, gate802inter5, gate802inter6, gate802inter7, gate802inter8, gate802inter9, gate802inter10, gate802inter11, gate802inter12, gate663inter0, gate663inter1, gate663inter2, gate663inter3, gate663inter4, gate663inter5, gate663inter6, gate663inter7, gate663inter8, gate663inter9, gate663inter10, gate663inter11, gate663inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate315inter0, gate315inter1, gate315inter2, gate315inter3, gate315inter4, gate315inter5, gate315inter6, gate315inter7, gate315inter8, gate315inter9, gate315inter10, gate315inter11, gate315inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate350inter0, gate350inter1, gate350inter2, gate350inter3, gate350inter4, gate350inter5, gate350inter6, gate350inter7, gate350inter8, gate350inter9, gate350inter10, gate350inter11, gate350inter12, gate321inter0, gate321inter1, gate321inter2, gate321inter3, gate321inter4, gate321inter5, gate321inter6, gate321inter7, gate321inter8, gate321inter9, gate321inter10, gate321inter11, gate321inter12, gate536inter0, gate536inter1, gate536inter2, gate536inter3, gate536inter4, gate536inter5, gate536inter6, gate536inter7, gate536inter8, gate536inter9, gate536inter10, gate536inter11, gate536inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate623inter0, gate623inter1, gate623inter2, gate623inter3, gate623inter4, gate623inter5, gate623inter6, gate623inter7, gate623inter8, gate623inter9, gate623inter10, gate623inter11, gate623inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );

  xor2  gate1581(.a(N91), .b(N66), .O(gate18inter0));
  nand2 gate1582(.a(gate18inter0), .b(s_100), .O(gate18inter1));
  and2  gate1583(.a(N91), .b(N66), .O(gate18inter2));
  inv1  gate1584(.a(s_100), .O(gate18inter3));
  inv1  gate1585(.a(s_101), .O(gate18inter4));
  nand2 gate1586(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1587(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1588(.a(N66), .O(gate18inter7));
  inv1  gate1589(.a(N91), .O(gate18inter8));
  nand2 gate1590(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1591(.a(s_101), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1592(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1593(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1594(.a(gate18inter12), .b(gate18inter1), .O(N252));
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );

  xor2  gate1651(.a(N331), .b(N306), .O(gate80inter0));
  nand2 gate1652(.a(gate80inter0), .b(s_110), .O(gate80inter1));
  and2  gate1653(.a(N331), .b(N306), .O(gate80inter2));
  inv1  gate1654(.a(s_110), .O(gate80inter3));
  inv1  gate1655(.a(s_111), .O(gate80inter4));
  nand2 gate1656(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1657(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1658(.a(N306), .O(gate80inter7));
  inv1  gate1659(.a(N331), .O(gate80inter8));
  nand2 gate1660(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1661(.a(s_111), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1662(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1663(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1664(.a(gate80inter12), .b(gate80inter1), .O(N555));
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );

  xor2  gate1679(.a(N300), .b(N256), .O(gate100inter0));
  nand2 gate1680(.a(gate100inter0), .b(s_114), .O(gate100inter1));
  and2  gate1681(.a(N300), .b(N256), .O(gate100inter2));
  inv1  gate1682(.a(s_114), .O(gate100inter3));
  inv1  gate1683(.a(s_115), .O(gate100inter4));
  nand2 gate1684(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1685(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1686(.a(N256), .O(gate100inter7));
  inv1  gate1687(.a(N300), .O(gate100inter8));
  nand2 gate1688(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1689(.a(s_115), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1690(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1691(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1692(.a(gate100inter12), .b(gate100inter1), .O(N612));
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );

  xor2  gate1707(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate1708(.a(gate245inter0), .b(s_118), .O(gate245inter1));
  and2  gate1709(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate1710(.a(s_118), .O(gate245inter3));
  inv1  gate1711(.a(s_119), .O(gate245inter4));
  nand2 gate1712(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1713(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1714(.a(N745), .O(gate245inter7));
  inv1  gate1715(.a(N1005), .O(gate245inter8));
  nand2 gate1716(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1717(.a(s_119), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1718(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1719(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1720(.a(gate245inter12), .b(gate245inter1), .O(N1130));
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );

  xor2  gate2169(.a(N938), .b(N1010), .O(gate271inter0));
  nand2 gate2170(.a(gate271inter0), .b(s_184), .O(gate271inter1));
  and2  gate2171(.a(N938), .b(N1010), .O(gate271inter2));
  inv1  gate2172(.a(s_184), .O(gate271inter3));
  inv1  gate2173(.a(s_185), .O(gate271inter4));
  nand2 gate2174(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2175(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2176(.a(N1010), .O(gate271inter7));
  inv1  gate2177(.a(N938), .O(gate271inter8));
  nand2 gate2178(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2179(.a(s_185), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2180(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2181(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2182(.a(gate271inter12), .b(gate271inter1), .O(N1206));
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate1329(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate1330(.a(gate277inter0), .b(s_64), .O(gate277inter1));
  and2  gate1331(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate1332(.a(s_64), .O(gate277inter3));
  inv1  gate1333(.a(s_65), .O(gate277inter4));
  nand2 gate1334(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1335(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1336(.a(N1019), .O(gate277inter7));
  inv1  gate1337(.a(N950), .O(gate277inter8));
  nand2 gate1338(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1339(.a(s_65), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1340(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1341(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1342(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );

  xor2  gate1189(.a(N980), .b(N1043), .O(gate294inter0));
  nand2 gate1190(.a(gate294inter0), .b(s_44), .O(gate294inter1));
  and2  gate1191(.a(N980), .b(N1043), .O(gate294inter2));
  inv1  gate1192(.a(s_44), .O(gate294inter3));
  inv1  gate1193(.a(s_45), .O(gate294inter4));
  nand2 gate1194(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1195(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1196(.a(N1043), .O(gate294inter7));
  inv1  gate1197(.a(N980), .O(gate294inter8));
  nand2 gate1198(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1199(.a(s_45), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1200(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1201(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1202(.a(gate294inter12), .b(gate294inter1), .O(N1229));
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );

  xor2  gate1231(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate1232(.a(gate297inter0), .b(s_50), .O(gate297inter1));
  and2  gate1233(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate1234(.a(s_50), .O(gate297inter3));
  inv1  gate1235(.a(s_51), .O(gate297inter4));
  nand2 gate1236(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate1237(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate1238(.a(N1119), .O(gate297inter7));
  inv1  gate1239(.a(N1120), .O(gate297inter8));
  nand2 gate1240(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate1241(.a(s_51), .b(gate297inter3), .O(gate297inter10));
  nor2  gate1242(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate1243(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate1244(.a(gate297inter12), .b(gate297inter1), .O(N1232));

  xor2  gate2267(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate2268(.a(gate298inter0), .b(s_198), .O(gate298inter1));
  and2  gate2269(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate2270(.a(s_198), .O(gate298inter3));
  inv1  gate2271(.a(s_199), .O(gate298inter4));
  nand2 gate2272(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate2273(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate2274(.a(N1121), .O(gate298inter7));
  inv1  gate2275(.a(N1122), .O(gate298inter8));
  nand2 gate2276(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate2277(.a(s_199), .b(gate298inter3), .O(gate298inter10));
  nor2  gate2278(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate2279(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate2280(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );

  xor2  gate2015(.a(N1001), .b(N1049), .O(gate303inter0));
  nand2 gate2016(.a(gate303inter0), .b(s_162), .O(gate303inter1));
  and2  gate2017(.a(N1001), .b(N1049), .O(gate303inter2));
  inv1  gate2018(.a(s_162), .O(gate303inter3));
  inv1  gate2019(.a(s_163), .O(gate303inter4));
  nand2 gate2020(.a(gate303inter4), .b(gate303inter3), .O(gate303inter5));
  nor2  gate2021(.a(gate303inter5), .b(gate303inter2), .O(gate303inter6));
  inv1  gate2022(.a(N1049), .O(gate303inter7));
  inv1  gate2023(.a(N1001), .O(gate303inter8));
  nand2 gate2024(.a(gate303inter8), .b(gate303inter7), .O(gate303inter9));
  nand2 gate2025(.a(s_163), .b(gate303inter3), .O(gate303inter10));
  nor2  gate2026(.a(gate303inter10), .b(gate303inter9), .O(gate303inter11));
  nor2  gate2027(.a(gate303inter11), .b(gate303inter6), .O(gate303inter12));
  nand2 gate2028(.a(gate303inter12), .b(gate303inter1), .O(N1242));
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );

  xor2  gate2001(.a(N1133), .b(N1132), .O(gate306inter0));
  nand2 gate2002(.a(gate306inter0), .b(s_160), .O(gate306inter1));
  and2  gate2003(.a(N1133), .b(N1132), .O(gate306inter2));
  inv1  gate2004(.a(s_160), .O(gate306inter3));
  inv1  gate2005(.a(s_161), .O(gate306inter4));
  nand2 gate2006(.a(gate306inter4), .b(gate306inter3), .O(gate306inter5));
  nor2  gate2007(.a(gate306inter5), .b(gate306inter2), .O(gate306inter6));
  inv1  gate2008(.a(N1132), .O(gate306inter7));
  inv1  gate2009(.a(N1133), .O(gate306inter8));
  nand2 gate2010(.a(gate306inter8), .b(gate306inter7), .O(gate306inter9));
  nand2 gate2011(.a(s_161), .b(gate306inter3), .O(gate306inter10));
  nor2  gate2012(.a(gate306inter10), .b(gate306inter9), .O(gate306inter11));
  nor2  gate2013(.a(gate306inter11), .b(gate306inter6), .O(gate306inter12));
  nand2 gate2014(.a(gate306inter12), .b(gate306inter1), .O(N1249));
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );

  xor2  gate1735(.a(N1205), .b(N688), .O(gate313inter0));
  nand2 gate1736(.a(gate313inter0), .b(s_122), .O(gate313inter1));
  and2  gate1737(.a(N1205), .b(N688), .O(gate313inter2));
  inv1  gate1738(.a(s_122), .O(gate313inter3));
  inv1  gate1739(.a(s_123), .O(gate313inter4));
  nand2 gate1740(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate1741(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate1742(.a(N688), .O(gate313inter7));
  inv1  gate1743(.a(N1205), .O(gate313inter8));
  nand2 gate1744(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate1745(.a(s_123), .b(gate313inter3), .O(gate313inter10));
  nor2  gate1746(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate1747(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate1748(.a(gate313inter12), .b(gate313inter1), .O(N1309));
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );

  xor2  gate2141(.a(N1209), .b(N694), .O(gate315inter0));
  nand2 gate2142(.a(gate315inter0), .b(s_180), .O(gate315inter1));
  and2  gate2143(.a(N1209), .b(N694), .O(gate315inter2));
  inv1  gate2144(.a(s_180), .O(gate315inter3));
  inv1  gate2145(.a(s_181), .O(gate315inter4));
  nand2 gate2146(.a(gate315inter4), .b(gate315inter3), .O(gate315inter5));
  nor2  gate2147(.a(gate315inter5), .b(gate315inter2), .O(gate315inter6));
  inv1  gate2148(.a(N694), .O(gate315inter7));
  inv1  gate2149(.a(N1209), .O(gate315inter8));
  nand2 gate2150(.a(gate315inter8), .b(gate315inter7), .O(gate315inter9));
  nand2 gate2151(.a(s_181), .b(gate315inter3), .O(gate315inter10));
  nor2  gate2152(.a(gate315inter10), .b(gate315inter9), .O(gate315inter11));
  nor2  gate2153(.a(gate315inter11), .b(gate315inter6), .O(gate315inter12));
  nand2 gate2154(.a(gate315inter12), .b(gate315inter1), .O(N1311));

  xor2  gate1819(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate1820(.a(gate316inter0), .b(s_134), .O(gate316inter1));
  and2  gate1821(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate1822(.a(s_134), .O(gate316inter3));
  inv1  gate1823(.a(s_135), .O(gate316inter4));
  nand2 gate1824(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate1825(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate1826(.a(N697), .O(gate316inter7));
  inv1  gate1827(.a(N1211), .O(gate316inter8));
  nand2 gate1828(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate1829(.a(s_135), .b(gate316inter3), .O(gate316inter10));
  nor2  gate1830(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate1831(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate1832(.a(gate316inter12), .b(gate316inter1), .O(N1312));

  xor2  gate1371(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate1372(.a(gate317inter0), .b(s_70), .O(gate317inter1));
  and2  gate1373(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate1374(.a(s_70), .O(gate317inter3));
  inv1  gate1375(.a(s_71), .O(gate317inter4));
  nand2 gate1376(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate1377(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate1378(.a(N700), .O(gate317inter7));
  inv1  gate1379(.a(N1213), .O(gate317inter8));
  nand2 gate1380(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate1381(.a(s_71), .b(gate317inter3), .O(gate317inter10));
  nor2  gate1382(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate1383(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate1384(.a(gate317inter12), .b(gate317inter1), .O(N1313));
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );

  xor2  gate2197(.a(N1225), .b(N712), .O(gate321inter0));
  nand2 gate2198(.a(gate321inter0), .b(s_188), .O(gate321inter1));
  and2  gate2199(.a(N1225), .b(N712), .O(gate321inter2));
  inv1  gate2200(.a(s_188), .O(gate321inter3));
  inv1  gate2201(.a(s_189), .O(gate321inter4));
  nand2 gate2202(.a(gate321inter4), .b(gate321inter3), .O(gate321inter5));
  nor2  gate2203(.a(gate321inter5), .b(gate321inter2), .O(gate321inter6));
  inv1  gate2204(.a(N712), .O(gate321inter7));
  inv1  gate2205(.a(N1225), .O(gate321inter8));
  nand2 gate2206(.a(gate321inter8), .b(gate321inter7), .O(gate321inter9));
  nand2 gate2207(.a(s_189), .b(gate321inter3), .O(gate321inter10));
  nor2  gate2208(.a(gate321inter10), .b(gate321inter9), .O(gate321inter11));
  nor2  gate2209(.a(gate321inter11), .b(gate321inter6), .O(gate321inter12));
  nand2 gate2210(.a(gate321inter12), .b(gate321inter1), .O(N1317));

  xor2  gate1623(.a(N1228), .b(N715), .O(gate322inter0));
  nand2 gate1624(.a(gate322inter0), .b(s_106), .O(gate322inter1));
  and2  gate1625(.a(N1228), .b(N715), .O(gate322inter2));
  inv1  gate1626(.a(s_106), .O(gate322inter3));
  inv1  gate1627(.a(s_107), .O(gate322inter4));
  nand2 gate1628(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate1629(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate1630(.a(N715), .O(gate322inter7));
  inv1  gate1631(.a(N1228), .O(gate322inter8));
  nand2 gate1632(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate1633(.a(s_107), .b(gate322inter3), .O(gate322inter10));
  nor2  gate1634(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate1635(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate1636(.a(gate322inter12), .b(gate322inter1), .O(N1318));
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );

  xor2  gate1973(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate1974(.a(gate326inter0), .b(s_156), .O(gate326inter1));
  and2  gate1975(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate1976(.a(s_156), .O(gate326inter3));
  inv1  gate1977(.a(s_157), .O(gate326inter4));
  nand2 gate1978(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate1979(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate1980(.a(N733), .O(gate326inter7));
  inv1  gate1981(.a(N1241), .O(gate326inter8));
  nand2 gate1982(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate1983(.a(s_157), .b(gate326inter3), .O(gate326inter10));
  nor2  gate1984(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate1985(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate1986(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );

  xor2  gate2225(.a(N1210), .b(N1311), .O(gate337inter0));
  nand2 gate2226(.a(gate337inter0), .b(s_192), .O(gate337inter1));
  and2  gate2227(.a(N1210), .b(N1311), .O(gate337inter2));
  inv1  gate2228(.a(s_192), .O(gate337inter3));
  inv1  gate2229(.a(s_193), .O(gate337inter4));
  nand2 gate2230(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate2231(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate2232(.a(N1311), .O(gate337inter7));
  inv1  gate2233(.a(N1210), .O(gate337inter8));
  nand2 gate2234(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate2235(.a(s_193), .b(gate337inter3), .O(gate337inter10));
  nor2  gate2236(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate2237(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate2238(.a(gate337inter12), .b(gate337inter1), .O(N1358));
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );

  xor2  gate951(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate952(.a(gate342inter0), .b(s_10), .O(gate342inter1));
  and2  gate953(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate954(.a(s_10), .O(gate342inter3));
  inv1  gate955(.a(s_11), .O(gate342inter4));
  nand2 gate956(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate957(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate958(.a(N1316), .O(gate342inter7));
  inv1  gate959(.a(N1224), .O(gate342inter8));
  nand2 gate960(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate961(.a(s_11), .b(gate342inter3), .O(gate342inter10));
  nor2  gate962(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate963(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate964(.a(gate342inter12), .b(gate342inter1), .O(N1373));
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );

  xor2  gate1497(.a(N1231), .b(N1322), .O(gate345inter0));
  nand2 gate1498(.a(gate345inter0), .b(s_88), .O(gate345inter1));
  and2  gate1499(.a(N1231), .b(N1322), .O(gate345inter2));
  inv1  gate1500(.a(s_88), .O(gate345inter3));
  inv1  gate1501(.a(s_89), .O(gate345inter4));
  nand2 gate1502(.a(gate345inter4), .b(gate345inter3), .O(gate345inter5));
  nor2  gate1503(.a(gate345inter5), .b(gate345inter2), .O(gate345inter6));
  inv1  gate1504(.a(N1322), .O(gate345inter7));
  inv1  gate1505(.a(N1231), .O(gate345inter8));
  nand2 gate1506(.a(gate345inter8), .b(gate345inter7), .O(gate345inter9));
  nand2 gate1507(.a(s_89), .b(gate345inter3), .O(gate345inter10));
  nor2  gate1508(.a(gate345inter10), .b(gate345inter9), .O(gate345inter11));
  nor2  gate1509(.a(gate345inter11), .b(gate345inter6), .O(gate345inter12));
  nand2 gate1510(.a(gate345inter12), .b(gate345inter1), .O(N1383));
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate1049(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate1050(.a(gate347inter0), .b(s_24), .O(gate347inter1));
  and2  gate1051(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate1052(.a(s_24), .O(gate347inter3));
  inv1  gate1053(.a(s_25), .O(gate347inter4));
  nand2 gate1054(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate1055(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate1056(.a(N1232), .O(gate347inter7));
  inv1  gate1057(.a(N990), .O(gate347inter8));
  nand2 gate1058(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate1059(.a(s_25), .b(gate347inter3), .O(gate347inter10));
  nor2  gate1060(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate1061(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate1062(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );

  xor2  gate2183(.a(N1239), .b(N1327), .O(gate350inter0));
  nand2 gate2184(.a(gate350inter0), .b(s_186), .O(gate350inter1));
  and2  gate2185(.a(N1239), .b(N1327), .O(gate350inter2));
  inv1  gate2186(.a(s_186), .O(gate350inter3));
  inv1  gate2187(.a(s_187), .O(gate350inter4));
  nand2 gate2188(.a(gate350inter4), .b(gate350inter3), .O(gate350inter5));
  nor2  gate2189(.a(gate350inter5), .b(gate350inter2), .O(gate350inter6));
  inv1  gate2190(.a(N1327), .O(gate350inter7));
  inv1  gate2191(.a(N1239), .O(gate350inter8));
  nand2 gate2192(.a(gate350inter8), .b(gate350inter7), .O(gate350inter9));
  nand2 gate2193(.a(s_187), .b(gate350inter3), .O(gate350inter10));
  nor2  gate2194(.a(gate350inter10), .b(gate350inter9), .O(gate350inter11));
  nor2  gate2195(.a(gate350inter11), .b(gate350inter6), .O(gate350inter12));
  nand2 gate2196(.a(gate350inter12), .b(gate350inter1), .O(N1390));
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );

  xor2  gate1805(.a(N1388), .b(N637), .O(gate362inter0));
  nand2 gate1806(.a(gate362inter0), .b(s_132), .O(gate362inter1));
  and2  gate1807(.a(N1388), .b(N637), .O(gate362inter2));
  inv1  gate1808(.a(s_132), .O(gate362inter3));
  inv1  gate1809(.a(s_133), .O(gate362inter4));
  nand2 gate1810(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate1811(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate1812(.a(N637), .O(gate362inter7));
  inv1  gate1813(.a(N1388), .O(gate362inter8));
  nand2 gate1814(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate1815(.a(s_133), .b(gate362inter3), .O(gate362inter10));
  nor2  gate1816(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate1817(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate1818(.a(gate362inter12), .b(gate362inter1), .O(N1434));

  xor2  gate1035(.a(N1396), .b(N640), .O(gate363inter0));
  nand2 gate1036(.a(gate363inter0), .b(s_22), .O(gate363inter1));
  and2  gate1037(.a(N1396), .b(N640), .O(gate363inter2));
  inv1  gate1038(.a(s_22), .O(gate363inter3));
  inv1  gate1039(.a(s_23), .O(gate363inter4));
  nand2 gate1040(.a(gate363inter4), .b(gate363inter3), .O(gate363inter5));
  nor2  gate1041(.a(gate363inter5), .b(gate363inter2), .O(gate363inter6));
  inv1  gate1042(.a(N640), .O(gate363inter7));
  inv1  gate1043(.a(N1396), .O(gate363inter8));
  nand2 gate1044(.a(gate363inter8), .b(gate363inter7), .O(gate363inter9));
  nand2 gate1045(.a(s_23), .b(gate363inter3), .O(gate363inter10));
  nor2  gate1046(.a(gate363inter10), .b(gate363inter9), .O(gate363inter11));
  nor2  gate1047(.a(gate363inter11), .b(gate363inter6), .O(gate363inter12));
  nand2 gate1048(.a(gate363inter12), .b(gate363inter1), .O(N1438));
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );

  xor2  gate1161(.a(N1148), .b(N1355), .O(gate366inter0));
  nand2 gate1162(.a(gate366inter0), .b(s_40), .O(gate366inter1));
  and2  gate1163(.a(N1148), .b(N1355), .O(gate366inter2));
  inv1  gate1164(.a(s_40), .O(gate366inter3));
  inv1  gate1165(.a(s_41), .O(gate366inter4));
  nand2 gate1166(.a(gate366inter4), .b(gate366inter3), .O(gate366inter5));
  nor2  gate1167(.a(gate366inter5), .b(gate366inter2), .O(gate366inter6));
  inv1  gate1168(.a(N1355), .O(gate366inter7));
  inv1  gate1169(.a(N1148), .O(gate366inter8));
  nand2 gate1170(.a(gate366inter8), .b(gate366inter7), .O(gate366inter9));
  nand2 gate1171(.a(s_41), .b(gate366inter3), .O(gate366inter10));
  nor2  gate1172(.a(gate366inter10), .b(gate366inter9), .O(gate366inter11));
  nor2  gate1173(.a(gate366inter11), .b(gate366inter6), .O(gate366inter12));
  nand2 gate1174(.a(gate366inter12), .b(gate366inter1), .O(N1443));
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );

  xor2  gate2085(.a(N1153), .b(N1367), .O(gate374inter0));
  nand2 gate2086(.a(gate374inter0), .b(s_172), .O(gate374inter1));
  and2  gate2087(.a(N1153), .b(N1367), .O(gate374inter2));
  inv1  gate2088(.a(s_172), .O(gate374inter3));
  inv1  gate2089(.a(s_173), .O(gate374inter4));
  nand2 gate2090(.a(gate374inter4), .b(gate374inter3), .O(gate374inter5));
  nor2  gate2091(.a(gate374inter5), .b(gate374inter2), .O(gate374inter6));
  inv1  gate2092(.a(N1367), .O(gate374inter7));
  inv1  gate2093(.a(N1153), .O(gate374inter8));
  nand2 gate2094(.a(gate374inter8), .b(gate374inter7), .O(gate374inter9));
  nand2 gate2095(.a(s_173), .b(gate374inter3), .O(gate374inter10));
  nor2  gate2096(.a(gate374inter10), .b(gate374inter9), .O(gate374inter11));
  nor2  gate2097(.a(gate374inter11), .b(gate374inter6), .O(gate374inter12));
  nand2 gate2098(.a(gate374inter12), .b(gate374inter1), .O(N1453));
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );

  xor2  gate1637(.a(N1157), .b(N1379), .O(gate380inter0));
  nand2 gate1638(.a(gate380inter0), .b(s_108), .O(gate380inter1));
  and2  gate1639(.a(N1157), .b(N1379), .O(gate380inter2));
  inv1  gate1640(.a(s_108), .O(gate380inter3));
  inv1  gate1641(.a(s_109), .O(gate380inter4));
  nand2 gate1642(.a(gate380inter4), .b(gate380inter3), .O(gate380inter5));
  nor2  gate1643(.a(gate380inter5), .b(gate380inter2), .O(gate380inter6));
  inv1  gate1644(.a(N1379), .O(gate380inter7));
  inv1  gate1645(.a(N1157), .O(gate380inter8));
  nand2 gate1646(.a(gate380inter8), .b(gate380inter7), .O(gate380inter9));
  nand2 gate1647(.a(s_109), .b(gate380inter3), .O(gate380inter10));
  nor2  gate1648(.a(gate380inter10), .b(gate380inter9), .O(gate380inter11));
  nor2  gate1649(.a(gate380inter11), .b(gate380inter6), .O(gate380inter12));
  nand2 gate1650(.a(gate380inter12), .b(gate380inter1), .O(N1459));
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );

  xor2  gate881(.a(N1412), .b(N1345), .O(gate385inter0));
  nand2 gate882(.a(gate385inter0), .b(s_0), .O(gate385inter1));
  and2  gate883(.a(N1412), .b(N1345), .O(gate385inter2));
  inv1  gate884(.a(s_0), .O(gate385inter3));
  inv1  gate885(.a(s_1), .O(gate385inter4));
  nand2 gate886(.a(gate385inter4), .b(gate385inter3), .O(gate385inter5));
  nor2  gate887(.a(gate385inter5), .b(gate385inter2), .O(gate385inter6));
  inv1  gate888(.a(N1345), .O(gate385inter7));
  inv1  gate889(.a(N1412), .O(gate385inter8));
  nand2 gate890(.a(gate385inter8), .b(gate385inter7), .O(gate385inter9));
  nand2 gate891(.a(s_1), .b(gate385inter3), .O(gate385inter10));
  nor2  gate892(.a(gate385inter10), .b(gate385inter9), .O(gate385inter11));
  nor2  gate893(.a(gate385inter11), .b(gate385inter6), .O(gate385inter12));
  nand2 gate894(.a(gate385inter12), .b(gate385inter1), .O(N1464));
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );

  xor2  gate1413(.a(N1433), .b(N1387), .O(gate390inter0));
  nand2 gate1414(.a(gate390inter0), .b(s_76), .O(gate390inter1));
  and2  gate1415(.a(N1433), .b(N1387), .O(gate390inter2));
  inv1  gate1416(.a(s_76), .O(gate390inter3));
  inv1  gate1417(.a(s_77), .O(gate390inter4));
  nand2 gate1418(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1419(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1420(.a(N1387), .O(gate390inter7));
  inv1  gate1421(.a(N1433), .O(gate390inter8));
  nand2 gate1422(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1423(.a(s_77), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1424(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1425(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1426(.a(gate390inter12), .b(gate390inter1), .O(N1472));
inv1 gate391( .a(N1390), .O(N1475) );

  xor2  gate1245(.a(N1240), .b(N1390), .O(gate392inter0));
  nand2 gate1246(.a(gate392inter0), .b(s_52), .O(gate392inter1));
  and2  gate1247(.a(N1240), .b(N1390), .O(gate392inter2));
  inv1  gate1248(.a(s_52), .O(gate392inter3));
  inv1  gate1249(.a(s_53), .O(gate392inter4));
  nand2 gate1250(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1251(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1252(.a(N1390), .O(gate392inter7));
  inv1  gate1253(.a(N1240), .O(gate392inter8));
  nand2 gate1254(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1255(.a(s_53), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1256(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1257(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1258(.a(gate392inter12), .b(gate392inter1), .O(N1476));
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );

  xor2  gate1889(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate1890(.a(gate402inter0), .b(s_144), .O(gate402inter1));
  and2  gate1891(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate1892(.a(s_144), .O(gate402inter3));
  inv1  gate1893(.a(s_145), .O(gate402inter4));
  nand2 gate1894(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1895(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1896(.a(N955), .O(gate402inter7));
  inv1  gate1897(.a(N1454), .O(gate402inter8));
  nand2 gate1898(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1899(.a(s_145), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1900(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1901(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1902(.a(gate402inter12), .b(gate402inter1), .O(N1493));

  xor2  gate1693(.a(N1456), .b(N951), .O(gate403inter0));
  nand2 gate1694(.a(gate403inter0), .b(s_116), .O(gate403inter1));
  and2  gate1695(.a(N1456), .b(N951), .O(gate403inter2));
  inv1  gate1696(.a(s_116), .O(gate403inter3));
  inv1  gate1697(.a(s_117), .O(gate403inter4));
  nand2 gate1698(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1699(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1700(.a(N951), .O(gate403inter7));
  inv1  gate1701(.a(N1456), .O(gate403inter8));
  nand2 gate1702(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1703(.a(s_117), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1704(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1705(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1706(.a(gate403inter12), .b(gate403inter1), .O(N1494));
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );

  xor2  gate1861(.a(N1468), .b(N965), .O(gate408inter0));
  nand2 gate1862(.a(gate408inter0), .b(s_140), .O(gate408inter1));
  and2  gate1863(.a(N1468), .b(N965), .O(gate408inter2));
  inv1  gate1864(.a(s_140), .O(gate408inter3));
  inv1  gate1865(.a(s_141), .O(gate408inter4));
  nand2 gate1866(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1867(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1868(.a(N965), .O(gate408inter7));
  inv1  gate1869(.a(N1468), .O(gate408inter8));
  nand2 gate1870(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1871(.a(s_141), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1872(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1873(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1874(.a(gate408inter12), .b(gate408inter1), .O(N1500));
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );

  xor2  gate1945(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate1946(.a(gate410inter0), .b(s_152), .O(gate410inter1));
  and2  gate1947(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate1948(.a(s_152), .O(gate410inter3));
  inv1  gate1949(.a(s_153), .O(gate410inter4));
  nand2 gate1950(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1951(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1952(.a(N994), .O(gate410inter7));
  inv1  gate1953(.a(N1475), .O(gate410inter8));
  nand2 gate1954(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1955(.a(s_153), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1956(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1957(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1958(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );

  xor2  gate1441(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate1442(.a(gate413inter0), .b(s_80), .O(gate413inter1));
  and2  gate1443(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate1444(.a(s_80), .O(gate413inter3));
  inv1  gate1445(.a(s_81), .O(gate413inter4));
  nand2 gate1446(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1447(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1448(.a(N1445), .O(gate413inter7));
  inv1  gate1449(.a(N1488), .O(gate413inter8));
  nand2 gate1450(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1451(.a(s_81), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1452(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1453(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1454(.a(gate413inter12), .b(gate413inter1), .O(N1514));

  xor2  gate1175(.a(N1489), .b(N1447), .O(gate414inter0));
  nand2 gate1176(.a(gate414inter0), .b(s_42), .O(gate414inter1));
  and2  gate1177(.a(N1489), .b(N1447), .O(gate414inter2));
  inv1  gate1178(.a(s_42), .O(gate414inter3));
  inv1  gate1179(.a(s_43), .O(gate414inter4));
  nand2 gate1180(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1181(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1182(.a(N1447), .O(gate414inter7));
  inv1  gate1183(.a(N1489), .O(gate414inter8));
  nand2 gate1184(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1185(.a(s_43), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1186(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1187(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1188(.a(gate414inter12), .b(gate414inter1), .O(N1517));
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );

  xor2  gate1959(.a(N1496), .b(N1459), .O(gate419inter0));
  nand2 gate1960(.a(gate419inter0), .b(s_154), .O(gate419inter1));
  and2  gate1961(.a(N1496), .b(N1459), .O(gate419inter2));
  inv1  gate1962(.a(s_154), .O(gate419inter3));
  inv1  gate1963(.a(s_155), .O(gate419inter4));
  nand2 gate1964(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1965(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1966(.a(N1459), .O(gate419inter7));
  inv1  gate1967(.a(N1496), .O(gate419inter8));
  nand2 gate1968(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1969(.a(s_155), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1970(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1971(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1972(.a(gate419inter12), .b(gate419inter1), .O(N1527));
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );

  xor2  gate979(.a(N1531), .b(N1484), .O(gate432inter0));
  nand2 gate980(.a(gate432inter0), .b(s_14), .O(gate432inter1));
  and2  gate981(.a(N1531), .b(N1484), .O(gate432inter2));
  inv1  gate982(.a(s_14), .O(gate432inter3));
  inv1  gate983(.a(s_15), .O(gate432inter4));
  nand2 gate984(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate985(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate986(.a(N1484), .O(gate432inter7));
  inv1  gate987(.a(N1531), .O(gate432inter8));
  nand2 gate988(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate989(.a(s_15), .b(gate432inter3), .O(gate432inter10));
  nor2  gate990(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate991(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate992(.a(gate432inter12), .b(gate432inter1), .O(N1567));

  xor2  gate1469(.a(N1532), .b(N1481), .O(gate433inter0));
  nand2 gate1470(.a(gate433inter0), .b(s_84), .O(gate433inter1));
  and2  gate1471(.a(N1532), .b(N1481), .O(gate433inter2));
  inv1  gate1472(.a(s_84), .O(gate433inter3));
  inv1  gate1473(.a(s_85), .O(gate433inter4));
  nand2 gate1474(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1475(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1476(.a(N1481), .O(gate433inter7));
  inv1  gate1477(.a(N1532), .O(gate433inter8));
  nand2 gate1478(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1479(.a(s_85), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1480(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1481(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1482(.a(gate433inter12), .b(gate433inter1), .O(N1568));
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );

  xor2  gate1847(.a(N893), .b(N1596), .O(gate462inter0));
  nand2 gate1848(.a(gate462inter0), .b(s_138), .O(gate462inter1));
  and2  gate1849(.a(N893), .b(N1596), .O(gate462inter2));
  inv1  gate1850(.a(s_138), .O(gate462inter3));
  inv1  gate1851(.a(s_139), .O(gate462inter4));
  nand2 gate1852(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1853(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1854(.a(N1596), .O(gate462inter7));
  inv1  gate1855(.a(N893), .O(gate462inter8));
  nand2 gate1856(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1857(.a(s_139), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1858(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1859(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1860(.a(gate462inter12), .b(gate462inter1), .O(N1671));
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );

  xor2  gate2239(.a(N1219), .b(N1609), .O(gate468inter0));
  nand2 gate2240(.a(gate468inter0), .b(s_194), .O(gate468inter1));
  and2  gate2241(.a(N1219), .b(N1609), .O(gate468inter2));
  inv1  gate2242(.a(s_194), .O(gate468inter3));
  inv1  gate2243(.a(s_195), .O(gate468inter4));
  nand2 gate2244(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2245(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2246(.a(N1609), .O(gate468inter7));
  inv1  gate2247(.a(N1219), .O(gate468inter8));
  nand2 gate2248(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2249(.a(s_195), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2250(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2251(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2252(.a(gate468inter12), .b(gate468inter1), .O(N1680));
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );

  xor2  gate2155(.a(N1672), .b(N643), .O(gate476inter0));
  nand2 gate2156(.a(gate476inter0), .b(s_182), .O(gate476inter1));
  and2  gate2157(.a(N1672), .b(N643), .O(gate476inter2));
  inv1  gate2158(.a(s_182), .O(gate476inter3));
  inv1  gate2159(.a(s_183), .O(gate476inter4));
  nand2 gate2160(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2161(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2162(.a(N643), .O(gate476inter7));
  inv1  gate2163(.a(N1672), .O(gate476inter8));
  nand2 gate2164(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2165(.a(s_183), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2166(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2167(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2168(.a(gate476inter12), .b(gate476inter1), .O(N1706));
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );

  xor2  gate1749(.a(N1593), .b(N1658), .O(gate486inter0));
  nand2 gate1750(.a(gate486inter0), .b(s_124), .O(gate486inter1));
  and2  gate1751(.a(N1593), .b(N1658), .O(gate486inter2));
  inv1  gate1752(.a(s_124), .O(gate486inter3));
  inv1  gate1753(.a(s_125), .O(gate486inter4));
  nand2 gate1754(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1755(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1756(.a(N1658), .O(gate486inter7));
  inv1  gate1757(.a(N1593), .O(gate486inter8));
  nand2 gate1758(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1759(.a(s_125), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1760(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1761(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1762(.a(gate486inter12), .b(gate486inter1), .O(N1720));
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );

  xor2  gate1091(.a(N1528), .b(N1685), .O(gate494inter0));
  nand2 gate1092(.a(gate494inter0), .b(s_30), .O(gate494inter1));
  and2  gate1093(.a(N1528), .b(N1685), .O(gate494inter2));
  inv1  gate1094(.a(s_30), .O(gate494inter3));
  inv1  gate1095(.a(s_31), .O(gate494inter4));
  nand2 gate1096(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1097(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1098(.a(N1685), .O(gate494inter7));
  inv1  gate1099(.a(N1528), .O(gate494inter8));
  nand2 gate1100(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1101(.a(s_31), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1102(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1103(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1104(.a(gate494inter12), .b(gate494inter1), .O(N1740));
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );

  xor2  gate1483(.a(N1711), .b(N1603), .O(gate498inter0));
  nand2 gate1484(.a(gate498inter0), .b(s_86), .O(gate498inter1));
  and2  gate1485(.a(N1711), .b(N1603), .O(gate498inter2));
  inv1  gate1486(.a(s_86), .O(gate498inter3));
  inv1  gate1487(.a(s_87), .O(gate498inter4));
  nand2 gate1488(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1489(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1490(.a(N1603), .O(gate498inter7));
  inv1  gate1491(.a(N1711), .O(gate498inter8));
  nand2 gate1492(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1493(.a(s_87), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1494(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1495(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1496(.a(gate498inter12), .b(gate498inter1), .O(N1747));
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate1021(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate1022(.a(gate503inter0), .b(s_20), .O(gate503inter1));
  and2  gate1023(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate1024(.a(s_20), .O(gate503inter3));
  inv1  gate1025(.a(s_21), .O(gate503inter4));
  nand2 gate1026(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1027(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1028(.a(N1697), .O(gate503inter7));
  inv1  gate1029(.a(N1727), .O(gate503inter8));
  nand2 gate1030(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1031(.a(s_21), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1032(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1033(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1034(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );

  xor2  gate895(.a(N1741), .b(N1472), .O(gate507inter0));
  nand2 gate896(.a(gate507inter0), .b(s_2), .O(gate507inter1));
  and2  gate897(.a(N1741), .b(N1472), .O(gate507inter2));
  inv1  gate898(.a(s_2), .O(gate507inter3));
  inv1  gate899(.a(s_3), .O(gate507inter4));
  nand2 gate900(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate901(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate902(.a(N1472), .O(gate507inter7));
  inv1  gate903(.a(N1741), .O(gate507inter8));
  nand2 gate904(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate905(.a(s_3), .b(gate507inter3), .O(gate507inter10));
  nor2  gate906(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate907(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate908(.a(gate507inter12), .b(gate507inter1), .O(N1769));

  xor2  gate1917(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate1918(.a(gate508inter0), .b(s_148), .O(gate508inter1));
  and2  gate1919(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate1920(.a(s_148), .O(gate508inter3));
  inv1  gate1921(.a(s_149), .O(gate508inter4));
  nand2 gate1922(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1923(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1924(.a(N1723), .O(gate508inter7));
  inv1  gate1925(.a(N1413), .O(gate508inter8));
  nand2 gate1926(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1927(.a(s_149), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1928(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1929(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1930(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1609(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1610(.a(gate513inter0), .b(s_104), .O(gate513inter1));
  and2  gate1611(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1612(.a(s_104), .O(gate513inter3));
  inv1  gate1613(.a(s_105), .O(gate513inter4));
  nand2 gate1614(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1615(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1616(.a(N1731), .O(gate513inter7));
  inv1  gate1617(.a(N1682), .O(gate513inter8));
  nand2 gate1618(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1619(.a(s_105), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1620(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1621(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1622(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );

  xor2  gate2211(.a(N1796), .b(N962), .O(gate536inter0));
  nand2 gate2212(.a(gate536inter0), .b(s_190), .O(gate536inter1));
  and2  gate2213(.a(N1796), .b(N962), .O(gate536inter2));
  inv1  gate2214(.a(s_190), .O(gate536inter3));
  inv1  gate2215(.a(s_191), .O(gate536inter4));
  nand2 gate2216(.a(gate536inter4), .b(gate536inter3), .O(gate536inter5));
  nor2  gate2217(.a(gate536inter5), .b(gate536inter2), .O(gate536inter6));
  inv1  gate2218(.a(N962), .O(gate536inter7));
  inv1  gate2219(.a(N1796), .O(gate536inter8));
  nand2 gate2220(.a(gate536inter8), .b(gate536inter7), .O(gate536inter9));
  nand2 gate2221(.a(s_191), .b(gate536inter3), .O(gate536inter10));
  nor2  gate2222(.a(gate536inter10), .b(gate536inter9), .O(gate536inter11));
  nor2  gate2223(.a(gate536inter11), .b(gate536inter6), .O(gate536inter12));
  nand2 gate2224(.a(gate536inter12), .b(gate536inter1), .O(N1825));
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );

  xor2  gate2071(.a(N1784), .b(N1809), .O(gate541inter0));
  nand2 gate2072(.a(gate541inter0), .b(s_170), .O(gate541inter1));
  and2  gate2073(.a(N1784), .b(N1809), .O(gate541inter2));
  inv1  gate2074(.a(s_170), .O(gate541inter3));
  inv1  gate2075(.a(s_171), .O(gate541inter4));
  nand2 gate2076(.a(gate541inter4), .b(gate541inter3), .O(gate541inter5));
  nor2  gate2077(.a(gate541inter5), .b(gate541inter2), .O(gate541inter6));
  inv1  gate2078(.a(N1809), .O(gate541inter7));
  inv1  gate2079(.a(N1784), .O(gate541inter8));
  nand2 gate2080(.a(gate541inter8), .b(gate541inter7), .O(gate541inter9));
  nand2 gate2081(.a(s_171), .b(gate541inter3), .O(gate541inter10));
  nor2  gate2082(.a(gate541inter10), .b(gate541inter9), .O(gate541inter11));
  nor2  gate2083(.a(gate541inter11), .b(gate541inter6), .O(gate541inter12));
  nand2 gate2084(.a(gate541inter12), .b(gate541inter1), .O(N1838));
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );

  xor2  gate1385(.a(N1825), .b(N1795), .O(gate545inter0));
  nand2 gate1386(.a(gate545inter0), .b(s_72), .O(gate545inter1));
  and2  gate1387(.a(N1825), .b(N1795), .O(gate545inter2));
  inv1  gate1388(.a(s_72), .O(gate545inter3));
  inv1  gate1389(.a(s_73), .O(gate545inter4));
  nand2 gate1390(.a(gate545inter4), .b(gate545inter3), .O(gate545inter5));
  nor2  gate1391(.a(gate545inter5), .b(gate545inter2), .O(gate545inter6));
  inv1  gate1392(.a(N1795), .O(gate545inter7));
  inv1  gate1393(.a(N1825), .O(gate545inter8));
  nand2 gate1394(.a(gate545inter8), .b(gate545inter7), .O(gate545inter9));
  nand2 gate1395(.a(s_73), .b(gate545inter3), .O(gate545inter10));
  nor2  gate1396(.a(gate545inter10), .b(gate545inter9), .O(gate545inter11));
  nor2  gate1397(.a(gate545inter11), .b(gate545inter6), .O(gate545inter12));
  nand2 gate1398(.a(gate545inter12), .b(gate545inter1), .O(N1850));
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );

  xor2  gate1455(.a(N1837), .b(N1808), .O(gate556inter0));
  nand2 gate1456(.a(gate556inter0), .b(s_82), .O(gate556inter1));
  and2  gate1457(.a(N1837), .b(N1808), .O(gate556inter2));
  inv1  gate1458(.a(s_82), .O(gate556inter3));
  inv1  gate1459(.a(s_83), .O(gate556inter4));
  nand2 gate1460(.a(gate556inter4), .b(gate556inter3), .O(gate556inter5));
  nor2  gate1461(.a(gate556inter5), .b(gate556inter2), .O(gate556inter6));
  inv1  gate1462(.a(N1808), .O(gate556inter7));
  inv1  gate1463(.a(N1837), .O(gate556inter8));
  nand2 gate1464(.a(gate556inter8), .b(gate556inter7), .O(gate556inter9));
  nand2 gate1465(.a(s_83), .b(gate556inter3), .O(gate556inter10));
  nor2  gate1466(.a(gate556inter10), .b(gate556inter9), .O(gate556inter11));
  nor2  gate1467(.a(gate556inter11), .b(gate556inter6), .O(gate556inter12));
  nand2 gate1468(.a(gate556inter12), .b(gate556inter1), .O(N1875));
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );

  xor2  gate1595(.a(N1852), .b(N1826), .O(gate561inter0));
  nand2 gate1596(.a(gate561inter0), .b(s_102), .O(gate561inter1));
  and2  gate1597(.a(N1852), .b(N1826), .O(gate561inter2));
  inv1  gate1598(.a(s_102), .O(gate561inter3));
  inv1  gate1599(.a(s_103), .O(gate561inter4));
  nand2 gate1600(.a(gate561inter4), .b(gate561inter3), .O(gate561inter5));
  nor2  gate1601(.a(gate561inter5), .b(gate561inter2), .O(gate561inter6));
  inv1  gate1602(.a(N1826), .O(gate561inter7));
  inv1  gate1603(.a(N1852), .O(gate561inter8));
  nand2 gate1604(.a(gate561inter8), .b(gate561inter7), .O(gate561inter9));
  nand2 gate1605(.a(s_103), .b(gate561inter3), .O(gate561inter10));
  nor2  gate1606(.a(gate561inter10), .b(gate561inter9), .O(gate561inter11));
  nor2  gate1607(.a(gate561inter11), .b(gate561inter6), .O(gate561inter12));
  nand2 gate1608(.a(gate561inter12), .b(gate561inter1), .O(N1884));

  xor2  gate1987(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate1988(.a(gate562inter0), .b(s_158), .O(gate562inter1));
  and2  gate1989(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate1990(.a(s_158), .O(gate562inter3));
  inv1  gate1991(.a(s_159), .O(gate562inter4));
  nand2 gate1992(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate1993(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate1994(.a(N1643), .O(gate562inter7));
  inv1  gate1995(.a(N1856), .O(gate562inter8));
  nand2 gate1996(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate1997(.a(s_159), .b(gate562inter3), .O(gate562inter10));
  nor2  gate1998(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate1999(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate2000(.a(gate562inter12), .b(gate562inter1), .O(N1885));
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate2281(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate2282(.a(gate565inter0), .b(s_200), .O(gate565inter1));
  and2  gate2283(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate2284(.a(s_200), .O(gate565inter3));
  inv1  gate2285(.a(s_201), .O(gate565inter4));
  nand2 gate2286(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate2287(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate2288(.a(N1838), .O(gate565inter7));
  inv1  gate2289(.a(N1785), .O(gate565inter8));
  nand2 gate2290(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate2291(.a(s_201), .b(gate565inter3), .O(gate565inter10));
  nor2  gate2292(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate2293(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate2294(.a(gate565inter12), .b(gate565inter1), .O(N1896));
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );

  xor2  gate1777(.a(N1885), .b(N1855), .O(gate572inter0));
  nand2 gate1778(.a(gate572inter0), .b(s_128), .O(gate572inter1));
  and2  gate1779(.a(N1885), .b(N1855), .O(gate572inter2));
  inv1  gate1780(.a(s_128), .O(gate572inter3));
  inv1  gate1781(.a(s_129), .O(gate572inter4));
  nand2 gate1782(.a(gate572inter4), .b(gate572inter3), .O(gate572inter5));
  nor2  gate1783(.a(gate572inter5), .b(gate572inter2), .O(gate572inter6));
  inv1  gate1784(.a(N1855), .O(gate572inter7));
  inv1  gate1785(.a(N1885), .O(gate572inter8));
  nand2 gate1786(.a(gate572inter8), .b(gate572inter7), .O(gate572inter9));
  nand2 gate1787(.a(s_129), .b(gate572inter3), .O(gate572inter10));
  nor2  gate1788(.a(gate572inter10), .b(gate572inter9), .O(gate572inter11));
  nor2  gate1789(.a(gate572inter11), .b(gate572inter6), .O(gate572inter12));
  nand2 gate1790(.a(gate572inter12), .b(gate572inter1), .O(N1913));
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );

  xor2  gate1357(.a(N1350), .b(N1953), .O(gate608inter0));
  nand2 gate1358(.a(gate608inter0), .b(s_68), .O(gate608inter1));
  and2  gate1359(.a(N1350), .b(N1953), .O(gate608inter2));
  inv1  gate1360(.a(s_68), .O(gate608inter3));
  inv1  gate1361(.a(s_69), .O(gate608inter4));
  nand2 gate1362(.a(gate608inter4), .b(gate608inter3), .O(gate608inter5));
  nor2  gate1363(.a(gate608inter5), .b(gate608inter2), .O(gate608inter6));
  inv1  gate1364(.a(N1953), .O(gate608inter7));
  inv1  gate1365(.a(N1350), .O(gate608inter8));
  nand2 gate1366(.a(gate608inter8), .b(gate608inter7), .O(gate608inter9));
  nand2 gate1367(.a(s_69), .b(gate608inter3), .O(gate608inter10));
  nor2  gate1368(.a(gate608inter10), .b(gate608inter9), .O(gate608inter11));
  nor2  gate1369(.a(gate608inter11), .b(gate608inter6), .O(gate608inter12));
  nand2 gate1370(.a(gate608inter12), .b(gate608inter1), .O(N2004));
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );

  xor2  gate1665(.a(N1978), .b(N670), .O(gate613inter0));
  nand2 gate1666(.a(gate613inter0), .b(s_112), .O(gate613inter1));
  and2  gate1667(.a(N1978), .b(N670), .O(gate613inter2));
  inv1  gate1668(.a(s_112), .O(gate613inter3));
  inv1  gate1669(.a(s_113), .O(gate613inter4));
  nand2 gate1670(.a(gate613inter4), .b(gate613inter3), .O(gate613inter5));
  nor2  gate1671(.a(gate613inter5), .b(gate613inter2), .O(gate613inter6));
  inv1  gate1672(.a(N670), .O(gate613inter7));
  inv1  gate1673(.a(N1978), .O(gate613inter8));
  nand2 gate1674(.a(gate613inter8), .b(gate613inter7), .O(gate613inter9));
  nand2 gate1675(.a(s_113), .b(gate613inter3), .O(gate613inter10));
  nor2  gate1676(.a(gate613inter10), .b(gate613inter9), .O(gate613inter11));
  nor2  gate1677(.a(gate613inter11), .b(gate613inter6), .O(gate613inter12));
  nand2 gate1678(.a(gate613inter12), .b(gate613inter1), .O(N2009));
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );

  xor2  gate1525(.a(N1923), .b(N1958), .O(gate616inter0));
  nand2 gate1526(.a(gate616inter0), .b(s_92), .O(gate616inter1));
  and2  gate1527(.a(N1923), .b(N1958), .O(gate616inter2));
  inv1  gate1528(.a(s_92), .O(gate616inter3));
  inv1  gate1529(.a(s_93), .O(gate616inter4));
  nand2 gate1530(.a(gate616inter4), .b(gate616inter3), .O(gate616inter5));
  nor2  gate1531(.a(gate616inter5), .b(gate616inter2), .O(gate616inter6));
  inv1  gate1532(.a(N1958), .O(gate616inter7));
  inv1  gate1533(.a(N1923), .O(gate616inter8));
  nand2 gate1534(.a(gate616inter8), .b(gate616inter7), .O(gate616inter9));
  nand2 gate1535(.a(s_93), .b(gate616inter3), .O(gate616inter10));
  nor2  gate1536(.a(gate616inter10), .b(gate616inter9), .O(gate616inter11));
  nor2  gate1537(.a(gate616inter11), .b(gate616inter6), .O(gate616inter12));
  nand2 gate1538(.a(gate616inter12), .b(gate616inter1), .O(N2014));
inv1 gate617( .a(N1961), .O(N2015) );

  xor2  gate937(.a(N1635), .b(N1961), .O(gate618inter0));
  nand2 gate938(.a(gate618inter0), .b(s_8), .O(gate618inter1));
  and2  gate939(.a(N1635), .b(N1961), .O(gate618inter2));
  inv1  gate940(.a(s_8), .O(gate618inter3));
  inv1  gate941(.a(s_9), .O(gate618inter4));
  nand2 gate942(.a(gate618inter4), .b(gate618inter3), .O(gate618inter5));
  nor2  gate943(.a(gate618inter5), .b(gate618inter2), .O(gate618inter6));
  inv1  gate944(.a(N1961), .O(gate618inter7));
  inv1  gate945(.a(N1635), .O(gate618inter8));
  nand2 gate946(.a(gate618inter8), .b(gate618inter7), .O(gate618inter9));
  nand2 gate947(.a(s_9), .b(gate618inter3), .O(gate618inter10));
  nor2  gate948(.a(gate618inter10), .b(gate618inter9), .O(gate618inter11));
  nor2  gate949(.a(gate618inter11), .b(gate618inter6), .O(gate618inter12));
  nand2 gate950(.a(gate618inter12), .b(gate618inter1), .O(N2016));
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );

  xor2  gate2253(.a(N1591), .b(N1987), .O(gate623inter0));
  nand2 gate2254(.a(gate623inter0), .b(s_196), .O(gate623inter1));
  and2  gate2255(.a(N1591), .b(N1987), .O(gate623inter2));
  inv1  gate2256(.a(s_196), .O(gate623inter3));
  inv1  gate2257(.a(s_197), .O(gate623inter4));
  nand2 gate2258(.a(gate623inter4), .b(gate623inter3), .O(gate623inter5));
  nor2  gate2259(.a(gate623inter5), .b(gate623inter2), .O(gate623inter6));
  inv1  gate2260(.a(N1987), .O(gate623inter7));
  inv1  gate2261(.a(N1591), .O(gate623inter8));
  nand2 gate2262(.a(gate623inter8), .b(gate623inter7), .O(gate623inter9));
  nand2 gate2263(.a(s_197), .b(gate623inter3), .O(gate623inter10));
  nor2  gate2264(.a(gate623inter10), .b(gate623inter9), .O(gate623inter11));
  nor2  gate2265(.a(gate623inter11), .b(gate623inter6), .O(gate623inter12));
  nand2 gate2266(.a(gate623inter12), .b(gate623inter1), .O(N2022));

  xor2  gate1105(.a(N2002), .b(N1440), .O(gate624inter0));
  nand2 gate1106(.a(gate624inter0), .b(s_32), .O(gate624inter1));
  and2  gate1107(.a(N2002), .b(N1440), .O(gate624inter2));
  inv1  gate1108(.a(s_32), .O(gate624inter3));
  inv1  gate1109(.a(s_33), .O(gate624inter4));
  nand2 gate1110(.a(gate624inter4), .b(gate624inter3), .O(gate624inter5));
  nor2  gate1111(.a(gate624inter5), .b(gate624inter2), .O(gate624inter6));
  inv1  gate1112(.a(N1440), .O(gate624inter7));
  inv1  gate1113(.a(N2002), .O(gate624inter8));
  nand2 gate1114(.a(gate624inter8), .b(gate624inter7), .O(gate624inter9));
  nand2 gate1115(.a(s_33), .b(gate624inter3), .O(gate624inter10));
  nor2  gate1116(.a(gate624inter10), .b(gate624inter9), .O(gate624inter11));
  nor2  gate1117(.a(gate624inter11), .b(gate624inter6), .O(gate624inter12));
  nand2 gate1118(.a(gate624inter12), .b(gate624inter1), .O(N2023));
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );

  xor2  gate1147(.a(N2007), .b(N1258), .O(gate626inter0));
  nand2 gate1148(.a(gate626inter0), .b(s_38), .O(gate626inter1));
  and2  gate1149(.a(N2007), .b(N1258), .O(gate626inter2));
  inv1  gate1150(.a(s_38), .O(gate626inter3));
  inv1  gate1151(.a(s_39), .O(gate626inter4));
  nand2 gate1152(.a(gate626inter4), .b(gate626inter3), .O(gate626inter5));
  nor2  gate1153(.a(gate626inter5), .b(gate626inter2), .O(gate626inter6));
  inv1  gate1154(.a(N1258), .O(gate626inter7));
  inv1  gate1155(.a(N2007), .O(gate626inter8));
  nand2 gate1156(.a(gate626inter8), .b(gate626inter7), .O(gate626inter9));
  nand2 gate1157(.a(s_39), .b(gate626inter3), .O(gate626inter10));
  nor2  gate1158(.a(gate626inter10), .b(gate626inter9), .O(gate626inter11));
  nor2  gate1159(.a(gate626inter11), .b(gate626inter6), .O(gate626inter12));
  nand2 gate1160(.a(gate626inter12), .b(gate626inter1), .O(N2025));
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );

  xor2  gate1133(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1134(.a(gate628inter0), .b(s_36), .O(gate628inter1));
  and2  gate1135(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1136(.a(s_36), .O(gate628inter3));
  inv1  gate1137(.a(s_37), .O(gate628inter4));
  nand2 gate1138(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1139(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1140(.a(N1977), .O(gate628inter7));
  inv1  gate1141(.a(N2009), .O(gate628inter8));
  nand2 gate1142(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1143(.a(s_37), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1144(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1145(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1146(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );

  xor2  gate1511(.a(N2015), .b(N1571), .O(gate632inter0));
  nand2 gate1512(.a(gate632inter0), .b(s_90), .O(gate632inter1));
  and2  gate1513(.a(N2015), .b(N1571), .O(gate632inter2));
  inv1  gate1514(.a(s_90), .O(gate632inter3));
  inv1  gate1515(.a(s_91), .O(gate632inter4));
  nand2 gate1516(.a(gate632inter4), .b(gate632inter3), .O(gate632inter5));
  nor2  gate1517(.a(gate632inter5), .b(gate632inter2), .O(gate632inter6));
  inv1  gate1518(.a(N1571), .O(gate632inter7));
  inv1  gate1519(.a(N2015), .O(gate632inter8));
  nand2 gate1520(.a(gate632inter8), .b(gate632inter7), .O(gate632inter9));
  nand2 gate1521(.a(s_91), .b(gate632inter3), .O(gate632inter10));
  nor2  gate1522(.a(gate632inter10), .b(gate632inter9), .O(gate632inter11));
  nor2  gate1523(.a(gate632inter11), .b(gate632inter6), .O(gate632inter12));
  nand2 gate1524(.a(gate632inter12), .b(gate632inter1), .O(N2037));

  xor2  gate1315(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate1316(.a(gate633inter0), .b(s_62), .O(gate633inter1));
  and2  gate1317(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate1318(.a(s_62), .O(gate633inter3));
  inv1  gate1319(.a(s_63), .O(gate633inter4));
  nand2 gate1320(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate1321(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate1322(.a(N2020), .O(gate633inter7));
  inv1  gate1323(.a(N2000), .O(gate633inter8));
  nand2 gate1324(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate1325(.a(s_63), .b(gate633inter3), .O(gate633inter10));
  nor2  gate1326(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate1327(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate1328(.a(gate633inter12), .b(gate633inter1), .O(N2038));
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );

  xor2  gate1903(.a(N2016), .b(N2037), .O(gate640inter0));
  nand2 gate1904(.a(gate640inter0), .b(s_146), .O(gate640inter1));
  and2  gate1905(.a(N2016), .b(N2037), .O(gate640inter2));
  inv1  gate1906(.a(s_146), .O(gate640inter3));
  inv1  gate1907(.a(s_147), .O(gate640inter4));
  nand2 gate1908(.a(gate640inter4), .b(gate640inter3), .O(gate640inter5));
  nor2  gate1909(.a(gate640inter5), .b(gate640inter2), .O(gate640inter6));
  inv1  gate1910(.a(N2037), .O(gate640inter7));
  inv1  gate1911(.a(N2016), .O(gate640inter8));
  nand2 gate1912(.a(gate640inter8), .b(gate640inter7), .O(gate640inter9));
  nand2 gate1913(.a(s_147), .b(gate640inter3), .O(gate640inter10));
  nor2  gate1914(.a(gate640inter10), .b(gate640inter9), .O(gate640inter11));
  nor2  gate1915(.a(gate640inter11), .b(gate640inter6), .O(gate640inter12));
  nand2 gate1916(.a(gate640inter12), .b(gate640inter1), .O(N2055));
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );

  xor2  gate2113(.a(N915), .b(N2151), .O(gate663inter0));
  nand2 gate2114(.a(gate663inter0), .b(s_176), .O(gate663inter1));
  and2  gate2115(.a(N915), .b(N2151), .O(gate663inter2));
  inv1  gate2116(.a(s_176), .O(gate663inter3));
  inv1  gate2117(.a(s_177), .O(gate663inter4));
  nand2 gate2118(.a(gate663inter4), .b(gate663inter3), .O(gate663inter5));
  nor2  gate2119(.a(gate663inter5), .b(gate663inter2), .O(gate663inter6));
  inv1  gate2120(.a(N2151), .O(gate663inter7));
  inv1  gate2121(.a(N915), .O(gate663inter8));
  nand2 gate2122(.a(gate663inter8), .b(gate663inter7), .O(gate663inter9));
  nand2 gate2123(.a(s_177), .b(gate663inter3), .O(gate663inter10));
  nor2  gate2124(.a(gate663inter10), .b(gate663inter9), .O(gate663inter11));
  nor2  gate2125(.a(gate663inter11), .b(gate663inter6), .O(gate663inter12));
  nand2 gate2126(.a(gate663inter12), .b(gate663inter1), .O(N2214));
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );

  xor2  gate965(.a(N2227), .b(N661), .O(gate679inter0));
  nand2 gate966(.a(gate679inter0), .b(s_12), .O(gate679inter1));
  and2  gate967(.a(N2227), .b(N661), .O(gate679inter2));
  inv1  gate968(.a(s_12), .O(gate679inter3));
  inv1  gate969(.a(s_13), .O(gate679inter4));
  nand2 gate970(.a(gate679inter4), .b(gate679inter3), .O(gate679inter5));
  nor2  gate971(.a(gate679inter5), .b(gate679inter2), .O(gate679inter6));
  inv1  gate972(.a(N661), .O(gate679inter7));
  inv1  gate973(.a(N2227), .O(gate679inter8));
  nand2 gate974(.a(gate679inter8), .b(gate679inter7), .O(gate679inter9));
  nand2 gate975(.a(s_13), .b(gate679inter3), .O(gate679inter10));
  nor2  gate976(.a(gate679inter10), .b(gate679inter9), .O(gate679inter11));
  nor2  gate977(.a(gate679inter11), .b(gate679inter6), .O(gate679inter12));
  nand2 gate978(.a(gate679inter12), .b(gate679inter1), .O(N2234));
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );

  xor2  gate1763(.a(N2231), .b(N2216), .O(gate682inter0));
  nand2 gate1764(.a(gate682inter0), .b(s_126), .O(gate682inter1));
  and2  gate1765(.a(N2231), .b(N2216), .O(gate682inter2));
  inv1  gate1766(.a(s_126), .O(gate682inter3));
  inv1  gate1767(.a(s_127), .O(gate682inter4));
  nand2 gate1768(.a(gate682inter4), .b(gate682inter3), .O(gate682inter5));
  nor2  gate1769(.a(gate682inter5), .b(gate682inter2), .O(gate682inter6));
  inv1  gate1770(.a(N2216), .O(gate682inter7));
  inv1  gate1771(.a(N2231), .O(gate682inter8));
  nand2 gate1772(.a(gate682inter8), .b(gate682inter7), .O(gate682inter9));
  nand2 gate1773(.a(s_127), .b(gate682inter3), .O(gate682inter10));
  nor2  gate1774(.a(gate682inter10), .b(gate682inter9), .O(gate682inter11));
  nor2  gate1775(.a(gate682inter11), .b(gate682inter6), .O(gate682inter12));
  nand2 gate1776(.a(gate682inter12), .b(gate682inter1), .O(N2237));
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );

  xor2  gate1539(.a(N2235), .b(N2228), .O(gate686inter0));
  nand2 gate1540(.a(gate686inter0), .b(s_94), .O(gate686inter1));
  and2  gate1541(.a(N2235), .b(N2228), .O(gate686inter2));
  inv1  gate1542(.a(s_94), .O(gate686inter3));
  inv1  gate1543(.a(s_95), .O(gate686inter4));
  nand2 gate1544(.a(gate686inter4), .b(gate686inter3), .O(gate686inter5));
  nor2  gate1545(.a(gate686inter5), .b(gate686inter2), .O(gate686inter6));
  inv1  gate1546(.a(N2228), .O(gate686inter7));
  inv1  gate1547(.a(N2235), .O(gate686inter8));
  nand2 gate1548(.a(gate686inter8), .b(gate686inter7), .O(gate686inter9));
  nand2 gate1549(.a(s_95), .b(gate686inter3), .O(gate686inter10));
  nor2  gate1550(.a(gate686inter10), .b(gate686inter9), .O(gate686inter11));
  nor2  gate1551(.a(gate686inter11), .b(gate686inter6), .O(gate686inter12));
  nand2 gate1552(.a(gate686inter12), .b(gate686inter1), .O(N2245));
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );

  xor2  gate1077(.a(N535), .b(N2561), .O(gate752inter0));
  nand2 gate1078(.a(gate752inter0), .b(s_28), .O(gate752inter1));
  and2  gate1079(.a(N535), .b(N2561), .O(gate752inter2));
  inv1  gate1080(.a(s_28), .O(gate752inter3));
  inv1  gate1081(.a(s_29), .O(gate752inter4));
  nand2 gate1082(.a(gate752inter4), .b(gate752inter3), .O(gate752inter5));
  nor2  gate1083(.a(gate752inter5), .b(gate752inter2), .O(gate752inter6));
  inv1  gate1084(.a(N2561), .O(gate752inter7));
  inv1  gate1085(.a(N535), .O(gate752inter8));
  nand2 gate1086(.a(gate752inter8), .b(gate752inter7), .O(gate752inter9));
  nand2 gate1087(.a(s_29), .b(gate752inter3), .O(gate752inter10));
  nor2  gate1088(.a(gate752inter10), .b(gate752inter9), .O(gate752inter11));
  nor2  gate1089(.a(gate752inter11), .b(gate752inter6), .O(gate752inter12));
  nand2 gate1090(.a(gate752inter12), .b(gate752inter1), .O(N2671));
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );

  xor2  gate923(.a(N548), .b(N2573), .O(gate760inter0));
  nand2 gate924(.a(gate760inter0), .b(s_6), .O(gate760inter1));
  and2  gate925(.a(N548), .b(N2573), .O(gate760inter2));
  inv1  gate926(.a(s_6), .O(gate760inter3));
  inv1  gate927(.a(s_7), .O(gate760inter4));
  nand2 gate928(.a(gate760inter4), .b(gate760inter3), .O(gate760inter5));
  nor2  gate929(.a(gate760inter5), .b(gate760inter2), .O(gate760inter6));
  inv1  gate930(.a(N2573), .O(gate760inter7));
  inv1  gate931(.a(N548), .O(gate760inter8));
  nand2 gate932(.a(gate760inter8), .b(gate760inter7), .O(gate760inter9));
  nand2 gate933(.a(s_7), .b(gate760inter3), .O(gate760inter10));
  nor2  gate934(.a(gate760inter10), .b(gate760inter9), .O(gate760inter11));
  nor2  gate935(.a(gate760inter11), .b(gate760inter6), .O(gate760inter12));
  nand2 gate936(.a(gate760inter12), .b(gate760inter1), .O(N2688));
inv1 gate761( .a(N2573), .O(N2689) );

  xor2  gate993(.a(N549), .b(N2576), .O(gate762inter0));
  nand2 gate994(.a(gate762inter0), .b(s_16), .O(gate762inter1));
  and2  gate995(.a(N549), .b(N2576), .O(gate762inter2));
  inv1  gate996(.a(s_16), .O(gate762inter3));
  inv1  gate997(.a(s_17), .O(gate762inter4));
  nand2 gate998(.a(gate762inter4), .b(gate762inter3), .O(gate762inter5));
  nor2  gate999(.a(gate762inter5), .b(gate762inter2), .O(gate762inter6));
  inv1  gate1000(.a(N2576), .O(gate762inter7));
  inv1  gate1001(.a(N549), .O(gate762inter8));
  nand2 gate1002(.a(gate762inter8), .b(gate762inter7), .O(gate762inter9));
  nand2 gate1003(.a(s_17), .b(gate762inter3), .O(gate762inter10));
  nor2  gate1004(.a(gate762inter10), .b(gate762inter9), .O(gate762inter11));
  nor2  gate1005(.a(gate762inter11), .b(gate762inter6), .O(gate762inter12));
  nand2 gate1006(.a(gate762inter12), .b(gate762inter1), .O(N2690));
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );

  xor2  gate1931(.a(N2672), .b(N346), .O(gate766inter0));
  nand2 gate1932(.a(gate766inter0), .b(s_150), .O(gate766inter1));
  and2  gate1933(.a(N2672), .b(N346), .O(gate766inter2));
  inv1  gate1934(.a(s_150), .O(gate766inter3));
  inv1  gate1935(.a(s_151), .O(gate766inter4));
  nand2 gate1936(.a(gate766inter4), .b(gate766inter3), .O(gate766inter5));
  nor2  gate1937(.a(gate766inter5), .b(gate766inter2), .O(gate766inter6));
  inv1  gate1938(.a(N346), .O(gate766inter7));
  inv1  gate1939(.a(N2672), .O(gate766inter8));
  nand2 gate1940(.a(gate766inter8), .b(gate766inter7), .O(gate766inter9));
  nand2 gate1941(.a(s_151), .b(gate766inter3), .O(gate766inter10));
  nor2  gate1942(.a(gate766inter10), .b(gate766inter9), .O(gate766inter11));
  nor2  gate1943(.a(gate766inter11), .b(gate766inter6), .O(gate766inter12));
  nand2 gate1944(.a(gate766inter12), .b(gate766inter1), .O(N2721));
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );

  xor2  gate1259(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate1260(.a(gate768inter0), .b(s_54), .O(gate768inter1));
  and2  gate1261(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate1262(.a(s_54), .O(gate768inter3));
  inv1  gate1263(.a(s_55), .O(gate768inter4));
  nand2 gate1264(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate1265(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate1266(.a(N352), .O(gate768inter7));
  inv1  gate1267(.a(N2676), .O(gate768inter8));
  nand2 gate1268(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate1269(.a(s_55), .b(gate768inter3), .O(gate768inter10));
  nor2  gate1270(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate1271(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate1272(.a(gate768inter12), .b(gate768inter1), .O(N2723));
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );

  xor2  gate1721(.a(N539), .b(N2642), .O(gate771inter0));
  nand2 gate1722(.a(gate771inter0), .b(s_120), .O(gate771inter1));
  and2  gate1723(.a(N539), .b(N2642), .O(gate771inter2));
  inv1  gate1724(.a(s_120), .O(gate771inter3));
  inv1  gate1725(.a(s_121), .O(gate771inter4));
  nand2 gate1726(.a(gate771inter4), .b(gate771inter3), .O(gate771inter5));
  nor2  gate1727(.a(gate771inter5), .b(gate771inter2), .O(gate771inter6));
  inv1  gate1728(.a(N2642), .O(gate771inter7));
  inv1  gate1729(.a(N539), .O(gate771inter8));
  nand2 gate1730(.a(gate771inter8), .b(gate771inter7), .O(gate771inter9));
  nand2 gate1731(.a(s_121), .b(gate771inter3), .O(gate771inter10));
  nor2  gate1732(.a(gate771inter10), .b(gate771inter9), .O(gate771inter11));
  nor2  gate1733(.a(gate771inter11), .b(gate771inter6), .O(gate771inter12));
  nand2 gate1734(.a(gate771inter12), .b(gate771inter1), .O(N2726));
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );

  xor2  gate1063(.a(N544), .b(N2655), .O(gate780inter0));
  nand2 gate1064(.a(gate780inter0), .b(s_26), .O(gate780inter1));
  and2  gate1065(.a(N544), .b(N2655), .O(gate780inter2));
  inv1  gate1066(.a(s_26), .O(gate780inter3));
  inv1  gate1067(.a(s_27), .O(gate780inter4));
  nand2 gate1068(.a(gate780inter4), .b(gate780inter3), .O(gate780inter5));
  nor2  gate1069(.a(gate780inter5), .b(gate780inter2), .O(gate780inter6));
  inv1  gate1070(.a(N2655), .O(gate780inter7));
  inv1  gate1071(.a(N544), .O(gate780inter8));
  nand2 gate1072(.a(gate780inter8), .b(gate780inter7), .O(gate780inter9));
  nand2 gate1073(.a(s_27), .b(gate780inter3), .O(gate780inter10));
  nor2  gate1074(.a(gate780inter10), .b(gate780inter9), .O(gate780inter11));
  nor2  gate1075(.a(gate780inter11), .b(gate780inter6), .O(gate780inter12));
  nand2 gate1076(.a(gate780inter12), .b(gate780inter1), .O(N2735));
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );

  xor2  gate1273(.a(N2723), .b(N2675), .O(gate797inter0));
  nand2 gate1274(.a(gate797inter0), .b(s_56), .O(gate797inter1));
  and2  gate1275(.a(N2723), .b(N2675), .O(gate797inter2));
  inv1  gate1276(.a(s_56), .O(gate797inter3));
  inv1  gate1277(.a(s_57), .O(gate797inter4));
  nand2 gate1278(.a(gate797inter4), .b(gate797inter3), .O(gate797inter5));
  nor2  gate1279(.a(gate797inter5), .b(gate797inter2), .O(gate797inter6));
  inv1  gate1280(.a(N2675), .O(gate797inter7));
  inv1  gate1281(.a(N2723), .O(gate797inter8));
  nand2 gate1282(.a(gate797inter8), .b(gate797inter7), .O(gate797inter9));
  nand2 gate1283(.a(s_57), .b(gate797inter3), .O(gate797inter10));
  nor2  gate1284(.a(gate797inter10), .b(gate797inter9), .O(gate797inter11));
  nor2  gate1285(.a(gate797inter11), .b(gate797inter6), .O(gate797inter12));
  nand2 gate1286(.a(gate797inter12), .b(gate797inter1), .O(N2756));
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );

  xor2  gate2057(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate2058(.a(gate799inter0), .b(s_168), .O(gate799inter1));
  and2  gate2059(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate2060(.a(s_168), .O(gate799inter3));
  inv1  gate2061(.a(s_169), .O(gate799inter4));
  nand2 gate2062(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate2063(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate2064(.a(N358), .O(gate799inter7));
  inv1  gate2065(.a(N2727), .O(gate799inter8));
  nand2 gate2066(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate2067(.a(s_169), .b(gate799inter3), .O(gate799inter10));
  nor2  gate2068(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate2069(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate2070(.a(gate799inter12), .b(gate799inter1), .O(N2758));
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );

  xor2  gate2099(.a(N2733), .b(N367), .O(gate802inter0));
  nand2 gate2100(.a(gate802inter0), .b(s_174), .O(gate802inter1));
  and2  gate2101(.a(N2733), .b(N367), .O(gate802inter2));
  inv1  gate2102(.a(s_174), .O(gate802inter3));
  inv1  gate2103(.a(s_175), .O(gate802inter4));
  nand2 gate2104(.a(gate802inter4), .b(gate802inter3), .O(gate802inter5));
  nor2  gate2105(.a(gate802inter5), .b(gate802inter2), .O(gate802inter6));
  inv1  gate2106(.a(N367), .O(gate802inter7));
  inv1  gate2107(.a(N2733), .O(gate802inter8));
  nand2 gate2108(.a(gate802inter8), .b(gate802inter7), .O(gate802inter9));
  nand2 gate2109(.a(s_175), .b(gate802inter3), .O(gate802inter10));
  nor2  gate2110(.a(gate802inter10), .b(gate802inter9), .O(gate802inter11));
  nor2  gate2111(.a(gate802inter11), .b(gate802inter6), .O(gate802inter12));
  nand2 gate2112(.a(gate802inter12), .b(gate802inter1), .O(N2761));
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );

  xor2  gate1203(.a(N2736), .b(N373), .O(gate804inter0));
  nand2 gate1204(.a(gate804inter0), .b(s_46), .O(gate804inter1));
  and2  gate1205(.a(N2736), .b(N373), .O(gate804inter2));
  inv1  gate1206(.a(s_46), .O(gate804inter3));
  inv1  gate1207(.a(s_47), .O(gate804inter4));
  nand2 gate1208(.a(gate804inter4), .b(gate804inter3), .O(gate804inter5));
  nor2  gate1209(.a(gate804inter5), .b(gate804inter2), .O(gate804inter6));
  inv1  gate1210(.a(N373), .O(gate804inter7));
  inv1  gate1211(.a(N2736), .O(gate804inter8));
  nand2 gate1212(.a(gate804inter8), .b(gate804inter7), .O(gate804inter9));
  nand2 gate1213(.a(s_47), .b(gate804inter3), .O(gate804inter10));
  nor2  gate1214(.a(gate804inter10), .b(gate804inter9), .O(gate804inter11));
  nor2  gate1215(.a(gate804inter11), .b(gate804inter6), .O(gate804inter12));
  nand2 gate1216(.a(gate804inter12), .b(gate804inter1), .O(N2763));

  xor2  gate1301(.a(N2738), .b(N376), .O(gate805inter0));
  nand2 gate1302(.a(gate805inter0), .b(s_60), .O(gate805inter1));
  and2  gate1303(.a(N2738), .b(N376), .O(gate805inter2));
  inv1  gate1304(.a(s_60), .O(gate805inter3));
  inv1  gate1305(.a(s_61), .O(gate805inter4));
  nand2 gate1306(.a(gate805inter4), .b(gate805inter3), .O(gate805inter5));
  nor2  gate1307(.a(gate805inter5), .b(gate805inter2), .O(gate805inter6));
  inv1  gate1308(.a(N376), .O(gate805inter7));
  inv1  gate1309(.a(N2738), .O(gate805inter8));
  nand2 gate1310(.a(gate805inter8), .b(gate805inter7), .O(gate805inter9));
  nand2 gate1311(.a(s_61), .b(gate805inter3), .O(gate805inter10));
  nor2  gate1312(.a(gate805inter10), .b(gate805inter9), .O(gate805inter11));
  nor2  gate1313(.a(gate805inter11), .b(gate805inter6), .O(gate805inter12));
  nand2 gate1314(.a(gate805inter12), .b(gate805inter1), .O(N2764));

  xor2  gate1833(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate1834(.a(gate806inter0), .b(s_136), .O(gate806inter1));
  and2  gate1835(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate1836(.a(s_136), .O(gate806inter3));
  inv1  gate1837(.a(s_137), .O(gate806inter4));
  nand2 gate1838(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate1839(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate1840(.a(N379), .O(gate806inter7));
  inv1  gate1841(.a(N2740), .O(gate806inter8));
  nand2 gate1842(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate1843(.a(s_137), .b(gate806inter3), .O(gate806inter10));
  nor2  gate1844(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate1845(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate1846(.a(gate806inter12), .b(gate806inter1), .O(N2765));
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );

  xor2  gate1343(.a(N2757), .b(N2724), .O(gate812inter0));
  nand2 gate1344(.a(gate812inter0), .b(s_66), .O(gate812inter1));
  and2  gate1345(.a(N2757), .b(N2724), .O(gate812inter2));
  inv1  gate1346(.a(s_66), .O(gate812inter3));
  inv1  gate1347(.a(s_67), .O(gate812inter4));
  nand2 gate1348(.a(gate812inter4), .b(gate812inter3), .O(gate812inter5));
  nor2  gate1349(.a(gate812inter5), .b(gate812inter2), .O(gate812inter6));
  inv1  gate1350(.a(N2724), .O(gate812inter7));
  inv1  gate1351(.a(N2757), .O(gate812inter8));
  nand2 gate1352(.a(gate812inter8), .b(gate812inter7), .O(gate812inter9));
  nand2 gate1353(.a(s_67), .b(gate812inter3), .O(gate812inter10));
  nor2  gate1354(.a(gate812inter10), .b(gate812inter9), .O(gate812inter11));
  nor2  gate1355(.a(gate812inter11), .b(gate812inter6), .O(gate812inter12));
  nand2 gate1356(.a(gate812inter12), .b(gate812inter1), .O(N2779));
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );

  xor2  gate1553(.a(N2764), .b(N2737), .O(gate818inter0));
  nand2 gate1554(.a(gate818inter0), .b(s_96), .O(gate818inter1));
  and2  gate1555(.a(N2764), .b(N2737), .O(gate818inter2));
  inv1  gate1556(.a(s_96), .O(gate818inter3));
  inv1  gate1557(.a(s_97), .O(gate818inter4));
  nand2 gate1558(.a(gate818inter4), .b(gate818inter3), .O(gate818inter5));
  nor2  gate1559(.a(gate818inter5), .b(gate818inter2), .O(gate818inter6));
  inv1  gate1560(.a(N2737), .O(gate818inter7));
  inv1  gate1561(.a(N2764), .O(gate818inter8));
  nand2 gate1562(.a(gate818inter8), .b(gate818inter7), .O(gate818inter9));
  nand2 gate1563(.a(s_97), .b(gate818inter3), .O(gate818inter10));
  nor2  gate1564(.a(gate818inter10), .b(gate818inter9), .O(gate818inter11));
  nor2  gate1565(.a(gate818inter11), .b(gate818inter6), .O(gate818inter12));
  nand2 gate1566(.a(gate818inter12), .b(gate818inter1), .O(N2785));
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );

  xor2  gate1007(.a(N2018), .b(N2773), .O(gate824inter0));
  nand2 gate1008(.a(gate824inter0), .b(s_18), .O(gate824inter1));
  and2  gate1009(.a(N2018), .b(N2773), .O(gate824inter2));
  inv1  gate1010(.a(s_18), .O(gate824inter3));
  inv1  gate1011(.a(s_19), .O(gate824inter4));
  nand2 gate1012(.a(gate824inter4), .b(gate824inter3), .O(gate824inter5));
  nor2  gate1013(.a(gate824inter5), .b(gate824inter2), .O(gate824inter6));
  inv1  gate1014(.a(N2773), .O(gate824inter7));
  inv1  gate1015(.a(N2018), .O(gate824inter8));
  nand2 gate1016(.a(gate824inter8), .b(gate824inter7), .O(gate824inter9));
  nand2 gate1017(.a(s_19), .b(gate824inter3), .O(gate824inter10));
  nor2  gate1018(.a(gate824inter10), .b(gate824inter9), .O(gate824inter11));
  nor2  gate1019(.a(gate824inter11), .b(gate824inter6), .O(gate824inter12));
  nand2 gate1020(.a(gate824inter12), .b(gate824inter1), .O(N2807));
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );

  xor2  gate1119(.a(N2808), .b(N1965), .O(gate834inter0));
  nand2 gate1120(.a(gate834inter0), .b(s_34), .O(gate834inter1));
  and2  gate1121(.a(N2808), .b(N1965), .O(gate834inter2));
  inv1  gate1122(.a(s_34), .O(gate834inter3));
  inv1  gate1123(.a(s_35), .O(gate834inter4));
  nand2 gate1124(.a(gate834inter4), .b(gate834inter3), .O(gate834inter5));
  nor2  gate1125(.a(gate834inter5), .b(gate834inter2), .O(gate834inter6));
  inv1  gate1126(.a(N1965), .O(gate834inter7));
  inv1  gate1127(.a(N2808), .O(gate834inter8));
  nand2 gate1128(.a(gate834inter8), .b(gate834inter7), .O(gate834inter9));
  nand2 gate1129(.a(s_35), .b(gate834inter3), .O(gate834inter10));
  nor2  gate1130(.a(gate834inter10), .b(gate834inter9), .O(gate834inter11));
  nor2  gate1131(.a(gate834inter11), .b(gate834inter6), .O(gate834inter12));
  nand2 gate1132(.a(gate834inter12), .b(gate834inter1), .O(N2827));

  xor2  gate1567(.a(N2810), .b(N1968), .O(gate835inter0));
  nand2 gate1568(.a(gate835inter0), .b(s_98), .O(gate835inter1));
  and2  gate1569(.a(N2810), .b(N1968), .O(gate835inter2));
  inv1  gate1570(.a(s_98), .O(gate835inter3));
  inv1  gate1571(.a(s_99), .O(gate835inter4));
  nand2 gate1572(.a(gate835inter4), .b(gate835inter3), .O(gate835inter5));
  nor2  gate1573(.a(gate835inter5), .b(gate835inter2), .O(gate835inter6));
  inv1  gate1574(.a(N1968), .O(gate835inter7));
  inv1  gate1575(.a(N2810), .O(gate835inter8));
  nand2 gate1576(.a(gate835inter8), .b(gate835inter7), .O(gate835inter9));
  nand2 gate1577(.a(s_99), .b(gate835inter3), .O(gate835inter10));
  nor2  gate1578(.a(gate835inter10), .b(gate835inter9), .O(gate835inter11));
  nor2  gate1579(.a(gate835inter11), .b(gate835inter6), .O(gate835inter12));
  nand2 gate1580(.a(gate835inter12), .b(gate835inter1), .O(N2828));
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );

  xor2  gate1875(.a(N2827), .b(N2807), .O(gate837inter0));
  nand2 gate1876(.a(gate837inter0), .b(s_142), .O(gate837inter1));
  and2  gate1877(.a(N2827), .b(N2807), .O(gate837inter2));
  inv1  gate1878(.a(s_142), .O(gate837inter3));
  inv1  gate1879(.a(s_143), .O(gate837inter4));
  nand2 gate1880(.a(gate837inter4), .b(gate837inter3), .O(gate837inter5));
  nor2  gate1881(.a(gate837inter5), .b(gate837inter2), .O(gate837inter6));
  inv1  gate1882(.a(N2807), .O(gate837inter7));
  inv1  gate1883(.a(N2827), .O(gate837inter8));
  nand2 gate1884(.a(gate837inter8), .b(gate837inter7), .O(gate837inter9));
  nand2 gate1885(.a(s_143), .b(gate837inter3), .O(gate837inter10));
  nor2  gate1886(.a(gate837inter10), .b(gate837inter9), .O(gate837inter11));
  nor2  gate1887(.a(gate837inter11), .b(gate837inter6), .O(gate837inter12));
  nand2 gate1888(.a(gate837inter12), .b(gate837inter1), .O(N2843));

  xor2  gate2043(.a(N2828), .b(N2809), .O(gate838inter0));
  nand2 gate2044(.a(gate838inter0), .b(s_166), .O(gate838inter1));
  and2  gate2045(.a(N2828), .b(N2809), .O(gate838inter2));
  inv1  gate2046(.a(s_166), .O(gate838inter3));
  inv1  gate2047(.a(s_167), .O(gate838inter4));
  nand2 gate2048(.a(gate838inter4), .b(gate838inter3), .O(gate838inter5));
  nor2  gate2049(.a(gate838inter5), .b(gate838inter2), .O(gate838inter6));
  inv1  gate2050(.a(N2809), .O(gate838inter7));
  inv1  gate2051(.a(N2828), .O(gate838inter8));
  nand2 gate2052(.a(gate838inter8), .b(gate838inter7), .O(gate838inter9));
  nand2 gate2053(.a(s_167), .b(gate838inter3), .O(gate838inter10));
  nor2  gate2054(.a(gate838inter10), .b(gate838inter9), .O(gate838inter11));
  nor2  gate2055(.a(gate838inter11), .b(gate838inter6), .O(gate838inter12));
  nand2 gate2056(.a(gate838inter12), .b(gate838inter1), .O(N2846));

  xor2  gate2127(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate2128(.a(gate839inter0), .b(s_178), .O(gate839inter1));
  and2  gate2129(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate2130(.a(s_178), .O(gate839inter3));
  inv1  gate2131(.a(s_179), .O(gate839inter4));
  nand2 gate2132(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate2133(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate2134(.a(N2812), .O(gate839inter7));
  inv1  gate2135(.a(N2076), .O(gate839inter8));
  nand2 gate2136(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate2137(.a(s_179), .b(gate839inter3), .O(gate839inter10));
  nor2  gate2138(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate2139(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate2140(.a(gate839inter12), .b(gate839inter1), .O(N2850));
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );

  xor2  gate1791(.a(N1938), .b(N2824), .O(gate843inter0));
  nand2 gate1792(.a(gate843inter0), .b(s_130), .O(gate843inter1));
  and2  gate1793(.a(N1938), .b(N2824), .O(gate843inter2));
  inv1  gate1794(.a(s_130), .O(gate843inter3));
  inv1  gate1795(.a(s_131), .O(gate843inter4));
  nand2 gate1796(.a(gate843inter4), .b(gate843inter3), .O(gate843inter5));
  nor2  gate1797(.a(gate843inter5), .b(gate843inter2), .O(gate843inter6));
  inv1  gate1798(.a(N2824), .O(gate843inter7));
  inv1  gate1799(.a(N1938), .O(gate843inter8));
  nand2 gate1800(.a(gate843inter8), .b(gate843inter7), .O(gate843inter9));
  nand2 gate1801(.a(s_131), .b(gate843inter3), .O(gate843inter10));
  nor2  gate1802(.a(gate843inter10), .b(gate843inter9), .O(gate843inter11));
  nor2  gate1803(.a(gate843inter11), .b(gate843inter6), .O(gate843inter12));
  nand2 gate1804(.a(gate843inter12), .b(gate843inter1), .O(N2854));
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );

  xor2  gate909(.a(N2857), .b(N2052), .O(gate851inter0));
  nand2 gate910(.a(gate851inter0), .b(s_4), .O(gate851inter1));
  and2  gate911(.a(N2857), .b(N2052), .O(gate851inter2));
  inv1  gate912(.a(s_4), .O(gate851inter3));
  inv1  gate913(.a(s_5), .O(gate851inter4));
  nand2 gate914(.a(gate851inter4), .b(gate851inter3), .O(gate851inter5));
  nor2  gate915(.a(gate851inter5), .b(gate851inter2), .O(gate851inter6));
  inv1  gate916(.a(N2052), .O(gate851inter7));
  inv1  gate917(.a(N2857), .O(gate851inter8));
  nand2 gate918(.a(gate851inter8), .b(gate851inter7), .O(gate851inter9));
  nand2 gate919(.a(s_5), .b(gate851inter3), .O(gate851inter10));
  nor2  gate920(.a(gate851inter10), .b(gate851inter9), .O(gate851inter11));
  nor2  gate921(.a(gate851inter11), .b(gate851inter6), .O(gate851inter12));
  nand2 gate922(.a(gate851inter12), .b(gate851inter1), .O(N2866));
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );

  xor2  gate1287(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1288(.a(gate856inter0), .b(s_58), .O(gate856inter1));
  and2  gate1289(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1290(.a(s_58), .O(gate856inter3));
  inv1  gate1291(.a(s_59), .O(gate856inter4));
  nand2 gate1292(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1293(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1294(.a(N2843), .O(gate856inter7));
  inv1  gate1295(.a(N886), .O(gate856inter8));
  nand2 gate1296(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1297(.a(s_59), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1298(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1299(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1300(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );

  xor2  gate1217(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate1218(.a(gate865inter0), .b(s_48), .O(gate865inter1));
  and2  gate1219(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate1220(.a(s_48), .O(gate865inter3));
  inv1  gate1221(.a(s_49), .O(gate865inter4));
  nand2 gate1222(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate1223(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate1224(.a(N2870), .O(gate865inter7));
  inv1  gate1225(.a(N2854), .O(gate865inter8));
  nand2 gate1226(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate1227(.a(s_49), .b(gate865inter3), .O(gate865inter10));
  nor2  gate1228(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate1229(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate1230(.a(gate865inter12), .b(gate865inter1), .O(N2880));
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate2029(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate2030(.a(gate874inter0), .b(s_164), .O(gate874inter1));
  and2  gate2031(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate2032(.a(s_164), .O(gate874inter3));
  inv1  gate2033(.a(s_165), .O(gate874inter4));
  nand2 gate2034(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate2035(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate2036(.a(N2871), .O(gate874inter7));
  inv1  gate2037(.a(N2881), .O(gate874inter8));
  nand2 gate2038(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate2039(.a(s_165), .b(gate874inter3), .O(gate874inter10));
  nor2  gate2040(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate2041(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate2042(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );

  xor2  gate1399(.a(N1461), .b(N2883), .O(gate876inter0));
  nand2 gate1400(.a(gate876inter0), .b(s_74), .O(gate876inter1));
  and2  gate1401(.a(N1461), .b(N2883), .O(gate876inter2));
  inv1  gate1402(.a(s_74), .O(gate876inter3));
  inv1  gate1403(.a(s_75), .O(gate876inter4));
  nand2 gate1404(.a(gate876inter4), .b(gate876inter3), .O(gate876inter5));
  nor2  gate1405(.a(gate876inter5), .b(gate876inter2), .O(gate876inter6));
  inv1  gate1406(.a(N2883), .O(gate876inter7));
  inv1  gate1407(.a(N1461), .O(gate876inter8));
  nand2 gate1408(.a(gate876inter8), .b(gate876inter7), .O(gate876inter9));
  nand2 gate1409(.a(s_75), .b(gate876inter3), .O(gate876inter10));
  nor2  gate1410(.a(gate876inter10), .b(gate876inter9), .O(gate876inter11));
  nor2  gate1411(.a(gate876inter11), .b(gate876inter6), .O(gate876inter12));
  nand2 gate1412(.a(gate876inter12), .b(gate876inter1), .O(N2895));
inv1 gate877( .a(N2883), .O(N2896) );

  xor2  gate1427(.a(N2896), .b(N1383), .O(gate878inter0));
  nand2 gate1428(.a(gate878inter0), .b(s_78), .O(gate878inter1));
  and2  gate1429(.a(N2896), .b(N1383), .O(gate878inter2));
  inv1  gate1430(.a(s_78), .O(gate878inter3));
  inv1  gate1431(.a(s_79), .O(gate878inter4));
  nand2 gate1432(.a(gate878inter4), .b(gate878inter3), .O(gate878inter5));
  nor2  gate1433(.a(gate878inter5), .b(gate878inter2), .O(gate878inter6));
  inv1  gate1434(.a(N1383), .O(gate878inter7));
  inv1  gate1435(.a(N2896), .O(gate878inter8));
  nand2 gate1436(.a(gate878inter8), .b(gate878inter7), .O(gate878inter9));
  nand2 gate1437(.a(s_79), .b(gate878inter3), .O(gate878inter10));
  nor2  gate1438(.a(gate878inter10), .b(gate878inter9), .O(gate878inter11));
  nor2  gate1439(.a(gate878inter11), .b(gate878inter6), .O(gate878inter12));
  nand2 gate1440(.a(gate878inter12), .b(gate878inter1), .O(N2897));
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule