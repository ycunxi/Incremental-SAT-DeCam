module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate623inter0, gate623inter1, gate623inter2, gate623inter3, gate623inter4, gate623inter5, gate623inter6, gate623inter7, gate623inter8, gate623inter9, gate623inter10, gate623inter11, gate623inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate345inter0, gate345inter1, gate345inter2, gate345inter3, gate345inter4, gate345inter5, gate345inter6, gate345inter7, gate345inter8, gate345inter9, gate345inter10, gate345inter11, gate345inter12, gate550inter0, gate550inter1, gate550inter2, gate550inter3, gate550inter4, gate550inter5, gate550inter6, gate550inter7, gate550inter8, gate550inter9, gate550inter10, gate550inter11, gate550inter12, gate669inter0, gate669inter1, gate669inter2, gate669inter3, gate669inter4, gate669inter5, gate669inter6, gate669inter7, gate669inter8, gate669inter9, gate669inter10, gate669inter11, gate669inter12, gate789inter0, gate789inter1, gate789inter2, gate789inter3, gate789inter4, gate789inter5, gate789inter6, gate789inter7, gate789inter8, gate789inter9, gate789inter10, gate789inter11, gate789inter12, gate338inter0, gate338inter1, gate338inter2, gate338inter3, gate338inter4, gate338inter5, gate338inter6, gate338inter7, gate338inter8, gate338inter9, gate338inter10, gate338inter11, gate338inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate600inter0, gate600inter1, gate600inter2, gate600inter3, gate600inter4, gate600inter5, gate600inter6, gate600inter7, gate600inter8, gate600inter9, gate600inter10, gate600inter11, gate600inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate306inter0, gate306inter1, gate306inter2, gate306inter3, gate306inter4, gate306inter5, gate306inter6, gate306inter7, gate306inter8, gate306inter9, gate306inter10, gate306inter11, gate306inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate526inter0, gate526inter1, gate526inter2, gate526inter3, gate526inter4, gate526inter5, gate526inter6, gate526inter7, gate526inter8, gate526inter9, gate526inter10, gate526inter11, gate526inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate523inter0, gate523inter1, gate523inter2, gate523inter3, gate523inter4, gate523inter5, gate523inter6, gate523inter7, gate523inter8, gate523inter9, gate523inter10, gate523inter11, gate523inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate587inter0, gate587inter1, gate587inter2, gate587inter3, gate587inter4, gate587inter5, gate587inter6, gate587inter7, gate587inter8, gate587inter9, gate587inter10, gate587inter11, gate587inter12, gate801inter0, gate801inter1, gate801inter2, gate801inter3, gate801inter4, gate801inter5, gate801inter6, gate801inter7, gate801inter8, gate801inter9, gate801inter10, gate801inter11, gate801inter12, gate637inter0, gate637inter1, gate637inter2, gate637inter3, gate637inter4, gate637inter5, gate637inter6, gate637inter7, gate637inter8, gate637inter9, gate637inter10, gate637inter11, gate637inter12, gate320inter0, gate320inter1, gate320inter2, gate320inter3, gate320inter4, gate320inter5, gate320inter6, gate320inter7, gate320inter8, gate320inter9, gate320inter10, gate320inter11, gate320inter12, gate380inter0, gate380inter1, gate380inter2, gate380inter3, gate380inter4, gate380inter5, gate380inter6, gate380inter7, gate380inter8, gate380inter9, gate380inter10, gate380inter11, gate380inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate329inter0, gate329inter1, gate329inter2, gate329inter3, gate329inter4, gate329inter5, gate329inter6, gate329inter7, gate329inter8, gate329inter9, gate329inter10, gate329inter11, gate329inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate534inter0, gate534inter1, gate534inter2, gate534inter3, gate534inter4, gate534inter5, gate534inter6, gate534inter7, gate534inter8, gate534inter9, gate534inter10, gate534inter11, gate534inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate819inter0, gate819inter1, gate819inter2, gate819inter3, gate819inter4, gate819inter5, gate819inter6, gate819inter7, gate819inter8, gate819inter9, gate819inter10, gate819inter11, gate819inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate540inter0, gate540inter1, gate540inter2, gate540inter3, gate540inter4, gate540inter5, gate540inter6, gate540inter7, gate540inter8, gate540inter9, gate540inter10, gate540inter11, gate540inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate775inter0, gate775inter1, gate775inter2, gate775inter3, gate775inter4, gate775inter5, gate775inter6, gate775inter7, gate775inter8, gate775inter9, gate775inter10, gate775inter11, gate775inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate862inter0, gate862inter1, gate862inter2, gate862inter3, gate862inter4, gate862inter5, gate862inter6, gate862inter7, gate862inter8, gate862inter9, gate862inter10, gate862inter11, gate862inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate353inter0, gate353inter1, gate353inter2, gate353inter3, gate353inter4, gate353inter5, gate353inter6, gate353inter7, gate353inter8, gate353inter9, gate353inter10, gate353inter11, gate353inter12, gate543inter0, gate543inter1, gate543inter2, gate543inter3, gate543inter4, gate543inter5, gate543inter6, gate543inter7, gate543inter8, gate543inter9, gate543inter10, gate543inter11, gate543inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate350inter0, gate350inter1, gate350inter2, gate350inter3, gate350inter4, gate350inter5, gate350inter6, gate350inter7, gate350inter8, gate350inter9, gate350inter10, gate350inter11, gate350inter12, gate867inter0, gate867inter1, gate867inter2, gate867inter3, gate867inter4, gate867inter5, gate867inter6, gate867inter7, gate867inter8, gate867inter9, gate867inter10, gate867inter11, gate867inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12, gate794inter0, gate794inter1, gate794inter2, gate794inter3, gate794inter4, gate794inter5, gate794inter6, gate794inter7, gate794inter8, gate794inter9, gate794inter10, gate794inter11, gate794inter12, gate852inter0, gate852inter1, gate852inter2, gate852inter3, gate852inter4, gate852inter5, gate852inter6, gate852inter7, gate852inter8, gate852inter9, gate852inter10, gate852inter11, gate852inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate864inter0, gate864inter1, gate864inter2, gate864inter3, gate864inter4, gate864inter5, gate864inter6, gate864inter7, gate864inter8, gate864inter9, gate864inter10, gate864inter11, gate864inter12, gate766inter0, gate766inter1, gate766inter2, gate766inter3, gate766inter4, gate766inter5, gate766inter6, gate766inter7, gate766inter8, gate766inter9, gate766inter10, gate766inter11, gate766inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate760inter0, gate760inter1, gate760inter2, gate760inter3, gate760inter4, gate760inter5, gate760inter6, gate760inter7, gate760inter8, gate760inter9, gate760inter10, gate760inter11, gate760inter12, gate516inter0, gate516inter1, gate516inter2, gate516inter3, gate516inter4, gate516inter5, gate516inter6, gate516inter7, gate516inter8, gate516inter9, gate516inter10, gate516inter11, gate516inter12, gate339inter0, gate339inter1, gate339inter2, gate339inter3, gate339inter4, gate339inter5, gate339inter6, gate339inter7, gate339inter8, gate339inter9, gate339inter10, gate339inter11, gate339inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate378inter0, gate378inter1, gate378inter2, gate378inter3, gate378inter4, gate378inter5, gate378inter6, gate378inter7, gate378inter8, gate378inter9, gate378inter10, gate378inter11, gate378inter12, gate802inter0, gate802inter1, gate802inter2, gate802inter3, gate802inter4, gate802inter5, gate802inter6, gate802inter7, gate802inter8, gate802inter9, gate802inter10, gate802inter11, gate802inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate640inter0, gate640inter1, gate640inter2, gate640inter3, gate640inter4, gate640inter5, gate640inter6, gate640inter7, gate640inter8, gate640inter9, gate640inter10, gate640inter11, gate640inter12, gate319inter0, gate319inter1, gate319inter2, gate319inter3, gate319inter4, gate319inter5, gate319inter6, gate319inter7, gate319inter8, gate319inter9, gate319inter10, gate319inter11, gate319inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate583inter0, gate583inter1, gate583inter2, gate583inter3, gate583inter4, gate583inter5, gate583inter6, gate583inter7, gate583inter8, gate583inter9, gate583inter10, gate583inter11, gate583inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12;



inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );

  xor2  gate1161(.a(N91), .b(N66), .O(gate18inter0));
  nand2 gate1162(.a(gate18inter0), .b(s_40), .O(gate18inter1));
  and2  gate1163(.a(N91), .b(N66), .O(gate18inter2));
  inv1  gate1164(.a(s_40), .O(gate18inter3));
  inv1  gate1165(.a(s_41), .O(gate18inter4));
  nand2 gate1166(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1167(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1168(.a(N66), .O(gate18inter7));
  inv1  gate1169(.a(N91), .O(gate18inter8));
  nand2 gate1170(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1171(.a(s_41), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1172(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1173(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1174(.a(gate18inter12), .b(gate18inter1), .O(N252));
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );

  xor2  gate1525(.a(N331), .b(N306), .O(gate76inter0));
  nand2 gate1526(.a(gate76inter0), .b(s_92), .O(gate76inter1));
  and2  gate1527(.a(N331), .b(N306), .O(gate76inter2));
  inv1  gate1528(.a(s_92), .O(gate76inter3));
  inv1  gate1529(.a(s_93), .O(gate76inter4));
  nand2 gate1530(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1531(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1532(.a(N306), .O(gate76inter7));
  inv1  gate1533(.a(N331), .O(gate76inter8));
  nand2 gate1534(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1535(.a(s_93), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1536(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1537(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1538(.a(gate76inter12), .b(gate76inter1), .O(N551));

  xor2  gate1455(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate1456(.a(gate77inter0), .b(s_82), .O(gate77inter1));
  and2  gate1457(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate1458(.a(s_82), .O(gate77inter3));
  inv1  gate1459(.a(s_83), .O(gate77inter4));
  nand2 gate1460(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1461(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1462(.a(N306), .O(gate77inter7));
  inv1  gate1463(.a(N331), .O(gate77inter8));
  nand2 gate1464(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1465(.a(s_83), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1466(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1467(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1468(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate1931(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate1932(.a(gate96inter0), .b(s_150), .O(gate96inter1));
  and2  gate1933(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate1934(.a(s_150), .O(gate96inter3));
  inv1  gate1935(.a(s_151), .O(gate96inter4));
  nand2 gate1936(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1937(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1938(.a(N326), .O(gate96inter7));
  inv1  gate1939(.a(N277), .O(gate96inter8));
  nand2 gate1940(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1941(.a(s_151), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1942(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1943(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1944(.a(gate96inter12), .b(gate96inter1), .O(N601));
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );

  xor2  gate1245(.a(N608), .b(N56), .O(gate163inter0));
  nand2 gate1246(.a(gate163inter0), .b(s_52), .O(gate163inter1));
  and2  gate1247(.a(N608), .b(N56), .O(gate163inter2));
  inv1  gate1248(.a(s_52), .O(gate163inter3));
  inv1  gate1249(.a(s_53), .O(gate163inter4));
  nand2 gate1250(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1251(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1252(.a(N56), .O(gate163inter7));
  inv1  gate1253(.a(N608), .O(gate163inter8));
  nand2 gate1254(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1255(.a(s_53), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1256(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1257(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1258(.a(gate163inter12), .b(gate163inter1), .O(N910));
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );

  xor2  gate1539(.a(N890), .b(N625), .O(gate235inter0));
  nand2 gate1540(.a(gate235inter0), .b(s_94), .O(gate235inter1));
  and2  gate1541(.a(N890), .b(N625), .O(gate235inter2));
  inv1  gate1542(.a(s_94), .O(gate235inter3));
  inv1  gate1543(.a(s_95), .O(gate235inter4));
  nand2 gate1544(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1545(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1546(.a(N625), .O(gate235inter7));
  inv1  gate1547(.a(N890), .O(gate235inter8));
  nand2 gate1548(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1549(.a(s_95), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1550(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1551(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1552(.a(gate235inter12), .b(gate235inter1), .O(N1063));
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );

  xor2  gate1091(.a(N988), .b(N721), .O(gate239inter0));
  nand2 gate1092(.a(gate239inter0), .b(s_30), .O(gate239inter1));
  and2  gate1093(.a(N988), .b(N721), .O(gate239inter2));
  inv1  gate1094(.a(s_30), .O(gate239inter3));
  inv1  gate1095(.a(s_31), .O(gate239inter4));
  nand2 gate1096(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1097(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1098(.a(N721), .O(gate239inter7));
  inv1  gate1099(.a(N988), .O(gate239inter8));
  nand2 gate1100(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1101(.a(s_31), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1102(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1103(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1104(.a(gate239inter12), .b(gate239inter1), .O(N1119));

  xor2  gate2197(.a(N989), .b(N718), .O(gate240inter0));
  nand2 gate2198(.a(gate240inter0), .b(s_188), .O(gate240inter1));
  and2  gate2199(.a(N989), .b(N718), .O(gate240inter2));
  inv1  gate2200(.a(s_188), .O(gate240inter3));
  inv1  gate2201(.a(s_189), .O(gate240inter4));
  nand2 gate2202(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2203(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2204(.a(N718), .O(gate240inter7));
  inv1  gate2205(.a(N989), .O(gate240inter8));
  nand2 gate2206(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2207(.a(s_189), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2208(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2209(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2210(.a(gate240inter12), .b(gate240inter1), .O(N1120));
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );

  xor2  gate881(.a(N1009), .b(N748), .O(gate248inter0));
  nand2 gate882(.a(gate248inter0), .b(s_0), .O(gate248inter1));
  and2  gate883(.a(N1009), .b(N748), .O(gate248inter2));
  inv1  gate884(.a(s_0), .O(gate248inter3));
  inv1  gate885(.a(s_1), .O(gate248inter4));
  nand2 gate886(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate887(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate888(.a(N748), .O(gate248inter7));
  inv1  gate889(.a(N1009), .O(gate248inter8));
  nand2 gate890(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate891(.a(s_1), .b(gate248inter3), .O(gate248inter10));
  nor2  gate892(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate893(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate894(.a(gate248inter12), .b(gate248inter1), .O(N1133));
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate1231(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate1232(.a(gate268inter0), .b(s_50), .O(gate268inter1));
  and2  gate1233(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate1234(.a(s_50), .O(gate268inter3));
  inv1  gate1235(.a(s_51), .O(gate268inter4));
  nand2 gate1236(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1237(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1238(.a(N921), .O(gate268inter7));
  inv1  gate1239(.a(N923), .O(gate268inter8));
  nand2 gate1240(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1241(.a(s_51), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1242(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1243(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1244(.a(gate268inter12), .b(gate268inter1), .O(N1171));
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate1063(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate1064(.a(gate275inter0), .b(s_26), .O(gate275inter1));
  and2  gate1065(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate1066(.a(s_26), .O(gate275inter3));
  inv1  gate1067(.a(s_27), .O(gate275inter4));
  nand2 gate1068(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1069(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1070(.a(N1016), .O(gate275inter7));
  inv1  gate1071(.a(N946), .O(gate275inter8));
  nand2 gate1072(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1073(.a(s_27), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1074(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1075(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1076(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );

  xor2  gate2155(.a(N958), .b(N1025), .O(gate281inter0));
  nand2 gate2156(.a(gate281inter0), .b(s_182), .O(gate281inter1));
  and2  gate2157(.a(N958), .b(N1025), .O(gate281inter2));
  inv1  gate2158(.a(s_182), .O(gate281inter3));
  inv1  gate2159(.a(s_183), .O(gate281inter4));
  nand2 gate2160(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2161(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2162(.a(N1025), .O(gate281inter7));
  inv1  gate2163(.a(N958), .O(gate281inter8));
  nand2 gate2164(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2165(.a(s_183), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2166(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2167(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2168(.a(gate281inter12), .b(gate281inter1), .O(N1216));
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );

  xor2  gate1805(.a(N984), .b(N981), .O(gate296inter0));
  nand2 gate1806(.a(gate296inter0), .b(s_132), .O(gate296inter1));
  and2  gate1807(.a(N984), .b(N981), .O(gate296inter2));
  inv1  gate1808(.a(s_132), .O(gate296inter3));
  inv1  gate1809(.a(s_133), .O(gate296inter4));
  nand2 gate1810(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1811(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1812(.a(N981), .O(gate296inter7));
  inv1  gate1813(.a(N984), .O(gate296inter8));
  nand2 gate1814(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1815(.a(s_133), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1816(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1817(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1818(.a(gate296inter12), .b(gate296inter1), .O(N1231));
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );

  xor2  gate1105(.a(N1133), .b(N1132), .O(gate306inter0));
  nand2 gate1106(.a(gate306inter0), .b(s_32), .O(gate306inter1));
  and2  gate1107(.a(N1133), .b(N1132), .O(gate306inter2));
  inv1  gate1108(.a(s_32), .O(gate306inter3));
  inv1  gate1109(.a(s_33), .O(gate306inter4));
  nand2 gate1110(.a(gate306inter4), .b(gate306inter3), .O(gate306inter5));
  nor2  gate1111(.a(gate306inter5), .b(gate306inter2), .O(gate306inter6));
  inv1  gate1112(.a(N1132), .O(gate306inter7));
  inv1  gate1113(.a(N1133), .O(gate306inter8));
  nand2 gate1114(.a(gate306inter8), .b(gate306inter7), .O(gate306inter9));
  nand2 gate1115(.a(s_33), .b(gate306inter3), .O(gate306inter10));
  nor2  gate1116(.a(gate306inter10), .b(gate306inter9), .O(gate306inter11));
  nor2  gate1117(.a(gate306inter11), .b(gate306inter6), .O(gate306inter12));
  nand2 gate1118(.a(gate306inter12), .b(gate306inter1), .O(N1249));
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );

  xor2  gate2085(.a(N1205), .b(N688), .O(gate313inter0));
  nand2 gate2086(.a(gate313inter0), .b(s_172), .O(gate313inter1));
  and2  gate2087(.a(N1205), .b(N688), .O(gate313inter2));
  inv1  gate2088(.a(s_172), .O(gate313inter3));
  inv1  gate2089(.a(s_173), .O(gate313inter4));
  nand2 gate2090(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate2091(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate2092(.a(N688), .O(gate313inter7));
  inv1  gate2093(.a(N1205), .O(gate313inter8));
  nand2 gate2094(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate2095(.a(s_173), .b(gate313inter3), .O(gate313inter10));
  nor2  gate2096(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate2097(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate2098(.a(gate313inter12), .b(gate313inter1), .O(N1309));
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );

  xor2  gate1833(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate1834(.a(gate316inter0), .b(s_136), .O(gate316inter1));
  and2  gate1835(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate1836(.a(s_136), .O(gate316inter3));
  inv1  gate1837(.a(s_137), .O(gate316inter4));
  nand2 gate1838(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate1839(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate1840(.a(N697), .O(gate316inter7));
  inv1  gate1841(.a(N1211), .O(gate316inter8));
  nand2 gate1842(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate1843(.a(s_137), .b(gate316inter3), .O(gate316inter10));
  nor2  gate1844(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate1845(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate1846(.a(gate316inter12), .b(gate316inter1), .O(N1312));

  xor2  gate1889(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate1890(.a(gate317inter0), .b(s_144), .O(gate317inter1));
  and2  gate1891(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate1892(.a(s_144), .O(gate317inter3));
  inv1  gate1893(.a(s_145), .O(gate317inter4));
  nand2 gate1894(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate1895(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate1896(.a(N700), .O(gate317inter7));
  inv1  gate1897(.a(N1213), .O(gate317inter8));
  nand2 gate1898(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate1899(.a(s_145), .b(gate317inter3), .O(gate317inter10));
  nor2  gate1900(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate1901(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate1902(.a(gate317inter12), .b(gate317inter1), .O(N1313));
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );

  xor2  gate2225(.a(N1220), .b(N706), .O(gate319inter0));
  nand2 gate2226(.a(gate319inter0), .b(s_192), .O(gate319inter1));
  and2  gate2227(.a(N1220), .b(N706), .O(gate319inter2));
  inv1  gate2228(.a(s_192), .O(gate319inter3));
  inv1  gate2229(.a(s_193), .O(gate319inter4));
  nand2 gate2230(.a(gate319inter4), .b(gate319inter3), .O(gate319inter5));
  nor2  gate2231(.a(gate319inter5), .b(gate319inter2), .O(gate319inter6));
  inv1  gate2232(.a(N706), .O(gate319inter7));
  inv1  gate2233(.a(N1220), .O(gate319inter8));
  nand2 gate2234(.a(gate319inter8), .b(gate319inter7), .O(gate319inter9));
  nand2 gate2235(.a(s_193), .b(gate319inter3), .O(gate319inter10));
  nor2  gate2236(.a(gate319inter10), .b(gate319inter9), .O(gate319inter11));
  nor2  gate2237(.a(gate319inter11), .b(gate319inter6), .O(gate319inter12));
  nand2 gate2238(.a(gate319inter12), .b(gate319inter1), .O(N1315));

  xor2  gate1329(.a(N1223), .b(N709), .O(gate320inter0));
  nand2 gate1330(.a(gate320inter0), .b(s_64), .O(gate320inter1));
  and2  gate1331(.a(N1223), .b(N709), .O(gate320inter2));
  inv1  gate1332(.a(s_64), .O(gate320inter3));
  inv1  gate1333(.a(s_65), .O(gate320inter4));
  nand2 gate1334(.a(gate320inter4), .b(gate320inter3), .O(gate320inter5));
  nor2  gate1335(.a(gate320inter5), .b(gate320inter2), .O(gate320inter6));
  inv1  gate1336(.a(N709), .O(gate320inter7));
  inv1  gate1337(.a(N1223), .O(gate320inter8));
  nand2 gate1338(.a(gate320inter8), .b(gate320inter7), .O(gate320inter9));
  nand2 gate1339(.a(s_65), .b(gate320inter3), .O(gate320inter10));
  nor2  gate1340(.a(gate320inter10), .b(gate320inter9), .O(gate320inter11));
  nor2  gate1341(.a(gate320inter11), .b(gate320inter6), .O(gate320inter12));
  nand2 gate1342(.a(gate320inter12), .b(gate320inter1), .O(N1316));
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );

  xor2  gate2029(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate2030(.a(gate326inter0), .b(s_164), .O(gate326inter1));
  and2  gate2031(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate2032(.a(s_164), .O(gate326inter3));
  inv1  gate2033(.a(s_165), .O(gate326inter4));
  nand2 gate2034(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate2035(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate2036(.a(N733), .O(gate326inter7));
  inv1  gate2037(.a(N1241), .O(gate326inter8));
  nand2 gate2038(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate2039(.a(s_165), .b(gate326inter3), .O(gate326inter10));
  nor2  gate2040(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate2041(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate2042(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );

  xor2  gate1609(.a(N1160), .b(N1267), .O(gate328inter0));
  nand2 gate1610(.a(gate328inter0), .b(s_104), .O(gate328inter1));
  and2  gate1611(.a(N1160), .b(N1267), .O(gate328inter2));
  inv1  gate1612(.a(s_104), .O(gate328inter3));
  inv1  gate1613(.a(s_105), .O(gate328inter4));
  nand2 gate1614(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate1615(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate1616(.a(N1267), .O(gate328inter7));
  inv1  gate1617(.a(N1160), .O(gate328inter8));
  nand2 gate1618(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate1619(.a(s_105), .b(gate328inter3), .O(gate328inter10));
  nor2  gate1620(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate1621(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate1622(.a(gate328inter12), .b(gate328inter1), .O(N1344));

  xor2  gate1371(.a(N894), .b(N1249), .O(gate329inter0));
  nand2 gate1372(.a(gate329inter0), .b(s_70), .O(gate329inter1));
  and2  gate1373(.a(N894), .b(N1249), .O(gate329inter2));
  inv1  gate1374(.a(s_70), .O(gate329inter3));
  inv1  gate1375(.a(s_71), .O(gate329inter4));
  nand2 gate1376(.a(gate329inter4), .b(gate329inter3), .O(gate329inter5));
  nor2  gate1377(.a(gate329inter5), .b(gate329inter2), .O(gate329inter6));
  inv1  gate1378(.a(N1249), .O(gate329inter7));
  inv1  gate1379(.a(N894), .O(gate329inter8));
  nand2 gate1380(.a(gate329inter8), .b(gate329inter7), .O(gate329inter9));
  nand2 gate1381(.a(s_71), .b(gate329inter3), .O(gate329inter10));
  nor2  gate1382(.a(gate329inter10), .b(gate329inter9), .O(gate329inter11));
  nor2  gate1383(.a(gate329inter11), .b(gate329inter6), .O(gate329inter12));
  nand2 gate1384(.a(gate329inter12), .b(gate329inter1), .O(N1345));
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );

  xor2  gate2043(.a(N1210), .b(N1311), .O(gate337inter0));
  nand2 gate2044(.a(gate337inter0), .b(s_166), .O(gate337inter1));
  and2  gate2045(.a(N1210), .b(N1311), .O(gate337inter2));
  inv1  gate2046(.a(s_166), .O(gate337inter3));
  inv1  gate2047(.a(s_167), .O(gate337inter4));
  nand2 gate2048(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate2049(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate2050(.a(N1311), .O(gate337inter7));
  inv1  gate2051(.a(N1210), .O(gate337inter8));
  nand2 gate2052(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate2053(.a(s_167), .b(gate337inter3), .O(gate337inter10));
  nor2  gate2054(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate2055(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate2056(.a(gate337inter12), .b(gate337inter1), .O(N1358));

  xor2  gate1007(.a(N1212), .b(N1312), .O(gate338inter0));
  nand2 gate1008(.a(gate338inter0), .b(s_18), .O(gate338inter1));
  and2  gate1009(.a(N1212), .b(N1312), .O(gate338inter2));
  inv1  gate1010(.a(s_18), .O(gate338inter3));
  inv1  gate1011(.a(s_19), .O(gate338inter4));
  nand2 gate1012(.a(gate338inter4), .b(gate338inter3), .O(gate338inter5));
  nor2  gate1013(.a(gate338inter5), .b(gate338inter2), .O(gate338inter6));
  inv1  gate1014(.a(N1312), .O(gate338inter7));
  inv1  gate1015(.a(N1212), .O(gate338inter8));
  nand2 gate1016(.a(gate338inter8), .b(gate338inter7), .O(gate338inter9));
  nand2 gate1017(.a(s_19), .b(gate338inter3), .O(gate338inter10));
  nor2  gate1018(.a(gate338inter10), .b(gate338inter9), .O(gate338inter11));
  nor2  gate1019(.a(gate338inter11), .b(gate338inter6), .O(gate338inter12));
  nand2 gate1020(.a(gate338inter12), .b(gate338inter1), .O(N1361));

  xor2  gate2141(.a(N1214), .b(N1313), .O(gate339inter0));
  nand2 gate2142(.a(gate339inter0), .b(s_180), .O(gate339inter1));
  and2  gate2143(.a(N1214), .b(N1313), .O(gate339inter2));
  inv1  gate2144(.a(s_180), .O(gate339inter3));
  inv1  gate2145(.a(s_181), .O(gate339inter4));
  nand2 gate2146(.a(gate339inter4), .b(gate339inter3), .O(gate339inter5));
  nor2  gate2147(.a(gate339inter5), .b(gate339inter2), .O(gate339inter6));
  inv1  gate2148(.a(N1313), .O(gate339inter7));
  inv1  gate2149(.a(N1214), .O(gate339inter8));
  nand2 gate2150(.a(gate339inter8), .b(gate339inter7), .O(gate339inter9));
  nand2 gate2151(.a(s_181), .b(gate339inter3), .O(gate339inter10));
  nor2  gate2152(.a(gate339inter10), .b(gate339inter9), .O(gate339inter11));
  nor2  gate2153(.a(gate339inter11), .b(gate339inter6), .O(gate339inter12));
  nand2 gate2154(.a(gate339inter12), .b(gate339inter1), .O(N1364));
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );

  xor2  gate951(.a(N1231), .b(N1322), .O(gate345inter0));
  nand2 gate952(.a(gate345inter0), .b(s_10), .O(gate345inter1));
  and2  gate953(.a(N1231), .b(N1322), .O(gate345inter2));
  inv1  gate954(.a(s_10), .O(gate345inter3));
  inv1  gate955(.a(s_11), .O(gate345inter4));
  nand2 gate956(.a(gate345inter4), .b(gate345inter3), .O(gate345inter5));
  nor2  gate957(.a(gate345inter5), .b(gate345inter2), .O(gate345inter6));
  inv1  gate958(.a(N1322), .O(gate345inter7));
  inv1  gate959(.a(N1231), .O(gate345inter8));
  nand2 gate960(.a(gate345inter8), .b(gate345inter7), .O(gate345inter9));
  nand2 gate961(.a(s_11), .b(gate345inter3), .O(gate345inter10));
  nor2  gate962(.a(gate345inter10), .b(gate345inter9), .O(gate345inter11));
  nor2  gate963(.a(gate345inter11), .b(gate345inter6), .O(gate345inter12));
  nand2 gate964(.a(gate345inter12), .b(gate345inter1), .O(N1383));
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate1273(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate1274(.a(gate347inter0), .b(s_56), .O(gate347inter1));
  and2  gate1275(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate1276(.a(s_56), .O(gate347inter3));
  inv1  gate1277(.a(s_57), .O(gate347inter4));
  nand2 gate1278(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate1279(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate1280(.a(N1232), .O(gate347inter7));
  inv1  gate1281(.a(N990), .O(gate347inter8));
  nand2 gate1282(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate1283(.a(s_57), .b(gate347inter3), .O(gate347inter10));
  nor2  gate1284(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate1285(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate1286(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );

  xor2  gate1959(.a(N1239), .b(N1327), .O(gate350inter0));
  nand2 gate1960(.a(gate350inter0), .b(s_154), .O(gate350inter1));
  and2  gate1961(.a(N1239), .b(N1327), .O(gate350inter2));
  inv1  gate1962(.a(s_154), .O(gate350inter3));
  inv1  gate1963(.a(s_155), .O(gate350inter4));
  nand2 gate1964(.a(gate350inter4), .b(gate350inter3), .O(gate350inter5));
  nor2  gate1965(.a(gate350inter5), .b(gate350inter2), .O(gate350inter6));
  inv1  gate1966(.a(N1327), .O(gate350inter7));
  inv1  gate1967(.a(N1239), .O(gate350inter8));
  nand2 gate1968(.a(gate350inter8), .b(gate350inter7), .O(gate350inter9));
  nand2 gate1969(.a(s_155), .b(gate350inter3), .O(gate350inter10));
  nor2  gate1970(.a(gate350inter10), .b(gate350inter9), .O(gate350inter11));
  nor2  gate1971(.a(gate350inter11), .b(gate350inter6), .O(gate350inter12));
  nand2 gate1972(.a(gate350inter12), .b(gate350inter1), .O(N1390));
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );

  xor2  gate1903(.a(N1004), .b(N1243), .O(gate353inter0));
  nand2 gate1904(.a(gate353inter0), .b(s_146), .O(gate353inter1));
  and2  gate1905(.a(N1004), .b(N1243), .O(gate353inter2));
  inv1  gate1906(.a(s_146), .O(gate353inter3));
  inv1  gate1907(.a(s_147), .O(gate353inter4));
  nand2 gate1908(.a(gate353inter4), .b(gate353inter3), .O(gate353inter5));
  nor2  gate1909(.a(gate353inter5), .b(gate353inter2), .O(gate353inter6));
  inv1  gate1910(.a(N1243), .O(gate353inter7));
  inv1  gate1911(.a(N1004), .O(gate353inter8));
  nand2 gate1912(.a(gate353inter8), .b(gate353inter7), .O(gate353inter9));
  nand2 gate1913(.a(s_147), .b(gate353inter3), .O(gate353inter10));
  nor2  gate1914(.a(gate353inter10), .b(gate353inter9), .O(gate353inter11));
  nor2  gate1915(.a(gate353inter11), .b(gate353inter6), .O(gate353inter12));
  nand2 gate1916(.a(gate353inter12), .b(gate353inter1), .O(N1397));
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate1357(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate1358(.a(gate376inter0), .b(s_68), .O(gate376inter1));
  and2  gate1359(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate1360(.a(s_68), .O(gate376inter3));
  inv1  gate1361(.a(s_69), .O(gate376inter4));
  nand2 gate1362(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate1363(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate1364(.a(N1364), .O(gate376inter7));
  inv1  gate1365(.a(N1154), .O(gate376inter8));
  nand2 gate1366(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate1367(.a(s_69), .b(gate376inter3), .O(gate376inter10));
  nor2  gate1368(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate1369(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate1370(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );

  xor2  gate2169(.a(N1156), .b(N1373), .O(gate378inter0));
  nand2 gate2170(.a(gate378inter0), .b(s_184), .O(gate378inter1));
  and2  gate2171(.a(N1156), .b(N1373), .O(gate378inter2));
  inv1  gate2172(.a(s_184), .O(gate378inter3));
  inv1  gate2173(.a(s_185), .O(gate378inter4));
  nand2 gate2174(.a(gate378inter4), .b(gate378inter3), .O(gate378inter5));
  nor2  gate2175(.a(gate378inter5), .b(gate378inter2), .O(gate378inter6));
  inv1  gate2176(.a(N1373), .O(gate378inter7));
  inv1  gate2177(.a(N1156), .O(gate378inter8));
  nand2 gate2178(.a(gate378inter8), .b(gate378inter7), .O(gate378inter9));
  nand2 gate2179(.a(s_185), .b(gate378inter3), .O(gate378inter10));
  nor2  gate2180(.a(gate378inter10), .b(gate378inter9), .O(gate378inter11));
  nor2  gate2181(.a(gate378inter11), .b(gate378inter6), .O(gate378inter12));
  nand2 gate2182(.a(gate378inter12), .b(gate378inter1), .O(N1457));
inv1 gate379( .a(N1373), .O(N1458) );

  xor2  gate1343(.a(N1157), .b(N1379), .O(gate380inter0));
  nand2 gate1344(.a(gate380inter0), .b(s_66), .O(gate380inter1));
  and2  gate1345(.a(N1157), .b(N1379), .O(gate380inter2));
  inv1  gate1346(.a(s_66), .O(gate380inter3));
  inv1  gate1347(.a(s_67), .O(gate380inter4));
  nand2 gate1348(.a(gate380inter4), .b(gate380inter3), .O(gate380inter5));
  nor2  gate1349(.a(gate380inter5), .b(gate380inter2), .O(gate380inter6));
  inv1  gate1350(.a(N1379), .O(gate380inter7));
  inv1  gate1351(.a(N1157), .O(gate380inter8));
  nand2 gate1352(.a(gate380inter8), .b(gate380inter7), .O(gate380inter9));
  nand2 gate1353(.a(s_67), .b(gate380inter3), .O(gate380inter10));
  nor2  gate1354(.a(gate380inter10), .b(gate380inter9), .O(gate380inter11));
  nor2  gate1355(.a(gate380inter11), .b(gate380inter6), .O(gate380inter12));
  nand2 gate1356(.a(gate380inter12), .b(gate380inter1), .O(N1459));
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate1567(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate1568(.a(gate383inter0), .b(s_98), .O(gate383inter1));
  and2  gate1569(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate1570(.a(s_98), .O(gate383inter3));
  inv1  gate1571(.a(s_99), .O(gate383inter4));
  nand2 gate1572(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate1573(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate1574(.a(N1393), .O(gate383inter7));
  inv1  gate1575(.a(N1161), .O(gate383inter8));
  nand2 gate1576(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate1577(.a(s_99), .b(gate383inter3), .O(gate383inter10));
  nor2  gate1578(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate1579(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate1580(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );

  xor2  gate1385(.a(N1222), .b(N1370), .O(gate387inter0));
  nand2 gate1386(.a(gate387inter0), .b(s_72), .O(gate387inter1));
  and2  gate1387(.a(N1222), .b(N1370), .O(gate387inter2));
  inv1  gate1388(.a(s_72), .O(gate387inter3));
  inv1  gate1389(.a(s_73), .O(gate387inter4));
  nand2 gate1390(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1391(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1392(.a(N1370), .O(gate387inter7));
  inv1  gate1393(.a(N1222), .O(gate387inter8));
  nand2 gate1394(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1395(.a(s_73), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1396(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1397(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1398(.a(gate387inter12), .b(gate387inter1), .O(N1469));
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );

  xor2  gate2253(.a(N1433), .b(N1387), .O(gate390inter0));
  nand2 gate2254(.a(gate390inter0), .b(s_196), .O(gate390inter1));
  and2  gate2255(.a(N1433), .b(N1387), .O(gate390inter2));
  inv1  gate2256(.a(s_196), .O(gate390inter3));
  inv1  gate2257(.a(s_197), .O(gate390inter4));
  nand2 gate2258(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2259(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2260(.a(N1387), .O(gate390inter7));
  inv1  gate2261(.a(N1433), .O(gate390inter8));
  nand2 gate2262(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2263(.a(s_197), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2264(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2265(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2266(.a(gate390inter12), .b(gate390inter1), .O(N1472));
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );

  xor2  gate1651(.a(N1434), .b(N1389), .O(gate393inter0));
  nand2 gate1652(.a(gate393inter0), .b(s_110), .O(gate393inter1));
  and2  gate1653(.a(N1434), .b(N1389), .O(gate393inter2));
  inv1  gate1654(.a(s_110), .O(gate393inter3));
  inv1  gate1655(.a(s_111), .O(gate393inter4));
  nand2 gate1656(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1657(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1658(.a(N1389), .O(gate393inter7));
  inv1  gate1659(.a(N1434), .O(gate393inter8));
  nand2 gate1660(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1661(.a(s_111), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1662(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1663(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1664(.a(gate393inter12), .b(gate393inter1), .O(N1478));
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );

  xor2  gate1021(.a(N1438), .b(N1397), .O(gate395inter0));
  nand2 gate1022(.a(gate395inter0), .b(s_20), .O(gate395inter1));
  and2  gate1023(.a(N1438), .b(N1397), .O(gate395inter2));
  inv1  gate1024(.a(s_20), .O(gate395inter3));
  inv1  gate1025(.a(s_21), .O(gate395inter4));
  nand2 gate1026(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1027(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1028(.a(N1397), .O(gate395inter7));
  inv1  gate1029(.a(N1438), .O(gate395inter8));
  nand2 gate1030(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1031(.a(s_21), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1032(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1033(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1034(.a(gate395inter12), .b(gate395inter1), .O(N1484));
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );

  xor2  gate1595(.a(N1448), .b(N943), .O(gate398inter0));
  nand2 gate1596(.a(gate398inter0), .b(s_102), .O(gate398inter1));
  and2  gate1597(.a(N1448), .b(N943), .O(gate398inter2));
  inv1  gate1598(.a(s_102), .O(gate398inter3));
  inv1  gate1599(.a(s_103), .O(gate398inter4));
  nand2 gate1600(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1601(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1602(.a(N943), .O(gate398inter7));
  inv1  gate1603(.a(N1448), .O(gate398inter8));
  nand2 gate1604(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1605(.a(s_103), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1606(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1607(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1608(.a(gate398inter12), .b(gate398inter1), .O(N1489));
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );

  xor2  gate1469(.a(N1460), .b(N977), .O(gate405inter0));
  nand2 gate1470(.a(gate405inter0), .b(s_84), .O(gate405inter1));
  and2  gate1471(.a(N1460), .b(N977), .O(gate405inter2));
  inv1  gate1472(.a(s_84), .O(gate405inter3));
  inv1  gate1473(.a(s_85), .O(gate405inter4));
  nand2 gate1474(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1475(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1476(.a(N977), .O(gate405inter7));
  inv1  gate1477(.a(N1460), .O(gate405inter8));
  nand2 gate1478(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1479(.a(s_85), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1480(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1481(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1482(.a(gate405inter12), .b(gate405inter1), .O(N1496));

  xor2  gate1945(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate1946(.a(gate406inter0), .b(s_152), .O(gate406inter1));
  and2  gate1947(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate1948(.a(s_152), .O(gate406inter3));
  inv1  gate1949(.a(s_153), .O(gate406inter4));
  nand2 gate1950(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1951(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1952(.a(N998), .O(gate406inter7));
  inv1  gate1953(.a(N1463), .O(gate406inter8));
  nand2 gate1954(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1955(.a(s_153), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1956(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1957(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1958(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );

  xor2  gate1189(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate1190(.a(gate410inter0), .b(s_44), .O(gate410inter1));
  and2  gate1191(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate1192(.a(s_44), .O(gate410inter3));
  inv1  gate1193(.a(s_45), .O(gate410inter4));
  nand2 gate1194(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1195(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1196(.a(N994), .O(gate410inter7));
  inv1  gate1197(.a(N1475), .O(gate410inter8));
  nand2 gate1198(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1199(.a(s_45), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1200(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1201(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1202(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );

  xor2  gate1791(.a(N1487), .b(N1443), .O(gate412inter0));
  nand2 gate1792(.a(gate412inter0), .b(s_130), .O(gate412inter1));
  and2  gate1793(.a(N1487), .b(N1443), .O(gate412inter2));
  inv1  gate1794(.a(s_130), .O(gate412inter3));
  inv1  gate1795(.a(s_131), .O(gate412inter4));
  nand2 gate1796(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1797(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1798(.a(N1443), .O(gate412inter7));
  inv1  gate1799(.a(N1487), .O(gate412inter8));
  nand2 gate1800(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1801(.a(s_131), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1802(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1803(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1804(.a(gate412inter12), .b(gate412inter1), .O(N1513));
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );

  xor2  gate1735(.a(N1530), .b(N1540), .O(gate440inter0));
  nand2 gate1736(.a(gate440inter0), .b(s_122), .O(gate440inter1));
  and2  gate1737(.a(N1530), .b(N1540), .O(gate440inter2));
  inv1  gate1738(.a(s_122), .O(gate440inter3));
  inv1  gate1739(.a(s_123), .O(gate440inter4));
  nand2 gate1740(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1741(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1742(.a(N1540), .O(gate440inter7));
  inv1  gate1743(.a(N1530), .O(gate440inter8));
  nand2 gate1744(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1745(.a(s_123), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1746(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1747(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1748(.a(gate440inter12), .b(gate440inter1), .O(N1594));
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );

  xor2  gate1511(.a(N1217), .b(N1606), .O(gate466inter0));
  nand2 gate1512(.a(gate466inter0), .b(s_90), .O(gate466inter1));
  and2  gate1513(.a(N1217), .b(N1606), .O(gate466inter2));
  inv1  gate1514(.a(s_90), .O(gate466inter3));
  inv1  gate1515(.a(s_91), .O(gate466inter4));
  nand2 gate1516(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1517(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1518(.a(N1606), .O(gate466inter7));
  inv1  gate1519(.a(N1217), .O(gate466inter8));
  nand2 gate1520(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1521(.a(s_91), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1522(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1523(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1524(.a(gate466inter12), .b(gate466inter1), .O(N1678));
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );

  xor2  gate1133(.a(N1639), .b(N1510), .O(gate473inter0));
  nand2 gate1134(.a(gate473inter0), .b(s_36), .O(gate473inter1));
  and2  gate1135(.a(N1639), .b(N1510), .O(gate473inter2));
  inv1  gate1136(.a(s_36), .O(gate473inter3));
  inv1  gate1137(.a(s_37), .O(gate473inter4));
  nand2 gate1138(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1139(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1140(.a(N1510), .O(gate473inter7));
  inv1  gate1141(.a(N1639), .O(gate473inter8));
  nand2 gate1142(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1143(.a(s_37), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1144(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1145(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1146(.a(gate473inter12), .b(gate473inter1), .O(N1688));
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );

  xor2  gate1203(.a(N1672), .b(N643), .O(gate476inter0));
  nand2 gate1204(.a(gate476inter0), .b(s_46), .O(gate476inter1));
  and2  gate1205(.a(N1672), .b(N643), .O(gate476inter2));
  inv1  gate1206(.a(s_46), .O(gate476inter3));
  inv1  gate1207(.a(s_47), .O(gate476inter4));
  nand2 gate1208(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1209(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1210(.a(N643), .O(gate476inter7));
  inv1  gate1211(.a(N1672), .O(gate476inter8));
  nand2 gate1212(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1213(.a(s_47), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1214(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1215(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1216(.a(gate476inter12), .b(gate476inter1), .O(N1706));
inv1 gate477( .a(N1643), .O(N1707) );

  xor2  gate1819(.a(N1675), .b(N1647), .O(gate478inter0));
  nand2 gate1820(.a(gate478inter0), .b(s_134), .O(gate478inter1));
  and2  gate1821(.a(N1675), .b(N1647), .O(gate478inter2));
  inv1  gate1822(.a(s_134), .O(gate478inter3));
  inv1  gate1823(.a(s_135), .O(gate478inter4));
  nand2 gate1824(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1825(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1826(.a(N1647), .O(gate478inter7));
  inv1  gate1827(.a(N1675), .O(gate478inter8));
  nand2 gate1828(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1829(.a(s_135), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1830(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1831(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1832(.a(gate478inter12), .b(gate478inter1), .O(N1708));
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );

  xor2  gate1707(.a(N1688), .b(N1638), .O(gate488inter0));
  nand2 gate1708(.a(gate488inter0), .b(s_118), .O(gate488inter1));
  and2  gate1709(.a(N1688), .b(N1638), .O(gate488inter2));
  inv1  gate1710(.a(s_118), .O(gate488inter3));
  inv1  gate1711(.a(s_119), .O(gate488inter4));
  nand2 gate1712(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1713(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1714(.a(N1638), .O(gate488inter7));
  inv1  gate1715(.a(N1688), .O(gate488inter8));
  nand2 gate1716(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1717(.a(s_119), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1718(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1719(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1720(.a(gate488inter12), .b(gate488inter1), .O(N1723));
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );

  xor2  gate1875(.a(N1709), .b(N1600), .O(gate497inter0));
  nand2 gate1876(.a(gate497inter0), .b(s_142), .O(gate497inter1));
  and2  gate1877(.a(N1709), .b(N1600), .O(gate497inter2));
  inv1  gate1878(.a(s_142), .O(gate497inter3));
  inv1  gate1879(.a(s_143), .O(gate497inter4));
  nand2 gate1880(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1881(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1882(.a(N1600), .O(gate497inter7));
  inv1  gate1883(.a(N1709), .O(gate497inter8));
  nand2 gate1884(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1885(.a(s_143), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1886(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1887(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1888(.a(gate497inter12), .b(gate497inter1), .O(N1746));
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );

  xor2  gate909(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate910(.a(gate499inter0), .b(s_4), .O(gate499inter1));
  and2  gate911(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate912(.a(s_4), .O(gate499inter3));
  inv1  gate913(.a(s_5), .O(gate499inter4));
  nand2 gate914(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate915(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate916(.a(N1678), .O(gate499inter7));
  inv1  gate917(.a(N1712), .O(gate499inter8));
  nand2 gate918(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate919(.a(s_5), .b(gate499inter3), .O(gate499inter10));
  nor2  gate920(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate921(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate922(.a(gate499inter12), .b(gate499inter1), .O(N1748));
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );

  xor2  gate1693(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate1694(.a(gate508inter0), .b(s_116), .O(gate508inter1));
  and2  gate1695(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate1696(.a(s_116), .O(gate508inter3));
  inv1  gate1697(.a(s_117), .O(gate508inter4));
  nand2 gate1698(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1699(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1700(.a(N1723), .O(gate508inter7));
  inv1  gate1701(.a(N1413), .O(gate508inter8));
  nand2 gate1702(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1703(.a(s_117), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1704(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1705(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1706(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );

  xor2  gate1427(.a(N1746), .b(N1708), .O(gate510inter0));
  nand2 gate1428(.a(gate510inter0), .b(s_78), .O(gate510inter1));
  and2  gate1429(.a(N1746), .b(N1708), .O(gate510inter2));
  inv1  gate1430(.a(s_78), .O(gate510inter3));
  inv1  gate1431(.a(s_79), .O(gate510inter4));
  nand2 gate1432(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1433(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1434(.a(N1708), .O(gate510inter7));
  inv1  gate1435(.a(N1746), .O(gate510inter8));
  nand2 gate1436(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1437(.a(s_79), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1438(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1439(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1440(.a(gate510inter12), .b(gate510inter1), .O(N1774));
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1665(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1666(.a(gate513inter0), .b(s_112), .O(gate513inter1));
  and2  gate1667(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1668(.a(s_112), .O(gate513inter3));
  inv1  gate1669(.a(s_113), .O(gate513inter4));
  nand2 gate1670(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1671(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1672(.a(N1731), .O(gate513inter7));
  inv1  gate1673(.a(N1682), .O(gate513inter8));
  nand2 gate1674(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1675(.a(s_113), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1676(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1677(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1678(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );

  xor2  gate2127(.a(N1683), .b(N1734), .O(gate516inter0));
  nand2 gate2128(.a(gate516inter0), .b(s_178), .O(gate516inter1));
  and2  gate2129(.a(N1683), .b(N1734), .O(gate516inter2));
  inv1  gate2130(.a(s_178), .O(gate516inter3));
  inv1  gate2131(.a(s_179), .O(gate516inter4));
  nand2 gate2132(.a(gate516inter4), .b(gate516inter3), .O(gate516inter5));
  nor2  gate2133(.a(gate516inter5), .b(gate516inter2), .O(gate516inter6));
  inv1  gate2134(.a(N1734), .O(gate516inter7));
  inv1  gate2135(.a(N1683), .O(gate516inter8));
  nand2 gate2136(.a(gate516inter8), .b(gate516inter7), .O(gate516inter9));
  nand2 gate2137(.a(s_179), .b(gate516inter3), .O(gate516inter10));
  nor2  gate2138(.a(gate516inter10), .b(gate516inter9), .O(gate516inter11));
  nor2  gate2139(.a(gate516inter11), .b(gate516inter6), .O(gate516inter12));
  nand2 gate2140(.a(gate516inter12), .b(gate516inter1), .O(N1787));
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );

  xor2  gate1623(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate1624(.a(gate520inter0), .b(s_106), .O(gate520inter1));
  and2  gate1625(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate1626(.a(s_106), .O(gate520inter3));
  inv1  gate1627(.a(s_107), .O(gate520inter4));
  nand2 gate1628(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate1629(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate1630(.a(N1751), .O(gate520inter7));
  inv1  gate1631(.a(N1155), .O(gate520inter8));
  nand2 gate1632(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate1633(.a(s_107), .b(gate520inter3), .O(gate520inter10));
  nor2  gate1634(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate1635(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate1636(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate1679(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate1680(.a(gate522inter0), .b(s_114), .O(gate522inter1));
  and2  gate1681(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate1682(.a(s_114), .O(gate522inter3));
  inv1  gate1683(.a(s_115), .O(gate522inter4));
  nand2 gate1684(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate1685(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate1686(.a(N1740), .O(gate522inter7));
  inv1  gate1687(.a(N1769), .O(gate522inter8));
  nand2 gate1688(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate1689(.a(s_115), .b(gate522inter3), .O(gate522inter10));
  nor2  gate1690(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate1691(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate1692(.a(gate522inter12), .b(gate522inter1), .O(N1798));

  xor2  gate1217(.a(N1773), .b(N1334), .O(gate523inter0));
  nand2 gate1218(.a(gate523inter0), .b(s_48), .O(gate523inter1));
  and2  gate1219(.a(N1773), .b(N1334), .O(gate523inter2));
  inv1  gate1220(.a(s_48), .O(gate523inter3));
  inv1  gate1221(.a(s_49), .O(gate523inter4));
  nand2 gate1222(.a(gate523inter4), .b(gate523inter3), .O(gate523inter5));
  nor2  gate1223(.a(gate523inter5), .b(gate523inter2), .O(gate523inter6));
  inv1  gate1224(.a(N1334), .O(gate523inter7));
  inv1  gate1225(.a(N1773), .O(gate523inter8));
  nand2 gate1226(.a(gate523inter8), .b(gate523inter7), .O(gate523inter9));
  nand2 gate1227(.a(s_49), .b(gate523inter3), .O(gate523inter10));
  nor2  gate1228(.a(gate523inter10), .b(gate523inter9), .O(gate523inter11));
  nor2  gate1229(.a(gate523inter11), .b(gate523inter6), .O(gate523inter12));
  nand2 gate1230(.a(gate523inter12), .b(gate523inter1), .O(N1801));
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );

  xor2  gate1175(.a(N1218), .b(N1748), .O(gate526inter0));
  nand2 gate1176(.a(gate526inter0), .b(s_42), .O(gate526inter1));
  and2  gate1177(.a(N1218), .b(N1748), .O(gate526inter2));
  inv1  gate1178(.a(s_42), .O(gate526inter3));
  inv1  gate1179(.a(s_43), .O(gate526inter4));
  nand2 gate1180(.a(gate526inter4), .b(gate526inter3), .O(gate526inter5));
  nor2  gate1181(.a(gate526inter5), .b(gate526inter2), .O(gate526inter6));
  inv1  gate1182(.a(N1748), .O(gate526inter7));
  inv1  gate1183(.a(N1218), .O(gate526inter8));
  nand2 gate1184(.a(gate526inter8), .b(gate526inter7), .O(gate526inter9));
  nand2 gate1185(.a(s_43), .b(gate526inter3), .O(gate526inter10));
  nor2  gate1186(.a(gate526inter10), .b(gate526inter9), .O(gate526inter11));
  nor2  gate1187(.a(gate526inter11), .b(gate526inter6), .O(gate526inter12));
  nand2 gate1188(.a(gate526inter12), .b(gate526inter1), .O(N1808));
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate2239(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate2240(.a(gate532inter0), .b(s_194), .O(gate532inter1));
  and2  gate2241(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate2242(.a(s_194), .O(gate532inter3));
  inv1  gate2243(.a(s_195), .O(gate532inter4));
  nand2 gate2244(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate2245(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate2246(.a(N1777), .O(gate532inter7));
  inv1  gate2247(.a(N1490), .O(gate532inter8));
  nand2 gate2248(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate2249(.a(s_195), .b(gate532inter3), .O(gate532inter10));
  nor2  gate2250(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate2251(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate2252(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );

  xor2  gate1441(.a(N1491), .b(N1774), .O(gate534inter0));
  nand2 gate1442(.a(gate534inter0), .b(s_80), .O(gate534inter1));
  and2  gate1443(.a(N1491), .b(N1774), .O(gate534inter2));
  inv1  gate1444(.a(s_80), .O(gate534inter3));
  inv1  gate1445(.a(s_81), .O(gate534inter4));
  nand2 gate1446(.a(gate534inter4), .b(gate534inter3), .O(gate534inter5));
  nor2  gate1447(.a(gate534inter5), .b(gate534inter2), .O(gate534inter6));
  inv1  gate1448(.a(N1774), .O(gate534inter7));
  inv1  gate1449(.a(N1491), .O(gate534inter8));
  nand2 gate1450(.a(gate534inter8), .b(gate534inter7), .O(gate534inter9));
  nand2 gate1451(.a(s_81), .b(gate534inter3), .O(gate534inter10));
  nor2  gate1452(.a(gate534inter10), .b(gate534inter9), .O(gate534inter11));
  nor2  gate1453(.a(gate534inter11), .b(gate534inter6), .O(gate534inter12));
  nand2 gate1454(.a(gate534inter12), .b(gate534inter1), .O(N1823));
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );

  xor2  gate1553(.a(N1807), .b(N959), .O(gate540inter0));
  nand2 gate1554(.a(gate540inter0), .b(s_96), .O(gate540inter1));
  and2  gate1555(.a(N1807), .b(N959), .O(gate540inter2));
  inv1  gate1556(.a(s_96), .O(gate540inter3));
  inv1  gate1557(.a(s_97), .O(gate540inter4));
  nand2 gate1558(.a(gate540inter4), .b(gate540inter3), .O(gate540inter5));
  nor2  gate1559(.a(gate540inter5), .b(gate540inter2), .O(gate540inter6));
  inv1  gate1560(.a(N959), .O(gate540inter7));
  inv1  gate1561(.a(N1807), .O(gate540inter8));
  nand2 gate1562(.a(gate540inter8), .b(gate540inter7), .O(gate540inter9));
  nand2 gate1563(.a(s_97), .b(gate540inter3), .O(gate540inter10));
  nor2  gate1564(.a(gate540inter10), .b(gate540inter9), .O(gate540inter11));
  nor2  gate1565(.a(gate540inter11), .b(gate540inter6), .O(gate540inter12));
  nand2 gate1566(.a(gate540inter12), .b(gate540inter1), .O(N1837));
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );

  xor2  gate1917(.a(N1822), .b(N1419), .O(gate543inter0));
  nand2 gate1918(.a(gate543inter0), .b(s_148), .O(gate543inter1));
  and2  gate1919(.a(N1822), .b(N1419), .O(gate543inter2));
  inv1  gate1920(.a(s_148), .O(gate543inter3));
  inv1  gate1921(.a(s_149), .O(gate543inter4));
  nand2 gate1922(.a(gate543inter4), .b(gate543inter3), .O(gate543inter5));
  nor2  gate1923(.a(gate543inter5), .b(gate543inter2), .O(gate543inter6));
  inv1  gate1924(.a(N1419), .O(gate543inter7));
  inv1  gate1925(.a(N1822), .O(gate543inter8));
  nand2 gate1926(.a(gate543inter8), .b(gate543inter7), .O(gate543inter9));
  nand2 gate1927(.a(s_149), .b(gate543inter3), .O(gate543inter10));
  nor2  gate1928(.a(gate543inter10), .b(gate543inter9), .O(gate543inter11));
  nor2  gate1929(.a(gate543inter11), .b(gate543inter6), .O(gate543inter12));
  nand2 gate1930(.a(gate543inter12), .b(gate543inter1), .O(N1848));

  xor2  gate923(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate924(.a(gate544inter0), .b(s_6), .O(gate544inter1));
  and2  gate925(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate926(.a(s_6), .O(gate544inter3));
  inv1  gate927(.a(s_7), .O(gate544inter4));
  nand2 gate928(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate929(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate930(.a(N1416), .O(gate544inter7));
  inv1  gate931(.a(N1824), .O(gate544inter8));
  nand2 gate932(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate933(.a(s_7), .b(gate544inter3), .O(gate544inter10));
  nor2  gate934(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate935(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate936(.a(gate544inter12), .b(gate544inter1), .O(N1849));
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );

  xor2  gate2281(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate2282(.a(gate546inter0), .b(s_200), .O(gate546inter1));
  and2  gate2283(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate2284(.a(s_200), .O(gate546inter3));
  inv1  gate2285(.a(s_201), .O(gate546inter4));
  nand2 gate2286(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate2287(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate2288(.a(N1319), .O(gate546inter7));
  inv1  gate2289(.a(N1827), .O(gate546inter8));
  nand2 gate2290(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate2291(.a(s_201), .b(gate546inter3), .O(gate546inter10));
  nor2  gate2292(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate2293(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate2294(.a(gate546inter12), .b(gate546inter1), .O(N1852));
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );

  xor2  gate965(.a(N290), .b(N1798), .O(gate550inter0));
  nand2 gate966(.a(gate550inter0), .b(s_12), .O(gate550inter1));
  and2  gate967(.a(N290), .b(N1798), .O(gate550inter2));
  inv1  gate968(.a(s_12), .O(gate550inter3));
  inv1  gate969(.a(s_13), .O(gate550inter4));
  nand2 gate970(.a(gate550inter4), .b(gate550inter3), .O(gate550inter5));
  nor2  gate971(.a(gate550inter5), .b(gate550inter2), .O(gate550inter6));
  inv1  gate972(.a(N1798), .O(gate550inter7));
  inv1  gate973(.a(N290), .O(gate550inter8));
  nand2 gate974(.a(gate550inter8), .b(gate550inter7), .O(gate550inter9));
  nand2 gate975(.a(s_13), .b(gate550inter3), .O(gate550inter10));
  nor2  gate976(.a(gate550inter10), .b(gate550inter9), .O(gate550inter11));
  nor2  gate977(.a(gate550inter11), .b(gate550inter6), .O(gate550inter12));
  nand2 gate978(.a(gate550inter12), .b(gate550inter1), .O(N1858));
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );

  xor2  gate1147(.a(N1848), .b(N1821), .O(gate557inter0));
  nand2 gate1148(.a(gate557inter0), .b(s_38), .O(gate557inter1));
  and2  gate1149(.a(N1848), .b(N1821), .O(gate557inter2));
  inv1  gate1150(.a(s_38), .O(gate557inter3));
  inv1  gate1151(.a(s_39), .O(gate557inter4));
  nand2 gate1152(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate1153(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate1154(.a(N1821), .O(gate557inter7));
  inv1  gate1155(.a(N1848), .O(gate557inter8));
  nand2 gate1156(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate1157(.a(s_39), .b(gate557inter3), .O(gate557inter10));
  nor2  gate1158(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate1159(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate1160(.a(gate557inter12), .b(gate557inter1), .O(N1878));
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );

  xor2  gate1861(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate1862(.a(gate562inter0), .b(s_140), .O(gate562inter1));
  and2  gate1863(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate1864(.a(s_140), .O(gate562inter3));
  inv1  gate1865(.a(s_141), .O(gate562inter4));
  nand2 gate1866(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate1867(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate1868(.a(N1643), .O(gate562inter7));
  inv1  gate1869(.a(N1856), .O(gate562inter8));
  nand2 gate1870(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate1871(.a(s_141), .b(gate562inter3), .O(gate562inter10));
  nor2  gate1872(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate1873(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate1874(.a(gate562inter12), .b(gate562inter1), .O(N1885));
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate1077(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate1078(.a(gate574inter0), .b(s_28), .O(gate574inter1));
  and2  gate1079(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate1080(.a(s_28), .O(gate574inter3));
  inv1  gate1081(.a(s_29), .O(gate574inter4));
  nand2 gate1082(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate1083(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate1084(.a(N1872), .O(gate574inter7));
  inv1  gate1085(.a(N919), .O(gate574inter8));
  nand2 gate1086(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate1087(.a(s_29), .b(gate574inter3), .O(gate574inter10));
  nor2  gate1088(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate1089(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate1090(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate1721(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate1722(.a(gate579inter0), .b(s_120), .O(gate579inter1));
  and2  gate1723(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate1724(.a(s_120), .O(gate579inter3));
  inv1  gate1725(.a(s_121), .O(gate579inter4));
  nand2 gate1726(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate1727(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate1728(.a(N1714), .O(gate579inter7));
  inv1  gate1729(.a(N1895), .O(gate579inter8));
  nand2 gate1730(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate1731(.a(s_121), .b(gate579inter3), .O(gate579inter10));
  nor2  gate1732(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate1733(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate1734(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );

  xor2  gate2267(.a(N1911), .b(N1882), .O(gate583inter0));
  nand2 gate2268(.a(gate583inter0), .b(s_198), .O(gate583inter1));
  and2  gate2269(.a(N1911), .b(N1882), .O(gate583inter2));
  inv1  gate2270(.a(s_198), .O(gate583inter3));
  inv1  gate2271(.a(s_199), .O(gate583inter4));
  nand2 gate2272(.a(gate583inter4), .b(gate583inter3), .O(gate583inter5));
  nor2  gate2273(.a(gate583inter5), .b(gate583inter2), .O(gate583inter6));
  inv1  gate2274(.a(N1882), .O(gate583inter7));
  inv1  gate2275(.a(N1911), .O(gate583inter8));
  nand2 gate2276(.a(gate583inter8), .b(gate583inter7), .O(gate583inter9));
  nand2 gate2277(.a(s_199), .b(gate583inter3), .O(gate583inter10));
  nor2  gate2278(.a(gate583inter10), .b(gate583inter9), .O(gate583inter11));
  nor2  gate2279(.a(gate583inter11), .b(gate583inter6), .O(gate583inter12));
  nand2 gate2280(.a(gate583inter12), .b(gate583inter1), .O(N1936));
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );

  xor2  gate1287(.a(N1922), .b(N676), .O(gate587inter0));
  nand2 gate1288(.a(gate587inter0), .b(s_58), .O(gate587inter1));
  and2  gate1289(.a(N1922), .b(N676), .O(gate587inter2));
  inv1  gate1290(.a(s_58), .O(gate587inter3));
  inv1  gate1291(.a(s_59), .O(gate587inter4));
  nand2 gate1292(.a(gate587inter4), .b(gate587inter3), .O(gate587inter5));
  nor2  gate1293(.a(gate587inter5), .b(gate587inter2), .O(gate587inter6));
  inv1  gate1294(.a(N676), .O(gate587inter7));
  inv1  gate1295(.a(N1922), .O(gate587inter8));
  nand2 gate1296(.a(gate587inter8), .b(gate587inter7), .O(gate587inter9));
  nand2 gate1297(.a(s_59), .b(gate587inter3), .O(gate587inter10));
  nor2  gate1298(.a(gate587inter10), .b(gate587inter9), .O(gate587inter11));
  nor2  gate1299(.a(gate587inter11), .b(gate587inter6), .O(gate587inter12));
  nand2 gate1300(.a(gate587inter12), .b(gate587inter1), .O(N1942));
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );

  xor2  gate1049(.a(N1941), .b(N1919), .O(gate600inter0));
  nand2 gate1050(.a(gate600inter0), .b(s_24), .O(gate600inter1));
  and2  gate1051(.a(N1941), .b(N1919), .O(gate600inter2));
  inv1  gate1052(.a(s_24), .O(gate600inter3));
  inv1  gate1053(.a(s_25), .O(gate600inter4));
  nand2 gate1054(.a(gate600inter4), .b(gate600inter3), .O(gate600inter5));
  nor2  gate1055(.a(gate600inter5), .b(gate600inter2), .O(gate600inter6));
  inv1  gate1056(.a(N1919), .O(gate600inter7));
  inv1  gate1057(.a(N1941), .O(gate600inter8));
  nand2 gate1058(.a(gate600inter8), .b(gate600inter7), .O(gate600inter9));
  nand2 gate1059(.a(s_25), .b(gate600inter3), .O(gate600inter10));
  nor2  gate1060(.a(gate600inter10), .b(gate600inter9), .O(gate600inter11));
  nor2  gate1061(.a(gate600inter11), .b(gate600inter6), .O(gate600inter12));
  nand2 gate1062(.a(gate600inter12), .b(gate600inter1), .O(N1979));
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );

  xor2  gate1581(.a(N1351), .b(N1950), .O(gate610inter0));
  nand2 gate1582(.a(gate610inter0), .b(s_100), .O(gate610inter1));
  and2  gate1583(.a(N1351), .b(N1950), .O(gate610inter2));
  inv1  gate1584(.a(s_100), .O(gate610inter3));
  inv1  gate1585(.a(s_101), .O(gate610inter4));
  nand2 gate1586(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate1587(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate1588(.a(N1950), .O(gate610inter7));
  inv1  gate1589(.a(N1351), .O(gate610inter8));
  nand2 gate1590(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate1591(.a(s_101), .b(gate610inter3), .O(gate610inter10));
  nor2  gate1592(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate1593(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate1594(.a(gate610inter12), .b(gate610inter1), .O(N2006));
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate1847(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate1848(.a(gate612inter0), .b(s_138), .O(gate612inter1));
  and2  gate1849(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate1850(.a(s_138), .O(gate612inter3));
  inv1  gate1851(.a(s_139), .O(gate612inter4));
  nand2 gate1852(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate1853(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate1854(.a(N673), .O(gate612inter7));
  inv1  gate1855(.a(N1976), .O(gate612inter8));
  nand2 gate1856(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate1857(.a(s_139), .b(gate612inter3), .O(gate612inter10));
  nor2  gate1858(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate1859(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate1860(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );

  xor2  gate895(.a(N1591), .b(N1987), .O(gate623inter0));
  nand2 gate896(.a(gate623inter0), .b(s_2), .O(gate623inter1));
  and2  gate897(.a(N1591), .b(N1987), .O(gate623inter2));
  inv1  gate898(.a(s_2), .O(gate623inter3));
  inv1  gate899(.a(s_3), .O(gate623inter4));
  nand2 gate900(.a(gate623inter4), .b(gate623inter3), .O(gate623inter5));
  nor2  gate901(.a(gate623inter5), .b(gate623inter2), .O(gate623inter6));
  inv1  gate902(.a(N1987), .O(gate623inter7));
  inv1  gate903(.a(N1591), .O(gate623inter8));
  nand2 gate904(.a(gate623inter8), .b(gate623inter7), .O(gate623inter9));
  nand2 gate905(.a(s_3), .b(gate623inter3), .O(gate623inter10));
  nor2  gate906(.a(gate623inter10), .b(gate623inter9), .O(gate623inter11));
  nor2  gate907(.a(gate623inter11), .b(gate623inter6), .O(gate623inter12));
  nand2 gate908(.a(gate623inter12), .b(gate623inter1), .O(N2022));
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );

  xor2  gate1413(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate1414(.a(gate627inter0), .b(s_76), .O(gate627inter1));
  and2  gate1415(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate1416(.a(s_76), .O(gate627inter3));
  inv1  gate1417(.a(s_77), .O(gate627inter4));
  nand2 gate1418(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate1419(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate1420(.a(N1975), .O(gate627inter7));
  inv1  gate1421(.a(N2008), .O(gate627inter8));
  nand2 gate1422(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate1423(.a(s_77), .b(gate627inter3), .O(gate627inter10));
  nor2  gate1424(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate1425(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate1426(.a(gate627inter12), .b(gate627inter1), .O(N2026));

  xor2  gate1035(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1036(.a(gate628inter0), .b(s_22), .O(gate628inter1));
  and2  gate1037(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1038(.a(s_22), .O(gate628inter3));
  inv1  gate1039(.a(s_23), .O(gate628inter4));
  nand2 gate1040(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1041(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1042(.a(N1977), .O(gate628inter7));
  inv1  gate1043(.a(N2009), .O(gate628inter8));
  nand2 gate1044(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1045(.a(s_23), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1046(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1047(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1048(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate1777(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate1778(.a(gate633inter0), .b(s_128), .O(gate633inter1));
  and2  gate1779(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate1780(.a(s_128), .O(gate633inter3));
  inv1  gate1781(.a(s_129), .O(gate633inter4));
  nand2 gate1782(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate1783(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate1784(.a(N2020), .O(gate633inter7));
  inv1  gate1785(.a(N2000), .O(gate633inter8));
  nand2 gate1786(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate1787(.a(s_129), .b(gate633inter3), .O(gate633inter10));
  nor2  gate1788(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate1789(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate1790(.a(gate633inter12), .b(gate633inter1), .O(N2038));

  xor2  gate1483(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate1484(.a(gate634inter0), .b(s_86), .O(gate634inter1));
  and2  gate1485(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate1486(.a(s_86), .O(gate634inter3));
  inv1  gate1487(.a(s_87), .O(gate634inter4));
  nand2 gate1488(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate1489(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate1490(.a(N1534), .O(gate634inter7));
  inv1  gate1491(.a(N2021), .O(gate634inter8));
  nand2 gate1492(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate1493(.a(s_87), .b(gate634inter3), .O(gate634inter10));
  nor2  gate1494(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate1495(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate1496(.a(gate634inter12), .b(gate634inter1), .O(N2039));
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );

  xor2  gate1315(.a(N2025), .b(N2006), .O(gate637inter0));
  nand2 gate1316(.a(gate637inter0), .b(s_62), .O(gate637inter1));
  and2  gate1317(.a(N2025), .b(N2006), .O(gate637inter2));
  inv1  gate1318(.a(s_62), .O(gate637inter3));
  inv1  gate1319(.a(s_63), .O(gate637inter4));
  nand2 gate1320(.a(gate637inter4), .b(gate637inter3), .O(gate637inter5));
  nor2  gate1321(.a(gate637inter5), .b(gate637inter2), .O(gate637inter6));
  inv1  gate1322(.a(N2006), .O(gate637inter7));
  inv1  gate1323(.a(N2025), .O(gate637inter8));
  nand2 gate1324(.a(gate637inter8), .b(gate637inter7), .O(gate637inter9));
  nand2 gate1325(.a(s_63), .b(gate637inter3), .O(gate637inter10));
  nor2  gate1326(.a(gate637inter10), .b(gate637inter9), .O(gate637inter11));
  nor2  gate1327(.a(gate637inter11), .b(gate637inter6), .O(gate637inter12));
  nand2 gate1328(.a(gate637inter12), .b(gate637inter1), .O(N2042));
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );

  xor2  gate2211(.a(N2016), .b(N2037), .O(gate640inter0));
  nand2 gate2212(.a(gate640inter0), .b(s_190), .O(gate640inter1));
  and2  gate2213(.a(N2016), .b(N2037), .O(gate640inter2));
  inv1  gate2214(.a(s_190), .O(gate640inter3));
  inv1  gate2215(.a(s_191), .O(gate640inter4));
  nand2 gate2216(.a(gate640inter4), .b(gate640inter3), .O(gate640inter5));
  nor2  gate2217(.a(gate640inter5), .b(gate640inter2), .O(gate640inter6));
  inv1  gate2218(.a(N2037), .O(gate640inter7));
  inv1  gate2219(.a(N2016), .O(gate640inter8));
  nand2 gate2220(.a(gate640inter8), .b(gate640inter7), .O(gate640inter9));
  nand2 gate2221(.a(s_191), .b(gate640inter3), .O(gate640inter10));
  nor2  gate2222(.a(gate640inter10), .b(gate640inter9), .O(gate640inter11));
  nor2  gate2223(.a(gate640inter11), .b(gate640inter6), .O(gate640inter12));
  nand2 gate2224(.a(gate640inter12), .b(gate640inter1), .O(N2055));
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate2099(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate2100(.a(gate667inter0), .b(s_174), .O(gate667inter1));
  and2  gate2101(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate2102(.a(s_174), .O(gate667inter3));
  inv1  gate2103(.a(s_175), .O(gate667inter4));
  nand2 gate2104(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate2105(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate2106(.a(N2199), .O(gate667inter7));
  inv1  gate2107(.a(N1348), .O(gate667inter8));
  nand2 gate2108(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate2109(.a(s_175), .b(gate667inter3), .O(gate667inter10));
  nor2  gate2110(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate2111(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate2112(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );

  xor2  gate979(.a(N1349), .b(N2196), .O(gate669inter0));
  nand2 gate980(.a(gate669inter0), .b(s_14), .O(gate669inter1));
  and2  gate981(.a(N1349), .b(N2196), .O(gate669inter2));
  inv1  gate982(.a(s_14), .O(gate669inter3));
  inv1  gate983(.a(s_15), .O(gate669inter4));
  nand2 gate984(.a(gate669inter4), .b(gate669inter3), .O(gate669inter5));
  nor2  gate985(.a(gate669inter5), .b(gate669inter2), .O(gate669inter6));
  inv1  gate986(.a(N2196), .O(gate669inter7));
  inv1  gate987(.a(N1349), .O(gate669inter8));
  nand2 gate988(.a(gate669inter8), .b(gate669inter7), .O(gate669inter9));
  nand2 gate989(.a(s_15), .b(gate669inter3), .O(gate669inter10));
  nor2  gate990(.a(gate669inter10), .b(gate669inter9), .O(gate669inter11));
  nor2  gate991(.a(gate669inter11), .b(gate669inter6), .O(gate669inter12));
  nand2 gate992(.a(gate669inter12), .b(gate669inter1), .O(N2224));
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate1119(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate1120(.a(gate671inter0), .b(s_34), .O(gate671inter1));
  and2  gate1121(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate1122(.a(s_34), .O(gate671inter3));
  inv1  gate1123(.a(s_35), .O(gate671inter4));
  nand2 gate1124(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate1125(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate1126(.a(N2205), .O(gate671inter7));
  inv1  gate1127(.a(N913), .O(gate671inter8));
  nand2 gate1128(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate1129(.a(s_35), .b(gate671inter3), .O(gate671inter10));
  nor2  gate1130(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate1131(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate1132(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate1399(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate1400(.a(gate754inter0), .b(s_74), .O(gate754inter1));
  and2  gate1401(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate1402(.a(s_74), .O(gate754inter3));
  inv1  gate1403(.a(s_75), .O(gate754inter4));
  nand2 gate1404(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1405(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1406(.a(N2564), .O(gate754inter7));
  inv1  gate1407(.a(N536), .O(gate754inter8));
  nand2 gate1408(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1409(.a(s_75), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1410(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1411(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1412(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );

  xor2  gate2113(.a(N548), .b(N2573), .O(gate760inter0));
  nand2 gate2114(.a(gate760inter0), .b(s_176), .O(gate760inter1));
  and2  gate2115(.a(N548), .b(N2573), .O(gate760inter2));
  inv1  gate2116(.a(s_176), .O(gate760inter3));
  inv1  gate2117(.a(s_177), .O(gate760inter4));
  nand2 gate2118(.a(gate760inter4), .b(gate760inter3), .O(gate760inter5));
  nor2  gate2119(.a(gate760inter5), .b(gate760inter2), .O(gate760inter6));
  inv1  gate2120(.a(N2573), .O(gate760inter7));
  inv1  gate2121(.a(N548), .O(gate760inter8));
  nand2 gate2122(.a(gate760inter8), .b(gate760inter7), .O(gate760inter9));
  nand2 gate2123(.a(s_177), .b(gate760inter3), .O(gate760inter10));
  nor2  gate2124(.a(gate760inter10), .b(gate760inter9), .O(gate760inter11));
  nor2  gate2125(.a(gate760inter11), .b(gate760inter6), .O(gate760inter12));
  nand2 gate2126(.a(gate760inter12), .b(gate760inter1), .O(N2688));
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );

  xor2  gate2071(.a(N2672), .b(N346), .O(gate766inter0));
  nand2 gate2072(.a(gate766inter0), .b(s_170), .O(gate766inter1));
  and2  gate2073(.a(N2672), .b(N346), .O(gate766inter2));
  inv1  gate2074(.a(s_170), .O(gate766inter3));
  inv1  gate2075(.a(s_171), .O(gate766inter4));
  nand2 gate2076(.a(gate766inter4), .b(gate766inter3), .O(gate766inter5));
  nor2  gate2077(.a(gate766inter5), .b(gate766inter2), .O(gate766inter6));
  inv1  gate2078(.a(N346), .O(gate766inter7));
  inv1  gate2079(.a(N2672), .O(gate766inter8));
  nand2 gate2080(.a(gate766inter8), .b(gate766inter7), .O(gate766inter9));
  nand2 gate2081(.a(s_171), .b(gate766inter3), .O(gate766inter10));
  nor2  gate2082(.a(gate766inter10), .b(gate766inter9), .O(gate766inter11));
  nor2  gate2083(.a(gate766inter11), .b(gate766inter6), .O(gate766inter12));
  nand2 gate2084(.a(gate766inter12), .b(gate766inter1), .O(N2721));
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate1259(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate1260(.a(gate773inter0), .b(s_54), .O(gate773inter1));
  and2  gate1261(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate1262(.a(s_54), .O(gate773inter3));
  inv1  gate1263(.a(s_55), .O(gate773inter4));
  nand2 gate1264(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate1265(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate1266(.a(N2645), .O(gate773inter7));
  inv1  gate1267(.a(N540), .O(gate773inter8));
  nand2 gate1268(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate1269(.a(s_55), .b(gate773inter3), .O(gate773inter10));
  nor2  gate1270(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate1271(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate1272(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );

  xor2  gate1637(.a(N541), .b(N2648), .O(gate775inter0));
  nand2 gate1638(.a(gate775inter0), .b(s_108), .O(gate775inter1));
  and2  gate1639(.a(N541), .b(N2648), .O(gate775inter2));
  inv1  gate1640(.a(s_108), .O(gate775inter3));
  inv1  gate1641(.a(s_109), .O(gate775inter4));
  nand2 gate1642(.a(gate775inter4), .b(gate775inter3), .O(gate775inter5));
  nor2  gate1643(.a(gate775inter5), .b(gate775inter2), .O(gate775inter6));
  inv1  gate1644(.a(N2648), .O(gate775inter7));
  inv1  gate1645(.a(N541), .O(gate775inter8));
  nand2 gate1646(.a(gate775inter8), .b(gate775inter7), .O(gate775inter9));
  nand2 gate1647(.a(s_109), .b(gate775inter3), .O(gate775inter10));
  nor2  gate1648(.a(gate775inter10), .b(gate775inter9), .O(gate775inter11));
  nor2  gate1649(.a(gate775inter11), .b(gate775inter6), .O(gate775inter12));
  nand2 gate1650(.a(gate775inter12), .b(gate775inter1), .O(N2730));
inv1 gate776( .a(N2648), .O(N2731) );

  xor2  gate1987(.a(N542), .b(N2651), .O(gate777inter0));
  nand2 gate1988(.a(gate777inter0), .b(s_158), .O(gate777inter1));
  and2  gate1989(.a(N542), .b(N2651), .O(gate777inter2));
  inv1  gate1990(.a(s_158), .O(gate777inter3));
  inv1  gate1991(.a(s_159), .O(gate777inter4));
  nand2 gate1992(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate1993(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate1994(.a(N2651), .O(gate777inter7));
  inv1  gate1995(.a(N542), .O(gate777inter8));
  nand2 gate1996(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate1997(.a(s_159), .b(gate777inter3), .O(gate777inter10));
  nor2  gate1998(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate1999(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate2000(.a(gate777inter12), .b(gate777inter1), .O(N2732));
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );

  xor2  gate993(.a(N2691), .b(N388), .O(gate789inter0));
  nand2 gate994(.a(gate789inter0), .b(s_16), .O(gate789inter1));
  and2  gate995(.a(N2691), .b(N388), .O(gate789inter2));
  inv1  gate996(.a(s_16), .O(gate789inter3));
  inv1  gate997(.a(s_17), .O(gate789inter4));
  nand2 gate998(.a(gate789inter4), .b(gate789inter3), .O(gate789inter5));
  nor2  gate999(.a(gate789inter5), .b(gate789inter2), .O(gate789inter6));
  inv1  gate1000(.a(N388), .O(gate789inter7));
  inv1  gate1001(.a(N2691), .O(gate789inter8));
  nand2 gate1002(.a(gate789inter8), .b(gate789inter7), .O(gate789inter9));
  nand2 gate1003(.a(s_17), .b(gate789inter3), .O(gate789inter10));
  nor2  gate1004(.a(gate789inter10), .b(gate789inter9), .O(gate789inter11));
  nor2  gate1005(.a(gate789inter11), .b(gate789inter6), .O(gate789inter12));
  nand2 gate1006(.a(gate789inter12), .b(gate789inter1), .O(N2744));
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );

  xor2  gate2001(.a(N2720), .b(N2669), .O(gate794inter0));
  nand2 gate2002(.a(gate794inter0), .b(s_160), .O(gate794inter1));
  and2  gate2003(.a(N2720), .b(N2669), .O(gate794inter2));
  inv1  gate2004(.a(s_160), .O(gate794inter3));
  inv1  gate2005(.a(s_161), .O(gate794inter4));
  nand2 gate2006(.a(gate794inter4), .b(gate794inter3), .O(gate794inter5));
  nor2  gate2007(.a(gate794inter5), .b(gate794inter2), .O(gate794inter6));
  inv1  gate2008(.a(N2669), .O(gate794inter7));
  inv1  gate2009(.a(N2720), .O(gate794inter8));
  nand2 gate2010(.a(gate794inter8), .b(gate794inter7), .O(gate794inter9));
  nand2 gate2011(.a(s_161), .b(gate794inter3), .O(gate794inter10));
  nor2  gate2012(.a(gate794inter10), .b(gate794inter9), .O(gate794inter11));
  nor2  gate2013(.a(gate794inter11), .b(gate794inter6), .O(gate794inter12));
  nand2 gate2014(.a(gate794inter12), .b(gate794inter1), .O(N2753));
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );

  xor2  gate1301(.a(N2731), .b(N364), .O(gate801inter0));
  nand2 gate1302(.a(gate801inter0), .b(s_60), .O(gate801inter1));
  and2  gate1303(.a(N2731), .b(N364), .O(gate801inter2));
  inv1  gate1304(.a(s_60), .O(gate801inter3));
  inv1  gate1305(.a(s_61), .O(gate801inter4));
  nand2 gate1306(.a(gate801inter4), .b(gate801inter3), .O(gate801inter5));
  nor2  gate1307(.a(gate801inter5), .b(gate801inter2), .O(gate801inter6));
  inv1  gate1308(.a(N364), .O(gate801inter7));
  inv1  gate1309(.a(N2731), .O(gate801inter8));
  nand2 gate1310(.a(gate801inter8), .b(gate801inter7), .O(gate801inter9));
  nand2 gate1311(.a(s_61), .b(gate801inter3), .O(gate801inter10));
  nor2  gate1312(.a(gate801inter10), .b(gate801inter9), .O(gate801inter11));
  nor2  gate1313(.a(gate801inter11), .b(gate801inter6), .O(gate801inter12));
  nand2 gate1314(.a(gate801inter12), .b(gate801inter1), .O(N2760));

  xor2  gate2183(.a(N2733), .b(N367), .O(gate802inter0));
  nand2 gate2184(.a(gate802inter0), .b(s_186), .O(gate802inter1));
  and2  gate2185(.a(N2733), .b(N367), .O(gate802inter2));
  inv1  gate2186(.a(s_186), .O(gate802inter3));
  inv1  gate2187(.a(s_187), .O(gate802inter4));
  nand2 gate2188(.a(gate802inter4), .b(gate802inter3), .O(gate802inter5));
  nor2  gate2189(.a(gate802inter5), .b(gate802inter2), .O(gate802inter6));
  inv1  gate2190(.a(N367), .O(gate802inter7));
  inv1  gate2191(.a(N2733), .O(gate802inter8));
  nand2 gate2192(.a(gate802inter8), .b(gate802inter7), .O(gate802inter9));
  nand2 gate2193(.a(s_187), .b(gate802inter3), .O(gate802inter10));
  nor2  gate2194(.a(gate802inter10), .b(gate802inter9), .O(gate802inter11));
  nor2  gate2195(.a(gate802inter11), .b(gate802inter6), .O(gate802inter12));
  nand2 gate2196(.a(gate802inter12), .b(gate802inter1), .O(N2761));
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );

  xor2  gate937(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate938(.a(gate813inter0), .b(s_8), .O(gate813inter1));
  and2  gate939(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate940(.a(s_8), .O(gate813inter3));
  inv1  gate941(.a(s_9), .O(gate813inter4));
  nand2 gate942(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate943(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate944(.a(N2726), .O(gate813inter7));
  inv1  gate945(.a(N2758), .O(gate813inter8));
  nand2 gate946(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate947(.a(s_9), .b(gate813inter3), .O(gate813inter10));
  nor2  gate948(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate949(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate950(.a(gate813inter12), .b(gate813inter1), .O(N2780));
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );

  xor2  gate1497(.a(N2765), .b(N2739), .O(gate819inter0));
  nand2 gate1498(.a(gate819inter0), .b(s_88), .O(gate819inter1));
  and2  gate1499(.a(N2765), .b(N2739), .O(gate819inter2));
  inv1  gate1500(.a(s_88), .O(gate819inter3));
  inv1  gate1501(.a(s_89), .O(gate819inter4));
  nand2 gate1502(.a(gate819inter4), .b(gate819inter3), .O(gate819inter5));
  nor2  gate1503(.a(gate819inter5), .b(gate819inter2), .O(gate819inter6));
  inv1  gate1504(.a(N2739), .O(gate819inter7));
  inv1  gate1505(.a(N2765), .O(gate819inter8));
  nand2 gate1506(.a(gate819inter8), .b(gate819inter7), .O(gate819inter9));
  nand2 gate1507(.a(s_89), .b(gate819inter3), .O(gate819inter10));
  nor2  gate1508(.a(gate819inter10), .b(gate819inter9), .O(gate819inter11));
  nor2  gate1509(.a(gate819inter11), .b(gate819inter6), .O(gate819inter12));
  nand2 gate1510(.a(gate819inter12), .b(gate819inter1), .O(N2786));
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );

  xor2  gate2015(.a(N2858), .b(N2055), .O(gate852inter0));
  nand2 gate2016(.a(gate852inter0), .b(s_162), .O(gate852inter1));
  and2  gate2017(.a(N2858), .b(N2055), .O(gate852inter2));
  inv1  gate2018(.a(s_162), .O(gate852inter3));
  inv1  gate2019(.a(s_163), .O(gate852inter4));
  nand2 gate2020(.a(gate852inter4), .b(gate852inter3), .O(gate852inter5));
  nor2  gate2021(.a(gate852inter5), .b(gate852inter2), .O(gate852inter6));
  inv1  gate2022(.a(N2055), .O(gate852inter7));
  inv1  gate2023(.a(N2858), .O(gate852inter8));
  nand2 gate2024(.a(gate852inter8), .b(gate852inter7), .O(gate852inter9));
  nand2 gate2025(.a(s_163), .b(gate852inter3), .O(gate852inter10));
  nor2  gate2026(.a(gate852inter10), .b(gate852inter9), .O(gate852inter11));
  nor2  gate2027(.a(gate852inter11), .b(gate852inter6), .O(gate852inter12));
  nand2 gate2028(.a(gate852inter12), .b(gate852inter1), .O(N2867));
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );

  xor2  gate1763(.a(N2851), .b(N2867), .O(gate862inter0));
  nand2 gate1764(.a(gate862inter0), .b(s_126), .O(gate862inter1));
  and2  gate1765(.a(N2851), .b(N2867), .O(gate862inter2));
  inv1  gate1766(.a(s_126), .O(gate862inter3));
  inv1  gate1767(.a(s_127), .O(gate862inter4));
  nand2 gate1768(.a(gate862inter4), .b(gate862inter3), .O(gate862inter5));
  nor2  gate1769(.a(gate862inter5), .b(gate862inter2), .O(gate862inter6));
  inv1  gate1770(.a(N2867), .O(gate862inter7));
  inv1  gate1771(.a(N2851), .O(gate862inter8));
  nand2 gate1772(.a(gate862inter8), .b(gate862inter7), .O(gate862inter9));
  nand2 gate1773(.a(s_127), .b(gate862inter3), .O(gate862inter10));
  nor2  gate1774(.a(gate862inter10), .b(gate862inter9), .O(gate862inter11));
  nor2  gate1775(.a(gate862inter11), .b(gate862inter6), .O(gate862inter12));
  nand2 gate1776(.a(gate862inter12), .b(gate862inter1), .O(N2877));
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );

  xor2  gate2057(.a(N2853), .b(N2869), .O(gate864inter0));
  nand2 gate2058(.a(gate864inter0), .b(s_168), .O(gate864inter1));
  and2  gate2059(.a(N2853), .b(N2869), .O(gate864inter2));
  inv1  gate2060(.a(s_168), .O(gate864inter3));
  inv1  gate2061(.a(s_169), .O(gate864inter4));
  nand2 gate2062(.a(gate864inter4), .b(gate864inter3), .O(gate864inter5));
  nor2  gate2063(.a(gate864inter5), .b(gate864inter2), .O(gate864inter6));
  inv1  gate2064(.a(N2869), .O(gate864inter7));
  inv1  gate2065(.a(N2853), .O(gate864inter8));
  nand2 gate2066(.a(gate864inter8), .b(gate864inter7), .O(gate864inter9));
  nand2 gate2067(.a(s_169), .b(gate864inter3), .O(gate864inter10));
  nor2  gate2068(.a(gate864inter10), .b(gate864inter9), .O(gate864inter11));
  nor2  gate2069(.a(gate864inter11), .b(gate864inter6), .O(gate864inter12));
  nand2 gate2070(.a(gate864inter12), .b(gate864inter1), .O(N2879));

  xor2  gate1749(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate1750(.a(gate865inter0), .b(s_124), .O(gate865inter1));
  and2  gate1751(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate1752(.a(s_124), .O(gate865inter3));
  inv1  gate1753(.a(s_125), .O(gate865inter4));
  nand2 gate1754(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate1755(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate1756(.a(N2870), .O(gate865inter7));
  inv1  gate1757(.a(N2854), .O(gate865inter8));
  nand2 gate1758(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate1759(.a(s_125), .b(gate865inter3), .O(gate865inter10));
  nor2  gate1760(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate1761(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate1762(.a(gate865inter12), .b(gate865inter1), .O(N2880));
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );

  xor2  gate1973(.a(N2874), .b(N685), .O(gate867inter0));
  nand2 gate1974(.a(gate867inter0), .b(s_156), .O(gate867inter1));
  and2  gate1975(.a(N2874), .b(N685), .O(gate867inter2));
  inv1  gate1976(.a(s_156), .O(gate867inter3));
  inv1  gate1977(.a(s_157), .O(gate867inter4));
  nand2 gate1978(.a(gate867inter4), .b(gate867inter3), .O(gate867inter5));
  nor2  gate1979(.a(gate867inter5), .b(gate867inter2), .O(gate867inter6));
  inv1  gate1980(.a(N685), .O(gate867inter7));
  inv1  gate1981(.a(N2874), .O(gate867inter8));
  nand2 gate1982(.a(gate867inter8), .b(gate867inter7), .O(gate867inter9));
  nand2 gate1983(.a(s_157), .b(gate867inter3), .O(gate867inter10));
  nor2  gate1984(.a(gate867inter10), .b(gate867inter9), .O(gate867inter11));
  nor2  gate1985(.a(gate867inter11), .b(gate867inter6), .O(gate867inter12));
  nand2 gate1986(.a(gate867inter12), .b(gate867inter1), .O(N2882));
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule