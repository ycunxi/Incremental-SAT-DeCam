module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1205(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1206(.a(gate9inter0), .b(s_94), .O(gate9inter1));
  and2  gate1207(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1208(.a(s_94), .O(gate9inter3));
  inv1  gate1209(.a(s_95), .O(gate9inter4));
  nand2 gate1210(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1211(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1212(.a(G1), .O(gate9inter7));
  inv1  gate1213(.a(G2), .O(gate9inter8));
  nand2 gate1214(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1215(.a(s_95), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1216(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1217(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1218(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate855(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate856(.a(gate11inter0), .b(s_44), .O(gate11inter1));
  and2  gate857(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate858(.a(s_44), .O(gate11inter3));
  inv1  gate859(.a(s_45), .O(gate11inter4));
  nand2 gate860(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate861(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate862(.a(G5), .O(gate11inter7));
  inv1  gate863(.a(G6), .O(gate11inter8));
  nand2 gate864(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate865(.a(s_45), .b(gate11inter3), .O(gate11inter10));
  nor2  gate866(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate867(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate868(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate771(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate772(.a(gate17inter0), .b(s_32), .O(gate17inter1));
  and2  gate773(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate774(.a(s_32), .O(gate17inter3));
  inv1  gate775(.a(s_33), .O(gate17inter4));
  nand2 gate776(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate777(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate778(.a(G17), .O(gate17inter7));
  inv1  gate779(.a(G18), .O(gate17inter8));
  nand2 gate780(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate781(.a(s_33), .b(gate17inter3), .O(gate17inter10));
  nor2  gate782(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate783(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate784(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1275(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1276(.a(gate27inter0), .b(s_104), .O(gate27inter1));
  and2  gate1277(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1278(.a(s_104), .O(gate27inter3));
  inv1  gate1279(.a(s_105), .O(gate27inter4));
  nand2 gate1280(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1281(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1282(.a(G2), .O(gate27inter7));
  inv1  gate1283(.a(G6), .O(gate27inter8));
  nand2 gate1284(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1285(.a(s_105), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1286(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1287(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1288(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1135(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1136(.a(gate43inter0), .b(s_84), .O(gate43inter1));
  and2  gate1137(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1138(.a(s_84), .O(gate43inter3));
  inv1  gate1139(.a(s_85), .O(gate43inter4));
  nand2 gate1140(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1141(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1142(.a(G3), .O(gate43inter7));
  inv1  gate1143(.a(G269), .O(gate43inter8));
  nand2 gate1144(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1145(.a(s_85), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1146(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1147(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1148(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate995(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate996(.a(gate44inter0), .b(s_64), .O(gate44inter1));
  and2  gate997(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate998(.a(s_64), .O(gate44inter3));
  inv1  gate999(.a(s_65), .O(gate44inter4));
  nand2 gate1000(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1001(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1002(.a(G4), .O(gate44inter7));
  inv1  gate1003(.a(G269), .O(gate44inter8));
  nand2 gate1004(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1005(.a(s_65), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1006(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1007(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1008(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate673(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate674(.a(gate46inter0), .b(s_18), .O(gate46inter1));
  and2  gate675(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate676(.a(s_18), .O(gate46inter3));
  inv1  gate677(.a(s_19), .O(gate46inter4));
  nand2 gate678(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate679(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate680(.a(G6), .O(gate46inter7));
  inv1  gate681(.a(G272), .O(gate46inter8));
  nand2 gate682(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate683(.a(s_19), .b(gate46inter3), .O(gate46inter10));
  nor2  gate684(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate685(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate686(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate561(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate562(.a(gate50inter0), .b(s_2), .O(gate50inter1));
  and2  gate563(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate564(.a(s_2), .O(gate50inter3));
  inv1  gate565(.a(s_3), .O(gate50inter4));
  nand2 gate566(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate567(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate568(.a(G10), .O(gate50inter7));
  inv1  gate569(.a(G278), .O(gate50inter8));
  nand2 gate570(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate571(.a(s_3), .b(gate50inter3), .O(gate50inter10));
  nor2  gate572(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate573(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate574(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1107(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1108(.a(gate70inter0), .b(s_80), .O(gate70inter1));
  and2  gate1109(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1110(.a(s_80), .O(gate70inter3));
  inv1  gate1111(.a(s_81), .O(gate70inter4));
  nand2 gate1112(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1113(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1114(.a(G30), .O(gate70inter7));
  inv1  gate1115(.a(G308), .O(gate70inter8));
  nand2 gate1116(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1117(.a(s_81), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1118(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1119(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1120(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate813(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate814(.a(gate74inter0), .b(s_38), .O(gate74inter1));
  and2  gate815(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate816(.a(s_38), .O(gate74inter3));
  inv1  gate817(.a(s_39), .O(gate74inter4));
  nand2 gate818(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate819(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate820(.a(G5), .O(gate74inter7));
  inv1  gate821(.a(G314), .O(gate74inter8));
  nand2 gate822(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate823(.a(s_39), .b(gate74inter3), .O(gate74inter10));
  nor2  gate824(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate825(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate826(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate939(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate940(.a(gate78inter0), .b(s_56), .O(gate78inter1));
  and2  gate941(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate942(.a(s_56), .O(gate78inter3));
  inv1  gate943(.a(s_57), .O(gate78inter4));
  nand2 gate944(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate945(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate946(.a(G6), .O(gate78inter7));
  inv1  gate947(.a(G320), .O(gate78inter8));
  nand2 gate948(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate949(.a(s_57), .b(gate78inter3), .O(gate78inter10));
  nor2  gate950(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate951(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate952(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1233(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1234(.a(gate79inter0), .b(s_98), .O(gate79inter1));
  and2  gate1235(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1236(.a(s_98), .O(gate79inter3));
  inv1  gate1237(.a(s_99), .O(gate79inter4));
  nand2 gate1238(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1239(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1240(.a(G10), .O(gate79inter7));
  inv1  gate1241(.a(G323), .O(gate79inter8));
  nand2 gate1242(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1243(.a(s_99), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1244(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1245(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1246(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate687(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate688(.a(gate87inter0), .b(s_20), .O(gate87inter1));
  and2  gate689(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate690(.a(s_20), .O(gate87inter3));
  inv1  gate691(.a(s_21), .O(gate87inter4));
  nand2 gate692(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate693(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate694(.a(G12), .O(gate87inter7));
  inv1  gate695(.a(G335), .O(gate87inter8));
  nand2 gate696(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate697(.a(s_21), .b(gate87inter3), .O(gate87inter10));
  nor2  gate698(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate699(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate700(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1121(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1122(.a(gate89inter0), .b(s_82), .O(gate89inter1));
  and2  gate1123(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1124(.a(s_82), .O(gate89inter3));
  inv1  gate1125(.a(s_83), .O(gate89inter4));
  nand2 gate1126(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1127(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1128(.a(G17), .O(gate89inter7));
  inv1  gate1129(.a(G338), .O(gate89inter8));
  nand2 gate1130(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1131(.a(s_83), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1132(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1133(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1134(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate785(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate786(.a(gate98inter0), .b(s_34), .O(gate98inter1));
  and2  gate787(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate788(.a(s_34), .O(gate98inter3));
  inv1  gate789(.a(s_35), .O(gate98inter4));
  nand2 gate790(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate791(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate792(.a(G23), .O(gate98inter7));
  inv1  gate793(.a(G350), .O(gate98inter8));
  nand2 gate794(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate795(.a(s_35), .b(gate98inter3), .O(gate98inter10));
  nor2  gate796(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate797(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate798(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate617(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate618(.a(gate99inter0), .b(s_10), .O(gate99inter1));
  and2  gate619(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate620(.a(s_10), .O(gate99inter3));
  inv1  gate621(.a(s_11), .O(gate99inter4));
  nand2 gate622(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate623(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate624(.a(G27), .O(gate99inter7));
  inv1  gate625(.a(G353), .O(gate99inter8));
  nand2 gate626(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate627(.a(s_11), .b(gate99inter3), .O(gate99inter10));
  nor2  gate628(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate629(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate630(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1065(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1066(.a(gate117inter0), .b(s_74), .O(gate117inter1));
  and2  gate1067(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1068(.a(s_74), .O(gate117inter3));
  inv1  gate1069(.a(s_75), .O(gate117inter4));
  nand2 gate1070(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1071(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1072(.a(G386), .O(gate117inter7));
  inv1  gate1073(.a(G387), .O(gate117inter8));
  nand2 gate1074(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1075(.a(s_75), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1076(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1077(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1078(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1163(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1164(.a(gate127inter0), .b(s_88), .O(gate127inter1));
  and2  gate1165(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1166(.a(s_88), .O(gate127inter3));
  inv1  gate1167(.a(s_89), .O(gate127inter4));
  nand2 gate1168(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1169(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1170(.a(G406), .O(gate127inter7));
  inv1  gate1171(.a(G407), .O(gate127inter8));
  nand2 gate1172(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1173(.a(s_89), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1174(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1175(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1176(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1093(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1094(.a(gate137inter0), .b(s_78), .O(gate137inter1));
  and2  gate1095(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1096(.a(s_78), .O(gate137inter3));
  inv1  gate1097(.a(s_79), .O(gate137inter4));
  nand2 gate1098(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1099(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1100(.a(G426), .O(gate137inter7));
  inv1  gate1101(.a(G429), .O(gate137inter8));
  nand2 gate1102(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1103(.a(s_79), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1104(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1105(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1106(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1247(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1248(.a(gate141inter0), .b(s_100), .O(gate141inter1));
  and2  gate1249(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1250(.a(s_100), .O(gate141inter3));
  inv1  gate1251(.a(s_101), .O(gate141inter4));
  nand2 gate1252(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1253(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1254(.a(G450), .O(gate141inter7));
  inv1  gate1255(.a(G453), .O(gate141inter8));
  nand2 gate1256(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1257(.a(s_101), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1258(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1259(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1260(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate575(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate576(.a(gate153inter0), .b(s_4), .O(gate153inter1));
  and2  gate577(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate578(.a(s_4), .O(gate153inter3));
  inv1  gate579(.a(s_5), .O(gate153inter4));
  nand2 gate580(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate581(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate582(.a(G426), .O(gate153inter7));
  inv1  gate583(.a(G522), .O(gate153inter8));
  nand2 gate584(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate585(.a(s_5), .b(gate153inter3), .O(gate153inter10));
  nor2  gate586(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate587(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate588(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate743(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate744(.a(gate155inter0), .b(s_28), .O(gate155inter1));
  and2  gate745(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate746(.a(s_28), .O(gate155inter3));
  inv1  gate747(.a(s_29), .O(gate155inter4));
  nand2 gate748(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate749(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate750(.a(G432), .O(gate155inter7));
  inv1  gate751(.a(G525), .O(gate155inter8));
  nand2 gate752(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate753(.a(s_29), .b(gate155inter3), .O(gate155inter10));
  nor2  gate754(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate755(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate756(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1037(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1038(.a(gate166inter0), .b(s_70), .O(gate166inter1));
  and2  gate1039(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1040(.a(s_70), .O(gate166inter3));
  inv1  gate1041(.a(s_71), .O(gate166inter4));
  nand2 gate1042(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1043(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1044(.a(G465), .O(gate166inter7));
  inv1  gate1045(.a(G540), .O(gate166inter8));
  nand2 gate1046(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1047(.a(s_71), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1048(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1049(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1050(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1289(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1290(.a(gate168inter0), .b(s_106), .O(gate168inter1));
  and2  gate1291(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1292(.a(s_106), .O(gate168inter3));
  inv1  gate1293(.a(s_107), .O(gate168inter4));
  nand2 gate1294(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1295(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1296(.a(G471), .O(gate168inter7));
  inv1  gate1297(.a(G543), .O(gate168inter8));
  nand2 gate1298(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1299(.a(s_107), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1300(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1301(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1302(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate911(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate912(.a(gate170inter0), .b(s_52), .O(gate170inter1));
  and2  gate913(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate914(.a(s_52), .O(gate170inter3));
  inv1  gate915(.a(s_53), .O(gate170inter4));
  nand2 gate916(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate917(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate918(.a(G477), .O(gate170inter7));
  inv1  gate919(.a(G546), .O(gate170inter8));
  nand2 gate920(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate921(.a(s_53), .b(gate170inter3), .O(gate170inter10));
  nor2  gate922(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate923(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate924(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1261(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1262(.a(gate178inter0), .b(s_102), .O(gate178inter1));
  and2  gate1263(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1264(.a(s_102), .O(gate178inter3));
  inv1  gate1265(.a(s_103), .O(gate178inter4));
  nand2 gate1266(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1267(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1268(.a(G501), .O(gate178inter7));
  inv1  gate1269(.a(G558), .O(gate178inter8));
  nand2 gate1270(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1271(.a(s_103), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1272(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1273(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1274(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate953(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate954(.a(gate180inter0), .b(s_58), .O(gate180inter1));
  and2  gate955(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate956(.a(s_58), .O(gate180inter3));
  inv1  gate957(.a(s_59), .O(gate180inter4));
  nand2 gate958(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate959(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate960(.a(G507), .O(gate180inter7));
  inv1  gate961(.a(G561), .O(gate180inter8));
  nand2 gate962(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate963(.a(s_59), .b(gate180inter3), .O(gate180inter10));
  nor2  gate964(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate965(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate966(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate757(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate758(.a(gate188inter0), .b(s_30), .O(gate188inter1));
  and2  gate759(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate760(.a(s_30), .O(gate188inter3));
  inv1  gate761(.a(s_31), .O(gate188inter4));
  nand2 gate762(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate763(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate764(.a(G576), .O(gate188inter7));
  inv1  gate765(.a(G577), .O(gate188inter8));
  nand2 gate766(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate767(.a(s_31), .b(gate188inter3), .O(gate188inter10));
  nor2  gate768(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate769(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate770(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate869(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate870(.a(gate191inter0), .b(s_46), .O(gate191inter1));
  and2  gate871(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate872(.a(s_46), .O(gate191inter3));
  inv1  gate873(.a(s_47), .O(gate191inter4));
  nand2 gate874(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate875(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate876(.a(G582), .O(gate191inter7));
  inv1  gate877(.a(G583), .O(gate191inter8));
  nand2 gate878(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate879(.a(s_47), .b(gate191inter3), .O(gate191inter10));
  nor2  gate880(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate881(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate882(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate659(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate660(.a(gate202inter0), .b(s_16), .O(gate202inter1));
  and2  gate661(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate662(.a(s_16), .O(gate202inter3));
  inv1  gate663(.a(s_17), .O(gate202inter4));
  nand2 gate664(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate665(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate666(.a(G612), .O(gate202inter7));
  inv1  gate667(.a(G617), .O(gate202inter8));
  nand2 gate668(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate669(.a(s_17), .b(gate202inter3), .O(gate202inter10));
  nor2  gate670(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate671(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate672(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate701(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate702(.a(gate205inter0), .b(s_22), .O(gate205inter1));
  and2  gate703(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate704(.a(s_22), .O(gate205inter3));
  inv1  gate705(.a(s_23), .O(gate205inter4));
  nand2 gate706(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate707(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate708(.a(G622), .O(gate205inter7));
  inv1  gate709(.a(G627), .O(gate205inter8));
  nand2 gate710(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate711(.a(s_23), .b(gate205inter3), .O(gate205inter10));
  nor2  gate712(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate713(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate714(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1051(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1052(.a(gate217inter0), .b(s_72), .O(gate217inter1));
  and2  gate1053(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1054(.a(s_72), .O(gate217inter3));
  inv1  gate1055(.a(s_73), .O(gate217inter4));
  nand2 gate1056(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1057(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1058(.a(G622), .O(gate217inter7));
  inv1  gate1059(.a(G678), .O(gate217inter8));
  nand2 gate1060(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1061(.a(s_73), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1062(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1063(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1064(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate589(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate590(.a(gate226inter0), .b(s_6), .O(gate226inter1));
  and2  gate591(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate592(.a(s_6), .O(gate226inter3));
  inv1  gate593(.a(s_7), .O(gate226inter4));
  nand2 gate594(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate595(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate596(.a(G692), .O(gate226inter7));
  inv1  gate597(.a(G693), .O(gate226inter8));
  nand2 gate598(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate599(.a(s_7), .b(gate226inter3), .O(gate226inter10));
  nor2  gate600(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate601(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate602(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate631(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate632(.a(gate233inter0), .b(s_12), .O(gate233inter1));
  and2  gate633(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate634(.a(s_12), .O(gate233inter3));
  inv1  gate635(.a(s_13), .O(gate233inter4));
  nand2 gate636(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate637(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate638(.a(G242), .O(gate233inter7));
  inv1  gate639(.a(G718), .O(gate233inter8));
  nand2 gate640(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate641(.a(s_13), .b(gate233inter3), .O(gate233inter10));
  nor2  gate642(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate643(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate644(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1219(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1220(.a(gate254inter0), .b(s_96), .O(gate254inter1));
  and2  gate1221(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1222(.a(s_96), .O(gate254inter3));
  inv1  gate1223(.a(s_97), .O(gate254inter4));
  nand2 gate1224(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1225(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1226(.a(G712), .O(gate254inter7));
  inv1  gate1227(.a(G748), .O(gate254inter8));
  nand2 gate1228(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1229(.a(s_97), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1230(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1231(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1232(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate981(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate982(.a(gate258inter0), .b(s_62), .O(gate258inter1));
  and2  gate983(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate984(.a(s_62), .O(gate258inter3));
  inv1  gate985(.a(s_63), .O(gate258inter4));
  nand2 gate986(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate987(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate988(.a(G756), .O(gate258inter7));
  inv1  gate989(.a(G757), .O(gate258inter8));
  nand2 gate990(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate991(.a(s_63), .b(gate258inter3), .O(gate258inter10));
  nor2  gate992(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate993(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate994(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate799(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate800(.a(gate266inter0), .b(s_36), .O(gate266inter1));
  and2  gate801(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate802(.a(s_36), .O(gate266inter3));
  inv1  gate803(.a(s_37), .O(gate266inter4));
  nand2 gate804(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate805(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate806(.a(G645), .O(gate266inter7));
  inv1  gate807(.a(G773), .O(gate266inter8));
  nand2 gate808(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate809(.a(s_37), .b(gate266inter3), .O(gate266inter10));
  nor2  gate810(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate811(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate812(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate547(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate548(.a(gate279inter0), .b(s_0), .O(gate279inter1));
  and2  gate549(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate550(.a(s_0), .O(gate279inter3));
  inv1  gate551(.a(s_1), .O(gate279inter4));
  nand2 gate552(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate553(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate554(.a(G651), .O(gate279inter7));
  inv1  gate555(.a(G803), .O(gate279inter8));
  nand2 gate556(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate557(.a(s_1), .b(gate279inter3), .O(gate279inter10));
  nor2  gate558(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate559(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate560(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1191(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1192(.a(gate280inter0), .b(s_92), .O(gate280inter1));
  and2  gate1193(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1194(.a(s_92), .O(gate280inter3));
  inv1  gate1195(.a(s_93), .O(gate280inter4));
  nand2 gate1196(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1197(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1198(.a(G779), .O(gate280inter7));
  inv1  gate1199(.a(G803), .O(gate280inter8));
  nand2 gate1200(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1201(.a(s_93), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1202(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1203(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1204(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate827(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate828(.a(gate285inter0), .b(s_40), .O(gate285inter1));
  and2  gate829(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate830(.a(s_40), .O(gate285inter3));
  inv1  gate831(.a(s_41), .O(gate285inter4));
  nand2 gate832(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate833(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate834(.a(G660), .O(gate285inter7));
  inv1  gate835(.a(G812), .O(gate285inter8));
  nand2 gate836(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate837(.a(s_41), .b(gate285inter3), .O(gate285inter10));
  nor2  gate838(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate839(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate840(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate897(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate898(.a(gate290inter0), .b(s_50), .O(gate290inter1));
  and2  gate899(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate900(.a(s_50), .O(gate290inter3));
  inv1  gate901(.a(s_51), .O(gate290inter4));
  nand2 gate902(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate903(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate904(.a(G820), .O(gate290inter7));
  inv1  gate905(.a(G821), .O(gate290inter8));
  nand2 gate906(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate907(.a(s_51), .b(gate290inter3), .O(gate290inter10));
  nor2  gate908(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate909(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate910(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1177(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1178(.a(gate388inter0), .b(s_90), .O(gate388inter1));
  and2  gate1179(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1180(.a(s_90), .O(gate388inter3));
  inv1  gate1181(.a(s_91), .O(gate388inter4));
  nand2 gate1182(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1183(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1184(.a(G2), .O(gate388inter7));
  inv1  gate1185(.a(G1039), .O(gate388inter8));
  nand2 gate1186(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1187(.a(s_91), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1188(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1189(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1190(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate925(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate926(.a(gate394inter0), .b(s_54), .O(gate394inter1));
  and2  gate927(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate928(.a(s_54), .O(gate394inter3));
  inv1  gate929(.a(s_55), .O(gate394inter4));
  nand2 gate930(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate931(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate932(.a(G8), .O(gate394inter7));
  inv1  gate933(.a(G1057), .O(gate394inter8));
  nand2 gate934(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate935(.a(s_55), .b(gate394inter3), .O(gate394inter10));
  nor2  gate936(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate937(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate938(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate645(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate646(.a(gate395inter0), .b(s_14), .O(gate395inter1));
  and2  gate647(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate648(.a(s_14), .O(gate395inter3));
  inv1  gate649(.a(s_15), .O(gate395inter4));
  nand2 gate650(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate651(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate652(.a(G9), .O(gate395inter7));
  inv1  gate653(.a(G1060), .O(gate395inter8));
  nand2 gate654(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate655(.a(s_15), .b(gate395inter3), .O(gate395inter10));
  nor2  gate656(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate657(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate658(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate967(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate968(.a(gate435inter0), .b(s_60), .O(gate435inter1));
  and2  gate969(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate970(.a(s_60), .O(gate435inter3));
  inv1  gate971(.a(s_61), .O(gate435inter4));
  nand2 gate972(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate973(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate974(.a(G9), .O(gate435inter7));
  inv1  gate975(.a(G1156), .O(gate435inter8));
  nand2 gate976(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate977(.a(s_61), .b(gate435inter3), .O(gate435inter10));
  nor2  gate978(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate979(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate980(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate715(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate716(.a(gate436inter0), .b(s_24), .O(gate436inter1));
  and2  gate717(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate718(.a(s_24), .O(gate436inter3));
  inv1  gate719(.a(s_25), .O(gate436inter4));
  nand2 gate720(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate721(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate722(.a(G1060), .O(gate436inter7));
  inv1  gate723(.a(G1156), .O(gate436inter8));
  nand2 gate724(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate725(.a(s_25), .b(gate436inter3), .O(gate436inter10));
  nor2  gate726(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate727(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate728(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate729(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate730(.a(gate440inter0), .b(s_26), .O(gate440inter1));
  and2  gate731(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate732(.a(s_26), .O(gate440inter3));
  inv1  gate733(.a(s_27), .O(gate440inter4));
  nand2 gate734(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate735(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate736(.a(G1066), .O(gate440inter7));
  inv1  gate737(.a(G1162), .O(gate440inter8));
  nand2 gate738(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate739(.a(s_27), .b(gate440inter3), .O(gate440inter10));
  nor2  gate740(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate741(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate742(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1317(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1318(.a(gate442inter0), .b(s_110), .O(gate442inter1));
  and2  gate1319(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1320(.a(s_110), .O(gate442inter3));
  inv1  gate1321(.a(s_111), .O(gate442inter4));
  nand2 gate1322(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1323(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1324(.a(G1069), .O(gate442inter7));
  inv1  gate1325(.a(G1165), .O(gate442inter8));
  nand2 gate1326(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1327(.a(s_111), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1328(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1329(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1330(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1009(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1010(.a(gate456inter0), .b(s_66), .O(gate456inter1));
  and2  gate1011(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1012(.a(s_66), .O(gate456inter3));
  inv1  gate1013(.a(s_67), .O(gate456inter4));
  nand2 gate1014(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1015(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1016(.a(G1090), .O(gate456inter7));
  inv1  gate1017(.a(G1186), .O(gate456inter8));
  nand2 gate1018(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1019(.a(s_67), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1020(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1021(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1022(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1079(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1080(.a(gate465inter0), .b(s_76), .O(gate465inter1));
  and2  gate1081(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1082(.a(s_76), .O(gate465inter3));
  inv1  gate1083(.a(s_77), .O(gate465inter4));
  nand2 gate1084(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1085(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1086(.a(G24), .O(gate465inter7));
  inv1  gate1087(.a(G1201), .O(gate465inter8));
  nand2 gate1088(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1089(.a(s_77), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1090(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1091(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1092(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1303(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1304(.a(gate484inter0), .b(s_108), .O(gate484inter1));
  and2  gate1305(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1306(.a(s_108), .O(gate484inter3));
  inv1  gate1307(.a(s_109), .O(gate484inter4));
  nand2 gate1308(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1309(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1310(.a(G1230), .O(gate484inter7));
  inv1  gate1311(.a(G1231), .O(gate484inter8));
  nand2 gate1312(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1313(.a(s_109), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1314(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1315(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1316(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate603(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate604(.a(gate486inter0), .b(s_8), .O(gate486inter1));
  and2  gate605(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate606(.a(s_8), .O(gate486inter3));
  inv1  gate607(.a(s_9), .O(gate486inter4));
  nand2 gate608(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate609(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate610(.a(G1234), .O(gate486inter7));
  inv1  gate611(.a(G1235), .O(gate486inter8));
  nand2 gate612(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate613(.a(s_9), .b(gate486inter3), .O(gate486inter10));
  nor2  gate614(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate615(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate616(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate883(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate884(.a(gate503inter0), .b(s_48), .O(gate503inter1));
  and2  gate885(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate886(.a(s_48), .O(gate503inter3));
  inv1  gate887(.a(s_49), .O(gate503inter4));
  nand2 gate888(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate889(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate890(.a(G1268), .O(gate503inter7));
  inv1  gate891(.a(G1269), .O(gate503inter8));
  nand2 gate892(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate893(.a(s_49), .b(gate503inter3), .O(gate503inter10));
  nor2  gate894(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate895(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate896(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate841(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate842(.a(gate506inter0), .b(s_42), .O(gate506inter1));
  and2  gate843(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate844(.a(s_42), .O(gate506inter3));
  inv1  gate845(.a(s_43), .O(gate506inter4));
  nand2 gate846(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate847(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate848(.a(G1274), .O(gate506inter7));
  inv1  gate849(.a(G1275), .O(gate506inter8));
  nand2 gate850(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate851(.a(s_43), .b(gate506inter3), .O(gate506inter10));
  nor2  gate852(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate853(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate854(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1149(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1150(.a(gate508inter0), .b(s_86), .O(gate508inter1));
  and2  gate1151(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1152(.a(s_86), .O(gate508inter3));
  inv1  gate1153(.a(s_87), .O(gate508inter4));
  nand2 gate1154(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1155(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1156(.a(G1278), .O(gate508inter7));
  inv1  gate1157(.a(G1279), .O(gate508inter8));
  nand2 gate1158(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1159(.a(s_87), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1160(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1161(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1162(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1023(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1024(.a(gate511inter0), .b(s_68), .O(gate511inter1));
  and2  gate1025(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1026(.a(s_68), .O(gate511inter3));
  inv1  gate1027(.a(s_69), .O(gate511inter4));
  nand2 gate1028(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1029(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1030(.a(G1284), .O(gate511inter7));
  inv1  gate1031(.a(G1285), .O(gate511inter8));
  nand2 gate1032(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1033(.a(s_69), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1034(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1035(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1036(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule