module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate427(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate428(.a(gate24inter0), .b(s_38), .O(gate24inter1));
  and2  gate429(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate430(.a(s_38), .O(gate24inter3));
  inv1  gate431(.a(s_39), .O(gate24inter4));
  nand2 gate432(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate433(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate434(.a(N130), .O(gate24inter7));
  inv1  gate435(.a(N43), .O(gate24inter8));
  nand2 gate436(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate437(.a(s_39), .b(gate24inter3), .O(gate24inter10));
  nor2  gate438(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate439(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate440(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate385(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate386(.a(gate27inter0), .b(s_32), .O(gate27inter1));
  and2  gate387(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate388(.a(s_32), .O(gate27inter3));
  inv1  gate389(.a(s_33), .O(gate27inter4));
  nand2 gate390(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate391(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate392(.a(N142), .O(gate27inter7));
  inv1  gate393(.a(N82), .O(gate27inter8));
  nand2 gate394(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate395(.a(s_33), .b(gate27inter3), .O(gate27inter10));
  nor2  gate396(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate397(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate398(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate357(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate358(.a(gate29inter0), .b(s_28), .O(gate29inter1));
  and2  gate359(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate360(.a(s_28), .O(gate29inter3));
  inv1  gate361(.a(s_29), .O(gate29inter4));
  nand2 gate362(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate363(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate364(.a(N150), .O(gate29inter7));
  inv1  gate365(.a(N108), .O(gate29inter8));
  nand2 gate366(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate367(.a(s_29), .b(gate29inter3), .O(gate29inter10));
  nor2  gate368(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate369(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate370(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate273(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate274(.a(gate38inter0), .b(s_16), .O(gate38inter1));
  and2  gate275(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate276(.a(s_16), .O(gate38inter3));
  inv1  gate277(.a(s_17), .O(gate38inter4));
  nand2 gate278(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate279(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate280(.a(N73), .O(gate38inter7));
  inv1  gate281(.a(N139), .O(gate38inter8));
  nand2 gate282(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate283(.a(s_17), .b(gate38inter3), .O(gate38inter10));
  nor2  gate284(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate285(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate286(.a(gate38inter12), .b(gate38inter1), .O(N191));
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate175(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate176(.a(gate41inter0), .b(s_2), .O(gate41inter1));
  and2  gate177(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate178(.a(s_2), .O(gate41inter3));
  inv1  gate179(.a(s_3), .O(gate41inter4));
  nand2 gate180(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate181(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate182(.a(N92), .O(gate41inter7));
  inv1  gate183(.a(N143), .O(gate41inter8));
  nand2 gate184(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate185(.a(s_3), .b(gate41inter3), .O(gate41inter10));
  nor2  gate186(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate187(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate188(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate315(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate316(.a(gate50inter0), .b(s_22), .O(gate50inter1));
  and2  gate317(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate318(.a(s_22), .O(gate50inter3));
  inv1  gate319(.a(s_23), .O(gate50inter4));
  nand2 gate320(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate321(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate322(.a(N203), .O(gate50inter7));
  inv1  gate323(.a(N154), .O(gate50inter8));
  nand2 gate324(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate325(.a(s_23), .b(gate50inter3), .O(gate50inter10));
  nor2  gate326(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate327(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate328(.a(gate50inter12), .b(gate50inter1), .O(N224));
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate301(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate302(.a(gate57inter0), .b(s_20), .O(gate57inter1));
  and2  gate303(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate304(.a(s_20), .O(gate57inter3));
  inv1  gate305(.a(s_21), .O(gate57inter4));
  nand2 gate306(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate307(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate308(.a(N203), .O(gate57inter7));
  inv1  gate309(.a(N174), .O(gate57inter8));
  nand2 gate310(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate311(.a(s_21), .b(gate57inter3), .O(gate57inter10));
  nor2  gate312(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate313(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate314(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate441(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate442(.a(gate62inter0), .b(s_40), .O(gate62inter1));
  and2  gate443(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate444(.a(s_40), .O(gate62inter3));
  inv1  gate445(.a(s_41), .O(gate62inter4));
  nand2 gate446(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate447(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate448(.a(N213), .O(gate62inter7));
  inv1  gate449(.a(N37), .O(gate62inter8));
  nand2 gate450(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate451(.a(s_41), .b(gate62inter3), .O(gate62inter10));
  nor2  gate452(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate453(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate454(.a(gate62inter12), .b(gate62inter1), .O(N254));
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate413(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate414(.a(gate65inter0), .b(s_36), .O(gate65inter1));
  and2  gate415(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate416(.a(s_36), .O(gate65inter3));
  inv1  gate417(.a(s_37), .O(gate65inter4));
  nand2 gate418(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate419(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate420(.a(N213), .O(gate65inter7));
  inv1  gate421(.a(N76), .O(gate65inter8));
  nand2 gate422(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate423(.a(s_37), .b(gate65inter3), .O(gate65inter10));
  nor2  gate424(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate425(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate426(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );

  xor2  gate329(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate330(.a(gate67inter0), .b(s_24), .O(gate67inter1));
  and2  gate331(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate332(.a(s_24), .O(gate67inter3));
  inv1  gate333(.a(s_25), .O(gate67inter4));
  nand2 gate334(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate335(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate336(.a(N213), .O(gate67inter7));
  inv1  gate337(.a(N102), .O(gate67inter8));
  nand2 gate338(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate339(.a(s_25), .b(gate67inter3), .O(gate67inter10));
  nor2  gate340(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate341(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate342(.a(gate67inter12), .b(gate67inter1), .O(N259));
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );

  xor2  gate189(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate190(.a(gate81inter0), .b(s_4), .O(gate81inter1));
  and2  gate191(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate192(.a(s_4), .O(gate81inter3));
  inv1  gate193(.a(s_5), .O(gate81inter4));
  nand2 gate194(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate195(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate196(.a(N236), .O(gate81inter7));
  inv1  gate197(.a(N190), .O(gate81inter8));
  nand2 gate198(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate199(.a(s_5), .b(gate81inter3), .O(gate81inter10));
  nor2  gate200(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate201(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate202(.a(gate81inter12), .b(gate81inter1), .O(N291));
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );

  xor2  gate245(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate246(.a(gate100inter0), .b(s_12), .O(gate100inter1));
  and2  gate247(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate248(.a(s_12), .O(gate100inter3));
  inv1  gate249(.a(s_13), .O(gate100inter4));
  nand2 gate250(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate251(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate252(.a(N309), .O(gate100inter7));
  inv1  gate253(.a(N264), .O(gate100inter8));
  nand2 gate254(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate255(.a(s_13), .b(gate100inter3), .O(gate100inter10));
  nor2  gate256(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate257(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate258(.a(gate100inter12), .b(gate100inter1), .O(N331));
xor2 gate101( .a(N309), .b(N267), .O(N332) );

  xor2  gate259(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate260(.a(gate102inter0), .b(s_14), .O(gate102inter1));
  and2  gate261(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate262(.a(s_14), .O(gate102inter3));
  inv1  gate263(.a(s_15), .O(gate102inter4));
  nand2 gate264(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate265(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate266(.a(N309), .O(gate102inter7));
  inv1  gate267(.a(N270), .O(gate102inter8));
  nand2 gate268(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate269(.a(s_15), .b(gate102inter3), .O(gate102inter10));
  nor2  gate270(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate271(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate272(.a(gate102inter12), .b(gate102inter1), .O(N333));
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate203(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate204(.a(gate110inter0), .b(s_6), .O(gate110inter1));
  and2  gate205(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate206(.a(s_6), .O(gate110inter3));
  inv1  gate207(.a(s_7), .O(gate110inter4));
  nand2 gate208(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate209(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate210(.a(N309), .O(gate110inter7));
  inv1  gate211(.a(N282), .O(gate110inter8));
  nand2 gate212(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate213(.a(s_7), .b(gate110inter3), .O(gate110inter10));
  nor2  gate214(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate215(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate216(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );

  xor2  gate161(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate162(.a(gate112inter0), .b(s_0), .O(gate112inter1));
  and2  gate163(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate164(.a(s_0), .O(gate112inter3));
  inv1  gate165(.a(s_1), .O(gate112inter4));
  nand2 gate166(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate167(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate168(.a(N309), .O(gate112inter7));
  inv1  gate169(.a(N285), .O(gate112inter8));
  nand2 gate170(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate171(.a(s_1), .b(gate112inter3), .O(gate112inter10));
  nor2  gate172(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate173(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate174(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );

  xor2  gate399(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate400(.a(gate116inter0), .b(s_34), .O(gate116inter1));
  and2  gate401(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate402(.a(s_34), .O(gate116inter3));
  inv1  gate403(.a(s_35), .O(gate116inter4));
  nand2 gate404(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate405(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate406(.a(N319), .O(gate116inter7));
  inv1  gate407(.a(N112), .O(gate116inter8));
  nand2 gate408(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate409(.a(s_35), .b(gate116inter3), .O(gate116inter10));
  nor2  gate410(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate411(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate412(.a(gate116inter12), .b(gate116inter1), .O(N347));

  xor2  gate287(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate288(.a(gate117inter0), .b(s_18), .O(gate117inter1));
  and2  gate289(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate290(.a(s_18), .O(gate117inter3));
  inv1  gate291(.a(s_19), .O(gate117inter4));
  nand2 gate292(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate293(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate294(.a(N330), .O(gate117inter7));
  inv1  gate295(.a(N300), .O(gate117inter8));
  nand2 gate296(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate297(.a(s_19), .b(gate117inter3), .O(gate117inter10));
  nor2  gate298(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate299(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate300(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate343(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate344(.a(gate120inter0), .b(s_26), .O(gate120inter1));
  and2  gate345(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate346(.a(s_26), .O(gate120inter3));
  inv1  gate347(.a(s_27), .O(gate120inter4));
  nand2 gate348(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate349(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate350(.a(N333), .O(gate120inter7));
  inv1  gate351(.a(N303), .O(gate120inter8));
  nand2 gate352(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate353(.a(s_27), .b(gate120inter3), .O(gate120inter10));
  nor2  gate354(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate355(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate356(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate371(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate372(.a(gate135inter0), .b(s_30), .O(gate135inter1));
  and2  gate373(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate374(.a(s_30), .O(gate135inter3));
  inv1  gate375(.a(s_31), .O(gate135inter4));
  nand2 gate376(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate377(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate378(.a(N360), .O(gate135inter7));
  inv1  gate379(.a(N92), .O(gate135inter8));
  nand2 gate380(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate381(.a(s_31), .b(gate135inter3), .O(gate135inter10));
  nor2  gate382(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate383(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate384(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate231(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate232(.a(gate153inter0), .b(s_10), .O(gate153inter1));
  and2  gate233(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate234(.a(s_10), .O(gate153inter3));
  inv1  gate235(.a(s_11), .O(gate153inter4));
  nand2 gate236(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate237(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate238(.a(N415), .O(gate153inter7));
  inv1  gate239(.a(N416), .O(gate153inter8));
  nand2 gate240(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate241(.a(s_11), .b(gate153inter3), .O(gate153inter10));
  nor2  gate242(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate243(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate244(.a(gate153inter12), .b(gate153inter1), .O(N421));

  xor2  gate217(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate218(.a(gate154inter0), .b(s_8), .O(gate154inter1));
  and2  gate219(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate220(.a(s_8), .O(gate154inter3));
  inv1  gate221(.a(s_9), .O(gate154inter4));
  nand2 gate222(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate223(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate224(.a(N386), .O(gate154inter7));
  inv1  gate225(.a(N417), .O(gate154inter8));
  nand2 gate226(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate227(.a(s_9), .b(gate154inter3), .O(gate154inter10));
  nor2  gate228(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate229(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate230(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule