module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1121(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1122(.a(gate12inter0), .b(s_82), .O(gate12inter1));
  and2  gate1123(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1124(.a(s_82), .O(gate12inter3));
  inv1  gate1125(.a(s_83), .O(gate12inter4));
  nand2 gate1126(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1127(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1128(.a(G7), .O(gate12inter7));
  inv1  gate1129(.a(G8), .O(gate12inter8));
  nand2 gate1130(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1131(.a(s_83), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1132(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1133(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1134(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1555(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1556(.a(gate15inter0), .b(s_144), .O(gate15inter1));
  and2  gate1557(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1558(.a(s_144), .O(gate15inter3));
  inv1  gate1559(.a(s_145), .O(gate15inter4));
  nand2 gate1560(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1561(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1562(.a(G13), .O(gate15inter7));
  inv1  gate1563(.a(G14), .O(gate15inter8));
  nand2 gate1564(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1565(.a(s_145), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1566(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1567(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1568(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate785(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate786(.a(gate30inter0), .b(s_34), .O(gate30inter1));
  and2  gate787(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate788(.a(s_34), .O(gate30inter3));
  inv1  gate789(.a(s_35), .O(gate30inter4));
  nand2 gate790(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate791(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate792(.a(G11), .O(gate30inter7));
  inv1  gate793(.a(G15), .O(gate30inter8));
  nand2 gate794(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate795(.a(s_35), .b(gate30inter3), .O(gate30inter10));
  nor2  gate796(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate797(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate798(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate771(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate772(.a(gate32inter0), .b(s_32), .O(gate32inter1));
  and2  gate773(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate774(.a(s_32), .O(gate32inter3));
  inv1  gate775(.a(s_33), .O(gate32inter4));
  nand2 gate776(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate777(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate778(.a(G12), .O(gate32inter7));
  inv1  gate779(.a(G16), .O(gate32inter8));
  nand2 gate780(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate781(.a(s_33), .b(gate32inter3), .O(gate32inter10));
  nor2  gate782(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate783(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate784(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate631(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate632(.a(gate36inter0), .b(s_12), .O(gate36inter1));
  and2  gate633(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate634(.a(s_12), .O(gate36inter3));
  inv1  gate635(.a(s_13), .O(gate36inter4));
  nand2 gate636(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate637(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate638(.a(G26), .O(gate36inter7));
  inv1  gate639(.a(G30), .O(gate36inter8));
  nand2 gate640(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate641(.a(s_13), .b(gate36inter3), .O(gate36inter10));
  nor2  gate642(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate643(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate644(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1639(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1640(.a(gate37inter0), .b(s_156), .O(gate37inter1));
  and2  gate1641(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1642(.a(s_156), .O(gate37inter3));
  inv1  gate1643(.a(s_157), .O(gate37inter4));
  nand2 gate1644(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1645(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1646(.a(G19), .O(gate37inter7));
  inv1  gate1647(.a(G23), .O(gate37inter8));
  nand2 gate1648(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1649(.a(s_157), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1650(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1651(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1652(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate715(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate716(.a(gate39inter0), .b(s_24), .O(gate39inter1));
  and2  gate717(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate718(.a(s_24), .O(gate39inter3));
  inv1  gate719(.a(s_25), .O(gate39inter4));
  nand2 gate720(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate721(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate722(.a(G20), .O(gate39inter7));
  inv1  gate723(.a(G24), .O(gate39inter8));
  nand2 gate724(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate725(.a(s_25), .b(gate39inter3), .O(gate39inter10));
  nor2  gate726(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate727(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate728(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate813(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate814(.a(gate50inter0), .b(s_38), .O(gate50inter1));
  and2  gate815(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate816(.a(s_38), .O(gate50inter3));
  inv1  gate817(.a(s_39), .O(gate50inter4));
  nand2 gate818(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate819(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate820(.a(G10), .O(gate50inter7));
  inv1  gate821(.a(G278), .O(gate50inter8));
  nand2 gate822(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate823(.a(s_39), .b(gate50inter3), .O(gate50inter10));
  nor2  gate824(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate825(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate826(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1331(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1332(.a(gate58inter0), .b(s_112), .O(gate58inter1));
  and2  gate1333(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1334(.a(s_112), .O(gate58inter3));
  inv1  gate1335(.a(s_113), .O(gate58inter4));
  nand2 gate1336(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1337(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1338(.a(G18), .O(gate58inter7));
  inv1  gate1339(.a(G290), .O(gate58inter8));
  nand2 gate1340(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1341(.a(s_113), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1342(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1343(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1344(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate547(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate548(.a(gate63inter0), .b(s_0), .O(gate63inter1));
  and2  gate549(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate550(.a(s_0), .O(gate63inter3));
  inv1  gate551(.a(s_1), .O(gate63inter4));
  nand2 gate552(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate553(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate554(.a(G23), .O(gate63inter7));
  inv1  gate555(.a(G299), .O(gate63inter8));
  nand2 gate556(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate557(.a(s_1), .b(gate63inter3), .O(gate63inter10));
  nor2  gate558(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate559(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate560(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1317(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1318(.a(gate64inter0), .b(s_110), .O(gate64inter1));
  and2  gate1319(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1320(.a(s_110), .O(gate64inter3));
  inv1  gate1321(.a(s_111), .O(gate64inter4));
  nand2 gate1322(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1323(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1324(.a(G24), .O(gate64inter7));
  inv1  gate1325(.a(G299), .O(gate64inter8));
  nand2 gate1326(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1327(.a(s_111), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1328(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1329(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1330(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1009(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1010(.a(gate85inter0), .b(s_66), .O(gate85inter1));
  and2  gate1011(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1012(.a(s_66), .O(gate85inter3));
  inv1  gate1013(.a(s_67), .O(gate85inter4));
  nand2 gate1014(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1015(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1016(.a(G4), .O(gate85inter7));
  inv1  gate1017(.a(G332), .O(gate85inter8));
  nand2 gate1018(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1019(.a(s_67), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1020(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1021(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1022(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate911(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate912(.a(gate90inter0), .b(s_52), .O(gate90inter1));
  and2  gate913(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate914(.a(s_52), .O(gate90inter3));
  inv1  gate915(.a(s_53), .O(gate90inter4));
  nand2 gate916(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate917(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate918(.a(G21), .O(gate90inter7));
  inv1  gate919(.a(G338), .O(gate90inter8));
  nand2 gate920(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate921(.a(s_53), .b(gate90inter3), .O(gate90inter10));
  nor2  gate922(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate923(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate924(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate617(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate618(.a(gate91inter0), .b(s_10), .O(gate91inter1));
  and2  gate619(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate620(.a(s_10), .O(gate91inter3));
  inv1  gate621(.a(s_11), .O(gate91inter4));
  nand2 gate622(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate623(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate624(.a(G25), .O(gate91inter7));
  inv1  gate625(.a(G341), .O(gate91inter8));
  nand2 gate626(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate627(.a(s_11), .b(gate91inter3), .O(gate91inter10));
  nor2  gate628(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate629(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate630(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1667(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1668(.a(gate100inter0), .b(s_160), .O(gate100inter1));
  and2  gate1669(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1670(.a(s_160), .O(gate100inter3));
  inv1  gate1671(.a(s_161), .O(gate100inter4));
  nand2 gate1672(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1673(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1674(.a(G31), .O(gate100inter7));
  inv1  gate1675(.a(G353), .O(gate100inter8));
  nand2 gate1676(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1677(.a(s_161), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1678(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1679(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1680(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1653(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1654(.a(gate104inter0), .b(s_158), .O(gate104inter1));
  and2  gate1655(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1656(.a(s_158), .O(gate104inter3));
  inv1  gate1657(.a(s_159), .O(gate104inter4));
  nand2 gate1658(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1659(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1660(.a(G32), .O(gate104inter7));
  inv1  gate1661(.a(G359), .O(gate104inter8));
  nand2 gate1662(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1663(.a(s_159), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1664(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1665(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1666(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate897(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate898(.a(gate106inter0), .b(s_50), .O(gate106inter1));
  and2  gate899(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate900(.a(s_50), .O(gate106inter3));
  inv1  gate901(.a(s_51), .O(gate106inter4));
  nand2 gate902(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate903(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate904(.a(G364), .O(gate106inter7));
  inv1  gate905(.a(G365), .O(gate106inter8));
  nand2 gate906(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate907(.a(s_51), .b(gate106inter3), .O(gate106inter10));
  nor2  gate908(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate909(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate910(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1401(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1402(.a(gate108inter0), .b(s_122), .O(gate108inter1));
  and2  gate1403(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1404(.a(s_122), .O(gate108inter3));
  inv1  gate1405(.a(s_123), .O(gate108inter4));
  nand2 gate1406(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1407(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1408(.a(G368), .O(gate108inter7));
  inv1  gate1409(.a(G369), .O(gate108inter8));
  nand2 gate1410(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1411(.a(s_123), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1412(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1413(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1414(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1135(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1136(.a(gate112inter0), .b(s_84), .O(gate112inter1));
  and2  gate1137(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1138(.a(s_84), .O(gate112inter3));
  inv1  gate1139(.a(s_85), .O(gate112inter4));
  nand2 gate1140(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1141(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1142(.a(G376), .O(gate112inter7));
  inv1  gate1143(.a(G377), .O(gate112inter8));
  nand2 gate1144(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1145(.a(s_85), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1146(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1147(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1148(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1149(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1150(.a(gate113inter0), .b(s_86), .O(gate113inter1));
  and2  gate1151(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1152(.a(s_86), .O(gate113inter3));
  inv1  gate1153(.a(s_87), .O(gate113inter4));
  nand2 gate1154(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1155(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1156(.a(G378), .O(gate113inter7));
  inv1  gate1157(.a(G379), .O(gate113inter8));
  nand2 gate1158(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1159(.a(s_87), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1160(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1161(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1162(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate827(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate828(.a(gate115inter0), .b(s_40), .O(gate115inter1));
  and2  gate829(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate830(.a(s_40), .O(gate115inter3));
  inv1  gate831(.a(s_41), .O(gate115inter4));
  nand2 gate832(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate833(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate834(.a(G382), .O(gate115inter7));
  inv1  gate835(.a(G383), .O(gate115inter8));
  nand2 gate836(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate837(.a(s_41), .b(gate115inter3), .O(gate115inter10));
  nor2  gate838(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate839(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate840(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1429(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1430(.a(gate117inter0), .b(s_126), .O(gate117inter1));
  and2  gate1431(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1432(.a(s_126), .O(gate117inter3));
  inv1  gate1433(.a(s_127), .O(gate117inter4));
  nand2 gate1434(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1435(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1436(.a(G386), .O(gate117inter7));
  inv1  gate1437(.a(G387), .O(gate117inter8));
  nand2 gate1438(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1439(.a(s_127), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1440(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1441(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1442(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1275(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1276(.a(gate128inter0), .b(s_104), .O(gate128inter1));
  and2  gate1277(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1278(.a(s_104), .O(gate128inter3));
  inv1  gate1279(.a(s_105), .O(gate128inter4));
  nand2 gate1280(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1281(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1282(.a(G408), .O(gate128inter7));
  inv1  gate1283(.a(G409), .O(gate128inter8));
  nand2 gate1284(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1285(.a(s_105), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1286(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1287(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1288(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1499(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1500(.a(gate132inter0), .b(s_136), .O(gate132inter1));
  and2  gate1501(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1502(.a(s_136), .O(gate132inter3));
  inv1  gate1503(.a(s_137), .O(gate132inter4));
  nand2 gate1504(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1505(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1506(.a(G416), .O(gate132inter7));
  inv1  gate1507(.a(G417), .O(gate132inter8));
  nand2 gate1508(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1509(.a(s_137), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1510(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1511(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1512(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1303(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1304(.a(gate133inter0), .b(s_108), .O(gate133inter1));
  and2  gate1305(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1306(.a(s_108), .O(gate133inter3));
  inv1  gate1307(.a(s_109), .O(gate133inter4));
  nand2 gate1308(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1309(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1310(.a(G418), .O(gate133inter7));
  inv1  gate1311(.a(G419), .O(gate133inter8));
  nand2 gate1312(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1313(.a(s_109), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1314(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1315(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1316(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate673(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate674(.a(gate136inter0), .b(s_18), .O(gate136inter1));
  and2  gate675(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate676(.a(s_18), .O(gate136inter3));
  inv1  gate677(.a(s_19), .O(gate136inter4));
  nand2 gate678(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate679(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate680(.a(G424), .O(gate136inter7));
  inv1  gate681(.a(G425), .O(gate136inter8));
  nand2 gate682(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate683(.a(s_19), .b(gate136inter3), .O(gate136inter10));
  nor2  gate684(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate685(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate686(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1247(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1248(.a(gate137inter0), .b(s_100), .O(gate137inter1));
  and2  gate1249(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1250(.a(s_100), .O(gate137inter3));
  inv1  gate1251(.a(s_101), .O(gate137inter4));
  nand2 gate1252(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1253(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1254(.a(G426), .O(gate137inter7));
  inv1  gate1255(.a(G429), .O(gate137inter8));
  nand2 gate1256(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1257(.a(s_101), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1258(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1259(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1260(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate701(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate702(.a(gate138inter0), .b(s_22), .O(gate138inter1));
  and2  gate703(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate704(.a(s_22), .O(gate138inter3));
  inv1  gate705(.a(s_23), .O(gate138inter4));
  nand2 gate706(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate707(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate708(.a(G432), .O(gate138inter7));
  inv1  gate709(.a(G435), .O(gate138inter8));
  nand2 gate710(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate711(.a(s_23), .b(gate138inter3), .O(gate138inter10));
  nor2  gate712(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate713(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate714(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1163(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1164(.a(gate139inter0), .b(s_88), .O(gate139inter1));
  and2  gate1165(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1166(.a(s_88), .O(gate139inter3));
  inv1  gate1167(.a(s_89), .O(gate139inter4));
  nand2 gate1168(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1169(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1170(.a(G438), .O(gate139inter7));
  inv1  gate1171(.a(G441), .O(gate139inter8));
  nand2 gate1172(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1173(.a(s_89), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1174(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1175(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1176(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate561(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate562(.a(gate143inter0), .b(s_2), .O(gate143inter1));
  and2  gate563(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate564(.a(s_2), .O(gate143inter3));
  inv1  gate565(.a(s_3), .O(gate143inter4));
  nand2 gate566(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate567(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate568(.a(G462), .O(gate143inter7));
  inv1  gate569(.a(G465), .O(gate143inter8));
  nand2 gate570(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate571(.a(s_3), .b(gate143inter3), .O(gate143inter10));
  nor2  gate572(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate573(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate574(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate855(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate856(.a(gate144inter0), .b(s_44), .O(gate144inter1));
  and2  gate857(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate858(.a(s_44), .O(gate144inter3));
  inv1  gate859(.a(s_45), .O(gate144inter4));
  nand2 gate860(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate861(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate862(.a(G468), .O(gate144inter7));
  inv1  gate863(.a(G471), .O(gate144inter8));
  nand2 gate864(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate865(.a(s_45), .b(gate144inter3), .O(gate144inter10));
  nor2  gate866(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate867(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate868(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate687(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate688(.a(gate152inter0), .b(s_20), .O(gate152inter1));
  and2  gate689(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate690(.a(s_20), .O(gate152inter3));
  inv1  gate691(.a(s_21), .O(gate152inter4));
  nand2 gate692(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate693(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate694(.a(G516), .O(gate152inter7));
  inv1  gate695(.a(G519), .O(gate152inter8));
  nand2 gate696(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate697(.a(s_21), .b(gate152inter3), .O(gate152inter10));
  nor2  gate698(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate699(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate700(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate603(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate604(.a(gate155inter0), .b(s_8), .O(gate155inter1));
  and2  gate605(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate606(.a(s_8), .O(gate155inter3));
  inv1  gate607(.a(s_9), .O(gate155inter4));
  nand2 gate608(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate609(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate610(.a(G432), .O(gate155inter7));
  inv1  gate611(.a(G525), .O(gate155inter8));
  nand2 gate612(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate613(.a(s_9), .b(gate155inter3), .O(gate155inter10));
  nor2  gate614(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate615(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate616(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate925(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate926(.a(gate156inter0), .b(s_54), .O(gate156inter1));
  and2  gate927(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate928(.a(s_54), .O(gate156inter3));
  inv1  gate929(.a(s_55), .O(gate156inter4));
  nand2 gate930(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate931(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate932(.a(G435), .O(gate156inter7));
  inv1  gate933(.a(G525), .O(gate156inter8));
  nand2 gate934(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate935(.a(s_55), .b(gate156inter3), .O(gate156inter10));
  nor2  gate936(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate937(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate938(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1611(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1612(.a(gate164inter0), .b(s_152), .O(gate164inter1));
  and2  gate1613(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1614(.a(s_152), .O(gate164inter3));
  inv1  gate1615(.a(s_153), .O(gate164inter4));
  nand2 gate1616(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1617(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1618(.a(G459), .O(gate164inter7));
  inv1  gate1619(.a(G537), .O(gate164inter8));
  nand2 gate1620(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1621(.a(s_153), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1622(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1623(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1624(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate1233(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1234(.a(gate165inter0), .b(s_98), .O(gate165inter1));
  and2  gate1235(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1236(.a(s_98), .O(gate165inter3));
  inv1  gate1237(.a(s_99), .O(gate165inter4));
  nand2 gate1238(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1239(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1240(.a(G462), .O(gate165inter7));
  inv1  gate1241(.a(G540), .O(gate165inter8));
  nand2 gate1242(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1243(.a(s_99), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1244(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1245(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1246(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1051(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1052(.a(gate166inter0), .b(s_72), .O(gate166inter1));
  and2  gate1053(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1054(.a(s_72), .O(gate166inter3));
  inv1  gate1055(.a(s_73), .O(gate166inter4));
  nand2 gate1056(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1057(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1058(.a(G465), .O(gate166inter7));
  inv1  gate1059(.a(G540), .O(gate166inter8));
  nand2 gate1060(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1061(.a(s_73), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1062(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1063(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1064(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1037(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1038(.a(gate170inter0), .b(s_70), .O(gate170inter1));
  and2  gate1039(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1040(.a(s_70), .O(gate170inter3));
  inv1  gate1041(.a(s_71), .O(gate170inter4));
  nand2 gate1042(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1043(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1044(.a(G477), .O(gate170inter7));
  inv1  gate1045(.a(G546), .O(gate170inter8));
  nand2 gate1046(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1047(.a(s_71), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1048(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1049(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1050(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate841(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate842(.a(gate173inter0), .b(s_42), .O(gate173inter1));
  and2  gate843(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate844(.a(s_42), .O(gate173inter3));
  inv1  gate845(.a(s_43), .O(gate173inter4));
  nand2 gate846(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate847(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate848(.a(G486), .O(gate173inter7));
  inv1  gate849(.a(G552), .O(gate173inter8));
  nand2 gate850(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate851(.a(s_43), .b(gate173inter3), .O(gate173inter10));
  nor2  gate852(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate853(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate854(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate967(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate968(.a(gate174inter0), .b(s_60), .O(gate174inter1));
  and2  gate969(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate970(.a(s_60), .O(gate174inter3));
  inv1  gate971(.a(s_61), .O(gate174inter4));
  nand2 gate972(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate973(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate974(.a(G489), .O(gate174inter7));
  inv1  gate975(.a(G552), .O(gate174inter8));
  nand2 gate976(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate977(.a(s_61), .b(gate174inter3), .O(gate174inter10));
  nor2  gate978(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate979(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate980(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1177(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1178(.a(gate175inter0), .b(s_90), .O(gate175inter1));
  and2  gate1179(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1180(.a(s_90), .O(gate175inter3));
  inv1  gate1181(.a(s_91), .O(gate175inter4));
  nand2 gate1182(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1183(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1184(.a(G492), .O(gate175inter7));
  inv1  gate1185(.a(G555), .O(gate175inter8));
  nand2 gate1186(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1187(.a(s_91), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1188(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1189(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1190(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate757(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate758(.a(gate188inter0), .b(s_30), .O(gate188inter1));
  and2  gate759(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate760(.a(s_30), .O(gate188inter3));
  inv1  gate761(.a(s_31), .O(gate188inter4));
  nand2 gate762(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate763(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate764(.a(G576), .O(gate188inter7));
  inv1  gate765(.a(G577), .O(gate188inter8));
  nand2 gate766(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate767(.a(s_31), .b(gate188inter3), .O(gate188inter10));
  nor2  gate768(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate769(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate770(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1345(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1346(.a(gate190inter0), .b(s_114), .O(gate190inter1));
  and2  gate1347(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1348(.a(s_114), .O(gate190inter3));
  inv1  gate1349(.a(s_115), .O(gate190inter4));
  nand2 gate1350(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1351(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1352(.a(G580), .O(gate190inter7));
  inv1  gate1353(.a(G581), .O(gate190inter8));
  nand2 gate1354(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1355(.a(s_115), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1356(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1357(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1358(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1107(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1108(.a(gate192inter0), .b(s_80), .O(gate192inter1));
  and2  gate1109(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1110(.a(s_80), .O(gate192inter3));
  inv1  gate1111(.a(s_81), .O(gate192inter4));
  nand2 gate1112(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1113(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1114(.a(G584), .O(gate192inter7));
  inv1  gate1115(.a(G585), .O(gate192inter8));
  nand2 gate1116(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1117(.a(s_81), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1118(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1119(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1120(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1205(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1206(.a(gate206inter0), .b(s_94), .O(gate206inter1));
  and2  gate1207(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1208(.a(s_94), .O(gate206inter3));
  inv1  gate1209(.a(s_95), .O(gate206inter4));
  nand2 gate1210(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1211(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1212(.a(G632), .O(gate206inter7));
  inv1  gate1213(.a(G637), .O(gate206inter8));
  nand2 gate1214(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1215(.a(s_95), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1216(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1217(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1218(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate743(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate744(.a(gate208inter0), .b(s_28), .O(gate208inter1));
  and2  gate745(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate746(.a(s_28), .O(gate208inter3));
  inv1  gate747(.a(s_29), .O(gate208inter4));
  nand2 gate748(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate749(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate750(.a(G627), .O(gate208inter7));
  inv1  gate751(.a(G637), .O(gate208inter8));
  nand2 gate752(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate753(.a(s_29), .b(gate208inter3), .O(gate208inter10));
  nor2  gate754(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate755(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate756(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1289(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1290(.a(gate209inter0), .b(s_106), .O(gate209inter1));
  and2  gate1291(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1292(.a(s_106), .O(gate209inter3));
  inv1  gate1293(.a(s_107), .O(gate209inter4));
  nand2 gate1294(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1295(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1296(.a(G602), .O(gate209inter7));
  inv1  gate1297(.a(G666), .O(gate209inter8));
  nand2 gate1298(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1299(.a(s_107), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1300(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1301(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1302(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate729(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate730(.a(gate219inter0), .b(s_26), .O(gate219inter1));
  and2  gate731(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate732(.a(s_26), .O(gate219inter3));
  inv1  gate733(.a(s_27), .O(gate219inter4));
  nand2 gate734(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate735(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate736(.a(G632), .O(gate219inter7));
  inv1  gate737(.a(G681), .O(gate219inter8));
  nand2 gate738(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate739(.a(s_27), .b(gate219inter3), .O(gate219inter10));
  nor2  gate740(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate741(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate742(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate659(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate660(.a(gate221inter0), .b(s_16), .O(gate221inter1));
  and2  gate661(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate662(.a(s_16), .O(gate221inter3));
  inv1  gate663(.a(s_17), .O(gate221inter4));
  nand2 gate664(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate665(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate666(.a(G622), .O(gate221inter7));
  inv1  gate667(.a(G684), .O(gate221inter8));
  nand2 gate668(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate669(.a(s_17), .b(gate221inter3), .O(gate221inter10));
  nor2  gate670(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate671(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate672(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate981(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate982(.a(gate224inter0), .b(s_62), .O(gate224inter1));
  and2  gate983(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate984(.a(s_62), .O(gate224inter3));
  inv1  gate985(.a(s_63), .O(gate224inter4));
  nand2 gate986(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate987(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate988(.a(G637), .O(gate224inter7));
  inv1  gate989(.a(G687), .O(gate224inter8));
  nand2 gate990(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate991(.a(s_63), .b(gate224inter3), .O(gate224inter10));
  nor2  gate992(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate993(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate994(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1583(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1584(.a(gate228inter0), .b(s_148), .O(gate228inter1));
  and2  gate1585(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1586(.a(s_148), .O(gate228inter3));
  inv1  gate1587(.a(s_149), .O(gate228inter4));
  nand2 gate1588(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1589(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1590(.a(G696), .O(gate228inter7));
  inv1  gate1591(.a(G697), .O(gate228inter8));
  nand2 gate1592(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1593(.a(s_149), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1594(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1595(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1596(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate869(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate870(.a(gate230inter0), .b(s_46), .O(gate230inter1));
  and2  gate871(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate872(.a(s_46), .O(gate230inter3));
  inv1  gate873(.a(s_47), .O(gate230inter4));
  nand2 gate874(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate875(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate876(.a(G700), .O(gate230inter7));
  inv1  gate877(.a(G701), .O(gate230inter8));
  nand2 gate878(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate879(.a(s_47), .b(gate230inter3), .O(gate230inter10));
  nor2  gate880(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate881(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate882(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1023(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1024(.a(gate243inter0), .b(s_68), .O(gate243inter1));
  and2  gate1025(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1026(.a(s_68), .O(gate243inter3));
  inv1  gate1027(.a(s_69), .O(gate243inter4));
  nand2 gate1028(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1029(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1030(.a(G245), .O(gate243inter7));
  inv1  gate1031(.a(G733), .O(gate243inter8));
  nand2 gate1032(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1033(.a(s_69), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1034(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1035(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1036(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate995(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate996(.a(gate259inter0), .b(s_64), .O(gate259inter1));
  and2  gate997(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate998(.a(s_64), .O(gate259inter3));
  inv1  gate999(.a(s_65), .O(gate259inter4));
  nand2 gate1000(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1001(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1002(.a(G758), .O(gate259inter7));
  inv1  gate1003(.a(G759), .O(gate259inter8));
  nand2 gate1004(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1005(.a(s_65), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1006(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1007(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1008(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate953(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate954(.a(gate262inter0), .b(s_58), .O(gate262inter1));
  and2  gate955(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate956(.a(s_58), .O(gate262inter3));
  inv1  gate957(.a(s_59), .O(gate262inter4));
  nand2 gate958(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate959(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate960(.a(G764), .O(gate262inter7));
  inv1  gate961(.a(G765), .O(gate262inter8));
  nand2 gate962(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate963(.a(s_59), .b(gate262inter3), .O(gate262inter10));
  nor2  gate964(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate965(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate966(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1261(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1262(.a(gate273inter0), .b(s_102), .O(gate273inter1));
  and2  gate1263(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1264(.a(s_102), .O(gate273inter3));
  inv1  gate1265(.a(s_103), .O(gate273inter4));
  nand2 gate1266(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1267(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1268(.a(G642), .O(gate273inter7));
  inv1  gate1269(.a(G794), .O(gate273inter8));
  nand2 gate1270(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1271(.a(s_103), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1272(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1273(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1274(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1443(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1444(.a(gate278inter0), .b(s_128), .O(gate278inter1));
  and2  gate1445(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1446(.a(s_128), .O(gate278inter3));
  inv1  gate1447(.a(s_129), .O(gate278inter4));
  nand2 gate1448(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1449(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1450(.a(G776), .O(gate278inter7));
  inv1  gate1451(.a(G800), .O(gate278inter8));
  nand2 gate1452(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1453(.a(s_129), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1454(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1455(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1456(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1093(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1094(.a(gate295inter0), .b(s_78), .O(gate295inter1));
  and2  gate1095(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1096(.a(s_78), .O(gate295inter3));
  inv1  gate1097(.a(s_79), .O(gate295inter4));
  nand2 gate1098(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1099(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1100(.a(G830), .O(gate295inter7));
  inv1  gate1101(.a(G831), .O(gate295inter8));
  nand2 gate1102(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1103(.a(s_79), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1104(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1105(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1106(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate883(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate884(.a(gate388inter0), .b(s_48), .O(gate388inter1));
  and2  gate885(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate886(.a(s_48), .O(gate388inter3));
  inv1  gate887(.a(s_49), .O(gate388inter4));
  nand2 gate888(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate889(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate890(.a(G2), .O(gate388inter7));
  inv1  gate891(.a(G1039), .O(gate388inter8));
  nand2 gate892(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate893(.a(s_49), .b(gate388inter3), .O(gate388inter10));
  nor2  gate894(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate895(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate896(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate939(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate940(.a(gate396inter0), .b(s_56), .O(gate396inter1));
  and2  gate941(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate942(.a(s_56), .O(gate396inter3));
  inv1  gate943(.a(s_57), .O(gate396inter4));
  nand2 gate944(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate945(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate946(.a(G10), .O(gate396inter7));
  inv1  gate947(.a(G1063), .O(gate396inter8));
  nand2 gate948(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate949(.a(s_57), .b(gate396inter3), .O(gate396inter10));
  nor2  gate950(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate951(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate952(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1387(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1388(.a(gate419inter0), .b(s_120), .O(gate419inter1));
  and2  gate1389(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1390(.a(s_120), .O(gate419inter3));
  inv1  gate1391(.a(s_121), .O(gate419inter4));
  nand2 gate1392(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1393(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1394(.a(G1), .O(gate419inter7));
  inv1  gate1395(.a(G1132), .O(gate419inter8));
  nand2 gate1396(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1397(.a(s_121), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1398(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1399(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1400(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1541(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1542(.a(gate432inter0), .b(s_142), .O(gate432inter1));
  and2  gate1543(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1544(.a(s_142), .O(gate432inter3));
  inv1  gate1545(.a(s_143), .O(gate432inter4));
  nand2 gate1546(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1547(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1548(.a(G1054), .O(gate432inter7));
  inv1  gate1549(.a(G1150), .O(gate432inter8));
  nand2 gate1550(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1551(.a(s_143), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1552(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1553(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1554(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1373(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1374(.a(gate433inter0), .b(s_118), .O(gate433inter1));
  and2  gate1375(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1376(.a(s_118), .O(gate433inter3));
  inv1  gate1377(.a(s_119), .O(gate433inter4));
  nand2 gate1378(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1379(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1380(.a(G8), .O(gate433inter7));
  inv1  gate1381(.a(G1153), .O(gate433inter8));
  nand2 gate1382(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1383(.a(s_119), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1384(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1385(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1386(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate645(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate646(.a(gate436inter0), .b(s_14), .O(gate436inter1));
  and2  gate647(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate648(.a(s_14), .O(gate436inter3));
  inv1  gate649(.a(s_15), .O(gate436inter4));
  nand2 gate650(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate651(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate652(.a(G1060), .O(gate436inter7));
  inv1  gate653(.a(G1156), .O(gate436inter8));
  nand2 gate654(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate655(.a(s_15), .b(gate436inter3), .O(gate436inter10));
  nor2  gate656(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate657(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate658(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1513(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1514(.a(gate437inter0), .b(s_138), .O(gate437inter1));
  and2  gate1515(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1516(.a(s_138), .O(gate437inter3));
  inv1  gate1517(.a(s_139), .O(gate437inter4));
  nand2 gate1518(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1519(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1520(.a(G10), .O(gate437inter7));
  inv1  gate1521(.a(G1159), .O(gate437inter8));
  nand2 gate1522(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1523(.a(s_139), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1524(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1525(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1526(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1485(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1486(.a(gate439inter0), .b(s_134), .O(gate439inter1));
  and2  gate1487(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1488(.a(s_134), .O(gate439inter3));
  inv1  gate1489(.a(s_135), .O(gate439inter4));
  nand2 gate1490(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1491(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1492(.a(G11), .O(gate439inter7));
  inv1  gate1493(.a(G1162), .O(gate439inter8));
  nand2 gate1494(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1495(.a(s_135), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1496(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1497(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1498(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate589(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate590(.a(gate441inter0), .b(s_6), .O(gate441inter1));
  and2  gate591(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate592(.a(s_6), .O(gate441inter3));
  inv1  gate593(.a(s_7), .O(gate441inter4));
  nand2 gate594(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate595(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate596(.a(G12), .O(gate441inter7));
  inv1  gate597(.a(G1165), .O(gate441inter8));
  nand2 gate598(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate599(.a(s_7), .b(gate441inter3), .O(gate441inter10));
  nor2  gate600(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate601(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate602(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1527(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1528(.a(gate445inter0), .b(s_140), .O(gate445inter1));
  and2  gate1529(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1530(.a(s_140), .O(gate445inter3));
  inv1  gate1531(.a(s_141), .O(gate445inter4));
  nand2 gate1532(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1533(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1534(.a(G14), .O(gate445inter7));
  inv1  gate1535(.a(G1171), .O(gate445inter8));
  nand2 gate1536(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1537(.a(s_141), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1538(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1539(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1540(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1569(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1570(.a(gate455inter0), .b(s_146), .O(gate455inter1));
  and2  gate1571(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1572(.a(s_146), .O(gate455inter3));
  inv1  gate1573(.a(s_147), .O(gate455inter4));
  nand2 gate1574(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1575(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1576(.a(G19), .O(gate455inter7));
  inv1  gate1577(.a(G1186), .O(gate455inter8));
  nand2 gate1578(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1579(.a(s_147), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1580(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1581(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1582(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1597(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1598(.a(gate458inter0), .b(s_150), .O(gate458inter1));
  and2  gate1599(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1600(.a(s_150), .O(gate458inter3));
  inv1  gate1601(.a(s_151), .O(gate458inter4));
  nand2 gate1602(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1603(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1604(.a(G1093), .O(gate458inter7));
  inv1  gate1605(.a(G1189), .O(gate458inter8));
  nand2 gate1606(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1607(.a(s_151), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1608(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1609(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1610(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1625(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1626(.a(gate461inter0), .b(s_154), .O(gate461inter1));
  and2  gate1627(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1628(.a(s_154), .O(gate461inter3));
  inv1  gate1629(.a(s_155), .O(gate461inter4));
  nand2 gate1630(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1631(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1632(.a(G22), .O(gate461inter7));
  inv1  gate1633(.a(G1195), .O(gate461inter8));
  nand2 gate1634(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1635(.a(s_155), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1636(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1637(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1638(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1415(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1416(.a(gate469inter0), .b(s_124), .O(gate469inter1));
  and2  gate1417(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1418(.a(s_124), .O(gate469inter3));
  inv1  gate1419(.a(s_125), .O(gate469inter4));
  nand2 gate1420(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1421(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1422(.a(G26), .O(gate469inter7));
  inv1  gate1423(.a(G1207), .O(gate469inter8));
  nand2 gate1424(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1425(.a(s_125), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1426(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1427(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1428(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1219(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1220(.a(gate472inter0), .b(s_96), .O(gate472inter1));
  and2  gate1221(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1222(.a(s_96), .O(gate472inter3));
  inv1  gate1223(.a(s_97), .O(gate472inter4));
  nand2 gate1224(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1225(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1226(.a(G1114), .O(gate472inter7));
  inv1  gate1227(.a(G1210), .O(gate472inter8));
  nand2 gate1228(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1229(.a(s_97), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1230(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1231(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1232(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1471(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1472(.a(gate474inter0), .b(s_132), .O(gate474inter1));
  and2  gate1473(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1474(.a(s_132), .O(gate474inter3));
  inv1  gate1475(.a(s_133), .O(gate474inter4));
  nand2 gate1476(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1477(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1478(.a(G1117), .O(gate474inter7));
  inv1  gate1479(.a(G1213), .O(gate474inter8));
  nand2 gate1480(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1481(.a(s_133), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1482(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1483(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1484(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1359(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1360(.a(gate475inter0), .b(s_116), .O(gate475inter1));
  and2  gate1361(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1362(.a(s_116), .O(gate475inter3));
  inv1  gate1363(.a(s_117), .O(gate475inter4));
  nand2 gate1364(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1365(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1366(.a(G29), .O(gate475inter7));
  inv1  gate1367(.a(G1216), .O(gate475inter8));
  nand2 gate1368(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1369(.a(s_117), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1370(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1371(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1372(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1079(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1080(.a(gate486inter0), .b(s_76), .O(gate486inter1));
  and2  gate1081(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1082(.a(s_76), .O(gate486inter3));
  inv1  gate1083(.a(s_77), .O(gate486inter4));
  nand2 gate1084(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1085(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1086(.a(G1234), .O(gate486inter7));
  inv1  gate1087(.a(G1235), .O(gate486inter8));
  nand2 gate1088(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1089(.a(s_77), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1090(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1091(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1092(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1191(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1192(.a(gate488inter0), .b(s_92), .O(gate488inter1));
  and2  gate1193(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1194(.a(s_92), .O(gate488inter3));
  inv1  gate1195(.a(s_93), .O(gate488inter4));
  nand2 gate1196(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1197(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1198(.a(G1238), .O(gate488inter7));
  inv1  gate1199(.a(G1239), .O(gate488inter8));
  nand2 gate1200(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1201(.a(s_93), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1202(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1203(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1204(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate575(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate576(.a(gate490inter0), .b(s_4), .O(gate490inter1));
  and2  gate577(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate578(.a(s_4), .O(gate490inter3));
  inv1  gate579(.a(s_5), .O(gate490inter4));
  nand2 gate580(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate581(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate582(.a(G1242), .O(gate490inter7));
  inv1  gate583(.a(G1243), .O(gate490inter8));
  nand2 gate584(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate585(.a(s_5), .b(gate490inter3), .O(gate490inter10));
  nor2  gate586(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate587(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate588(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1065(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1066(.a(gate495inter0), .b(s_74), .O(gate495inter1));
  and2  gate1067(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1068(.a(s_74), .O(gate495inter3));
  inv1  gate1069(.a(s_75), .O(gate495inter4));
  nand2 gate1070(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1071(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1072(.a(G1252), .O(gate495inter7));
  inv1  gate1073(.a(G1253), .O(gate495inter8));
  nand2 gate1074(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1075(.a(s_75), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1076(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1077(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1078(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1457(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1458(.a(gate499inter0), .b(s_130), .O(gate499inter1));
  and2  gate1459(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1460(.a(s_130), .O(gate499inter3));
  inv1  gate1461(.a(s_131), .O(gate499inter4));
  nand2 gate1462(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1463(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1464(.a(G1260), .O(gate499inter7));
  inv1  gate1465(.a(G1261), .O(gate499inter8));
  nand2 gate1466(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1467(.a(s_131), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1468(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1469(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1470(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate799(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate800(.a(gate501inter0), .b(s_36), .O(gate501inter1));
  and2  gate801(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate802(.a(s_36), .O(gate501inter3));
  inv1  gate803(.a(s_37), .O(gate501inter4));
  nand2 gate804(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate805(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate806(.a(G1264), .O(gate501inter7));
  inv1  gate807(.a(G1265), .O(gate501inter8));
  nand2 gate808(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate809(.a(s_37), .b(gate501inter3), .O(gate501inter10));
  nor2  gate810(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate811(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate812(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule