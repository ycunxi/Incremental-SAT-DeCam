module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1037(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1038(.a(gate13inter0), .b(s_70), .O(gate13inter1));
  and2  gate1039(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1040(.a(s_70), .O(gate13inter3));
  inv1  gate1041(.a(s_71), .O(gate13inter4));
  nand2 gate1042(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1043(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1044(.a(G9), .O(gate13inter7));
  inv1  gate1045(.a(G10), .O(gate13inter8));
  nand2 gate1046(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1047(.a(s_71), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1048(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1049(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1050(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1961(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1962(.a(gate14inter0), .b(s_202), .O(gate14inter1));
  and2  gate1963(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1964(.a(s_202), .O(gate14inter3));
  inv1  gate1965(.a(s_203), .O(gate14inter4));
  nand2 gate1966(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1967(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1968(.a(G11), .O(gate14inter7));
  inv1  gate1969(.a(G12), .O(gate14inter8));
  nand2 gate1970(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1971(.a(s_203), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1972(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1973(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1974(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1891(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1892(.a(gate15inter0), .b(s_192), .O(gate15inter1));
  and2  gate1893(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1894(.a(s_192), .O(gate15inter3));
  inv1  gate1895(.a(s_193), .O(gate15inter4));
  nand2 gate1896(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1897(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1898(.a(G13), .O(gate15inter7));
  inv1  gate1899(.a(G14), .O(gate15inter8));
  nand2 gate1900(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1901(.a(s_193), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1902(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1903(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1904(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1121(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1122(.a(gate19inter0), .b(s_82), .O(gate19inter1));
  and2  gate1123(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1124(.a(s_82), .O(gate19inter3));
  inv1  gate1125(.a(s_83), .O(gate19inter4));
  nand2 gate1126(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1127(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1128(.a(G21), .O(gate19inter7));
  inv1  gate1129(.a(G22), .O(gate19inter8));
  nand2 gate1130(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1131(.a(s_83), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1132(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1133(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1134(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1457(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1458(.a(gate21inter0), .b(s_130), .O(gate21inter1));
  and2  gate1459(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1460(.a(s_130), .O(gate21inter3));
  inv1  gate1461(.a(s_131), .O(gate21inter4));
  nand2 gate1462(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1463(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1464(.a(G25), .O(gate21inter7));
  inv1  gate1465(.a(G26), .O(gate21inter8));
  nand2 gate1466(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1467(.a(s_131), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1468(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1469(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1470(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1611(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1612(.a(gate34inter0), .b(s_152), .O(gate34inter1));
  and2  gate1613(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1614(.a(s_152), .O(gate34inter3));
  inv1  gate1615(.a(s_153), .O(gate34inter4));
  nand2 gate1616(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1617(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1618(.a(G25), .O(gate34inter7));
  inv1  gate1619(.a(G29), .O(gate34inter8));
  nand2 gate1620(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1621(.a(s_153), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1622(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1623(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1624(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate743(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate744(.a(gate38inter0), .b(s_28), .O(gate38inter1));
  and2  gate745(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate746(.a(s_28), .O(gate38inter3));
  inv1  gate747(.a(s_29), .O(gate38inter4));
  nand2 gate748(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate749(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate750(.a(G27), .O(gate38inter7));
  inv1  gate751(.a(G31), .O(gate38inter8));
  nand2 gate752(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate753(.a(s_29), .b(gate38inter3), .O(gate38inter10));
  nor2  gate754(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate755(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate756(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1821(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1822(.a(gate45inter0), .b(s_182), .O(gate45inter1));
  and2  gate1823(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1824(.a(s_182), .O(gate45inter3));
  inv1  gate1825(.a(s_183), .O(gate45inter4));
  nand2 gate1826(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1827(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1828(.a(G5), .O(gate45inter7));
  inv1  gate1829(.a(G272), .O(gate45inter8));
  nand2 gate1830(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1831(.a(s_183), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1832(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1833(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1834(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1093(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1094(.a(gate52inter0), .b(s_78), .O(gate52inter1));
  and2  gate1095(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1096(.a(s_78), .O(gate52inter3));
  inv1  gate1097(.a(s_79), .O(gate52inter4));
  nand2 gate1098(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1099(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1100(.a(G12), .O(gate52inter7));
  inv1  gate1101(.a(G281), .O(gate52inter8));
  nand2 gate1102(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1103(.a(s_79), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1104(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1105(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1106(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate855(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate856(.a(gate54inter0), .b(s_44), .O(gate54inter1));
  and2  gate857(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate858(.a(s_44), .O(gate54inter3));
  inv1  gate859(.a(s_45), .O(gate54inter4));
  nand2 gate860(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate861(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate862(.a(G14), .O(gate54inter7));
  inv1  gate863(.a(G284), .O(gate54inter8));
  nand2 gate864(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate865(.a(s_45), .b(gate54inter3), .O(gate54inter10));
  nor2  gate866(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate867(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate868(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1527(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1528(.a(gate58inter0), .b(s_140), .O(gate58inter1));
  and2  gate1529(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1530(.a(s_140), .O(gate58inter3));
  inv1  gate1531(.a(s_141), .O(gate58inter4));
  nand2 gate1532(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1533(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1534(.a(G18), .O(gate58inter7));
  inv1  gate1535(.a(G290), .O(gate58inter8));
  nand2 gate1536(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1537(.a(s_141), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1538(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1539(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1540(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate813(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate814(.a(gate61inter0), .b(s_38), .O(gate61inter1));
  and2  gate815(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate816(.a(s_38), .O(gate61inter3));
  inv1  gate817(.a(s_39), .O(gate61inter4));
  nand2 gate818(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate819(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate820(.a(G21), .O(gate61inter7));
  inv1  gate821(.a(G296), .O(gate61inter8));
  nand2 gate822(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate823(.a(s_39), .b(gate61inter3), .O(gate61inter10));
  nor2  gate824(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate825(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate826(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1247(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1248(.a(gate64inter0), .b(s_100), .O(gate64inter1));
  and2  gate1249(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1250(.a(s_100), .O(gate64inter3));
  inv1  gate1251(.a(s_101), .O(gate64inter4));
  nand2 gate1252(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1253(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1254(.a(G24), .O(gate64inter7));
  inv1  gate1255(.a(G299), .O(gate64inter8));
  nand2 gate1256(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1257(.a(s_101), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1258(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1259(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1260(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate547(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate548(.a(gate65inter0), .b(s_0), .O(gate65inter1));
  and2  gate549(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate550(.a(s_0), .O(gate65inter3));
  inv1  gate551(.a(s_1), .O(gate65inter4));
  nand2 gate552(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate553(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate554(.a(G25), .O(gate65inter7));
  inv1  gate555(.a(G302), .O(gate65inter8));
  nand2 gate556(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate557(.a(s_1), .b(gate65inter3), .O(gate65inter10));
  nor2  gate558(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate559(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate560(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate995(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate996(.a(gate73inter0), .b(s_64), .O(gate73inter1));
  and2  gate997(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate998(.a(s_64), .O(gate73inter3));
  inv1  gate999(.a(s_65), .O(gate73inter4));
  nand2 gate1000(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1001(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1002(.a(G1), .O(gate73inter7));
  inv1  gate1003(.a(G314), .O(gate73inter8));
  nand2 gate1004(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1005(.a(s_65), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1006(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1007(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1008(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1359(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1360(.a(gate74inter0), .b(s_116), .O(gate74inter1));
  and2  gate1361(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1362(.a(s_116), .O(gate74inter3));
  inv1  gate1363(.a(s_117), .O(gate74inter4));
  nand2 gate1364(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1365(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1366(.a(G5), .O(gate74inter7));
  inv1  gate1367(.a(G314), .O(gate74inter8));
  nand2 gate1368(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1369(.a(s_117), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1370(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1371(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1372(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1863(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1864(.a(gate75inter0), .b(s_188), .O(gate75inter1));
  and2  gate1865(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1866(.a(s_188), .O(gate75inter3));
  inv1  gate1867(.a(s_189), .O(gate75inter4));
  nand2 gate1868(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1869(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1870(.a(G9), .O(gate75inter7));
  inv1  gate1871(.a(G317), .O(gate75inter8));
  nand2 gate1872(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1873(.a(s_189), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1874(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1875(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1876(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate603(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate604(.a(gate89inter0), .b(s_8), .O(gate89inter1));
  and2  gate605(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate606(.a(s_8), .O(gate89inter3));
  inv1  gate607(.a(s_9), .O(gate89inter4));
  nand2 gate608(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate609(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate610(.a(G17), .O(gate89inter7));
  inv1  gate611(.a(G338), .O(gate89inter8));
  nand2 gate612(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate613(.a(s_9), .b(gate89inter3), .O(gate89inter10));
  nor2  gate614(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate615(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate616(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1597(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1598(.a(gate90inter0), .b(s_150), .O(gate90inter1));
  and2  gate1599(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1600(.a(s_150), .O(gate90inter3));
  inv1  gate1601(.a(s_151), .O(gate90inter4));
  nand2 gate1602(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1603(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1604(.a(G21), .O(gate90inter7));
  inv1  gate1605(.a(G338), .O(gate90inter8));
  nand2 gate1606(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1607(.a(s_151), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1608(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1609(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1610(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1723(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1724(.a(gate93inter0), .b(s_168), .O(gate93inter1));
  and2  gate1725(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1726(.a(s_168), .O(gate93inter3));
  inv1  gate1727(.a(s_169), .O(gate93inter4));
  nand2 gate1728(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1729(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1730(.a(G18), .O(gate93inter7));
  inv1  gate1731(.a(G344), .O(gate93inter8));
  nand2 gate1732(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1733(.a(s_169), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1734(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1735(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1736(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1429(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1430(.a(gate97inter0), .b(s_126), .O(gate97inter1));
  and2  gate1431(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1432(.a(s_126), .O(gate97inter3));
  inv1  gate1433(.a(s_127), .O(gate97inter4));
  nand2 gate1434(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1435(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1436(.a(G19), .O(gate97inter7));
  inv1  gate1437(.a(G350), .O(gate97inter8));
  nand2 gate1438(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1439(.a(s_127), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1440(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1441(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1442(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate897(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate898(.a(gate98inter0), .b(s_50), .O(gate98inter1));
  and2  gate899(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate900(.a(s_50), .O(gate98inter3));
  inv1  gate901(.a(s_51), .O(gate98inter4));
  nand2 gate902(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate903(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate904(.a(G23), .O(gate98inter7));
  inv1  gate905(.a(G350), .O(gate98inter8));
  nand2 gate906(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate907(.a(s_51), .b(gate98inter3), .O(gate98inter10));
  nor2  gate908(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate909(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate910(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate687(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate688(.a(gate99inter0), .b(s_20), .O(gate99inter1));
  and2  gate689(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate690(.a(s_20), .O(gate99inter3));
  inv1  gate691(.a(s_21), .O(gate99inter4));
  nand2 gate692(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate693(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate694(.a(G27), .O(gate99inter7));
  inv1  gate695(.a(G353), .O(gate99inter8));
  nand2 gate696(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate697(.a(s_21), .b(gate99inter3), .O(gate99inter10));
  nor2  gate698(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate699(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate700(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1331(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1332(.a(gate109inter0), .b(s_112), .O(gate109inter1));
  and2  gate1333(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1334(.a(s_112), .O(gate109inter3));
  inv1  gate1335(.a(s_113), .O(gate109inter4));
  nand2 gate1336(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1337(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1338(.a(G370), .O(gate109inter7));
  inv1  gate1339(.a(G371), .O(gate109inter8));
  nand2 gate1340(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1341(.a(s_113), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1342(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1343(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1344(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1975(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1976(.a(gate112inter0), .b(s_204), .O(gate112inter1));
  and2  gate1977(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1978(.a(s_204), .O(gate112inter3));
  inv1  gate1979(.a(s_205), .O(gate112inter4));
  nand2 gate1980(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1981(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1982(.a(G376), .O(gate112inter7));
  inv1  gate1983(.a(G377), .O(gate112inter8));
  nand2 gate1984(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1985(.a(s_205), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1986(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1987(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1988(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate575(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate576(.a(gate113inter0), .b(s_4), .O(gate113inter1));
  and2  gate577(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate578(.a(s_4), .O(gate113inter3));
  inv1  gate579(.a(s_5), .O(gate113inter4));
  nand2 gate580(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate581(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate582(.a(G378), .O(gate113inter7));
  inv1  gate583(.a(G379), .O(gate113inter8));
  nand2 gate584(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate585(.a(s_5), .b(gate113inter3), .O(gate113inter10));
  nor2  gate586(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate587(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate588(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1233(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1234(.a(gate116inter0), .b(s_98), .O(gate116inter1));
  and2  gate1235(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1236(.a(s_98), .O(gate116inter3));
  inv1  gate1237(.a(s_99), .O(gate116inter4));
  nand2 gate1238(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1239(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1240(.a(G384), .O(gate116inter7));
  inv1  gate1241(.a(G385), .O(gate116inter8));
  nand2 gate1242(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1243(.a(s_99), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1244(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1245(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1246(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1569(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1570(.a(gate119inter0), .b(s_146), .O(gate119inter1));
  and2  gate1571(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1572(.a(s_146), .O(gate119inter3));
  inv1  gate1573(.a(s_147), .O(gate119inter4));
  nand2 gate1574(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1575(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1576(.a(G390), .O(gate119inter7));
  inv1  gate1577(.a(G391), .O(gate119inter8));
  nand2 gate1578(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1579(.a(s_147), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1580(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1581(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1582(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1205(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1206(.a(gate123inter0), .b(s_94), .O(gate123inter1));
  and2  gate1207(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1208(.a(s_94), .O(gate123inter3));
  inv1  gate1209(.a(s_95), .O(gate123inter4));
  nand2 gate1210(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1211(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1212(.a(G398), .O(gate123inter7));
  inv1  gate1213(.a(G399), .O(gate123inter8));
  nand2 gate1214(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1215(.a(s_95), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1216(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1217(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1218(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate841(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate842(.a(gate126inter0), .b(s_42), .O(gate126inter1));
  and2  gate843(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate844(.a(s_42), .O(gate126inter3));
  inv1  gate845(.a(s_43), .O(gate126inter4));
  nand2 gate846(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate847(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate848(.a(G404), .O(gate126inter7));
  inv1  gate849(.a(G405), .O(gate126inter8));
  nand2 gate850(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate851(.a(s_43), .b(gate126inter3), .O(gate126inter10));
  nor2  gate852(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate853(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate854(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1653(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1654(.a(gate129inter0), .b(s_158), .O(gate129inter1));
  and2  gate1655(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1656(.a(s_158), .O(gate129inter3));
  inv1  gate1657(.a(s_159), .O(gate129inter4));
  nand2 gate1658(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1659(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1660(.a(G410), .O(gate129inter7));
  inv1  gate1661(.a(G411), .O(gate129inter8));
  nand2 gate1662(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1663(.a(s_159), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1664(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1665(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1666(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate799(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate800(.a(gate131inter0), .b(s_36), .O(gate131inter1));
  and2  gate801(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate802(.a(s_36), .O(gate131inter3));
  inv1  gate803(.a(s_37), .O(gate131inter4));
  nand2 gate804(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate805(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate806(.a(G414), .O(gate131inter7));
  inv1  gate807(.a(G415), .O(gate131inter8));
  nand2 gate808(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate809(.a(s_37), .b(gate131inter3), .O(gate131inter10));
  nor2  gate810(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate811(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate812(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1779(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1780(.a(gate140inter0), .b(s_176), .O(gate140inter1));
  and2  gate1781(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1782(.a(s_176), .O(gate140inter3));
  inv1  gate1783(.a(s_177), .O(gate140inter4));
  nand2 gate1784(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1785(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1786(.a(G444), .O(gate140inter7));
  inv1  gate1787(.a(G447), .O(gate140inter8));
  nand2 gate1788(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1789(.a(s_177), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1790(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1791(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1792(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1009(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1010(.a(gate143inter0), .b(s_66), .O(gate143inter1));
  and2  gate1011(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1012(.a(s_66), .O(gate143inter3));
  inv1  gate1013(.a(s_67), .O(gate143inter4));
  nand2 gate1014(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1015(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1016(.a(G462), .O(gate143inter7));
  inv1  gate1017(.a(G465), .O(gate143inter8));
  nand2 gate1018(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1019(.a(s_67), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1020(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1021(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1022(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1947(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1948(.a(gate147inter0), .b(s_200), .O(gate147inter1));
  and2  gate1949(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1950(.a(s_200), .O(gate147inter3));
  inv1  gate1951(.a(s_201), .O(gate147inter4));
  nand2 gate1952(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1953(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1954(.a(G486), .O(gate147inter7));
  inv1  gate1955(.a(G489), .O(gate147inter8));
  nand2 gate1956(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1957(.a(s_201), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1958(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1959(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1960(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1163(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1164(.a(gate149inter0), .b(s_88), .O(gate149inter1));
  and2  gate1165(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1166(.a(s_88), .O(gate149inter3));
  inv1  gate1167(.a(s_89), .O(gate149inter4));
  nand2 gate1168(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1169(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1170(.a(G498), .O(gate149inter7));
  inv1  gate1171(.a(G501), .O(gate149inter8));
  nand2 gate1172(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1173(.a(s_89), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1174(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1175(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1176(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1079(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1080(.a(gate151inter0), .b(s_76), .O(gate151inter1));
  and2  gate1081(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1082(.a(s_76), .O(gate151inter3));
  inv1  gate1083(.a(s_77), .O(gate151inter4));
  nand2 gate1084(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1085(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1086(.a(G510), .O(gate151inter7));
  inv1  gate1087(.a(G513), .O(gate151inter8));
  nand2 gate1088(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1089(.a(s_77), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1090(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1091(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1092(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate771(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate772(.a(gate155inter0), .b(s_32), .O(gate155inter1));
  and2  gate773(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate774(.a(s_32), .O(gate155inter3));
  inv1  gate775(.a(s_33), .O(gate155inter4));
  nand2 gate776(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate777(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate778(.a(G432), .O(gate155inter7));
  inv1  gate779(.a(G525), .O(gate155inter8));
  nand2 gate780(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate781(.a(s_33), .b(gate155inter3), .O(gate155inter10));
  nor2  gate782(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate783(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate784(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate981(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate982(.a(gate156inter0), .b(s_62), .O(gate156inter1));
  and2  gate983(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate984(.a(s_62), .O(gate156inter3));
  inv1  gate985(.a(s_63), .O(gate156inter4));
  nand2 gate986(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate987(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate988(.a(G435), .O(gate156inter7));
  inv1  gate989(.a(G525), .O(gate156inter8));
  nand2 gate990(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate991(.a(s_63), .b(gate156inter3), .O(gate156inter10));
  nor2  gate992(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate993(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate994(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1387(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1388(.a(gate157inter0), .b(s_120), .O(gate157inter1));
  and2  gate1389(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1390(.a(s_120), .O(gate157inter3));
  inv1  gate1391(.a(s_121), .O(gate157inter4));
  nand2 gate1392(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1393(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1394(.a(G438), .O(gate157inter7));
  inv1  gate1395(.a(G528), .O(gate157inter8));
  nand2 gate1396(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1397(.a(s_121), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1398(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1399(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1400(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate631(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate632(.a(gate160inter0), .b(s_12), .O(gate160inter1));
  and2  gate633(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate634(.a(s_12), .O(gate160inter3));
  inv1  gate635(.a(s_13), .O(gate160inter4));
  nand2 gate636(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate637(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate638(.a(G447), .O(gate160inter7));
  inv1  gate639(.a(G531), .O(gate160inter8));
  nand2 gate640(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate641(.a(s_13), .b(gate160inter3), .O(gate160inter10));
  nor2  gate642(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate643(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate644(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1107(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1108(.a(gate162inter0), .b(s_80), .O(gate162inter1));
  and2  gate1109(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1110(.a(s_80), .O(gate162inter3));
  inv1  gate1111(.a(s_81), .O(gate162inter4));
  nand2 gate1112(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1113(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1114(.a(G453), .O(gate162inter7));
  inv1  gate1115(.a(G534), .O(gate162inter8));
  nand2 gate1116(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1117(.a(s_81), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1118(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1119(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1120(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2003(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2004(.a(gate163inter0), .b(s_208), .O(gate163inter1));
  and2  gate2005(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2006(.a(s_208), .O(gate163inter3));
  inv1  gate2007(.a(s_209), .O(gate163inter4));
  nand2 gate2008(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2009(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2010(.a(G456), .O(gate163inter7));
  inv1  gate2011(.a(G537), .O(gate163inter8));
  nand2 gate2012(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2013(.a(s_209), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2014(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2015(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2016(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1051(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1052(.a(gate169inter0), .b(s_72), .O(gate169inter1));
  and2  gate1053(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1054(.a(s_72), .O(gate169inter3));
  inv1  gate1055(.a(s_73), .O(gate169inter4));
  nand2 gate1056(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1057(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1058(.a(G474), .O(gate169inter7));
  inv1  gate1059(.a(G546), .O(gate169inter8));
  nand2 gate1060(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1061(.a(s_73), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1062(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1063(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1064(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate659(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate660(.a(gate175inter0), .b(s_16), .O(gate175inter1));
  and2  gate661(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate662(.a(s_16), .O(gate175inter3));
  inv1  gate663(.a(s_17), .O(gate175inter4));
  nand2 gate664(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate665(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate666(.a(G492), .O(gate175inter7));
  inv1  gate667(.a(G555), .O(gate175inter8));
  nand2 gate668(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate669(.a(s_17), .b(gate175inter3), .O(gate175inter10));
  nor2  gate670(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate671(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate672(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate715(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate716(.a(gate178inter0), .b(s_24), .O(gate178inter1));
  and2  gate717(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate718(.a(s_24), .O(gate178inter3));
  inv1  gate719(.a(s_25), .O(gate178inter4));
  nand2 gate720(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate721(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate722(.a(G501), .O(gate178inter7));
  inv1  gate723(.a(G558), .O(gate178inter8));
  nand2 gate724(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate725(.a(s_25), .b(gate178inter3), .O(gate178inter10));
  nor2  gate726(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate727(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate728(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1149(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1150(.a(gate180inter0), .b(s_86), .O(gate180inter1));
  and2  gate1151(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1152(.a(s_86), .O(gate180inter3));
  inv1  gate1153(.a(s_87), .O(gate180inter4));
  nand2 gate1154(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1155(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1156(.a(G507), .O(gate180inter7));
  inv1  gate1157(.a(G561), .O(gate180inter8));
  nand2 gate1158(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1159(.a(s_87), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1160(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1161(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1162(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1317(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1318(.a(gate182inter0), .b(s_110), .O(gate182inter1));
  and2  gate1319(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1320(.a(s_110), .O(gate182inter3));
  inv1  gate1321(.a(s_111), .O(gate182inter4));
  nand2 gate1322(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1323(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1324(.a(G513), .O(gate182inter7));
  inv1  gate1325(.a(G564), .O(gate182inter8));
  nand2 gate1326(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1327(.a(s_111), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1328(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1329(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1330(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate869(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate870(.a(gate184inter0), .b(s_46), .O(gate184inter1));
  and2  gate871(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate872(.a(s_46), .O(gate184inter3));
  inv1  gate873(.a(s_47), .O(gate184inter4));
  nand2 gate874(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate875(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate876(.a(G519), .O(gate184inter7));
  inv1  gate877(.a(G567), .O(gate184inter8));
  nand2 gate878(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate879(.a(s_47), .b(gate184inter3), .O(gate184inter10));
  nor2  gate880(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate881(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate882(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1373(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1374(.a(gate187inter0), .b(s_118), .O(gate187inter1));
  and2  gate1375(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1376(.a(s_118), .O(gate187inter3));
  inv1  gate1377(.a(s_119), .O(gate187inter4));
  nand2 gate1378(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1379(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1380(.a(G574), .O(gate187inter7));
  inv1  gate1381(.a(G575), .O(gate187inter8));
  nand2 gate1382(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1383(.a(s_119), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1384(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1385(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1386(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1191(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1192(.a(gate188inter0), .b(s_92), .O(gate188inter1));
  and2  gate1193(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1194(.a(s_92), .O(gate188inter3));
  inv1  gate1195(.a(s_93), .O(gate188inter4));
  nand2 gate1196(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1197(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1198(.a(G576), .O(gate188inter7));
  inv1  gate1199(.a(G577), .O(gate188inter8));
  nand2 gate1200(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1201(.a(s_93), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1202(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1203(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1204(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate785(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate786(.a(gate195inter0), .b(s_34), .O(gate195inter1));
  and2  gate787(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate788(.a(s_34), .O(gate195inter3));
  inv1  gate789(.a(s_35), .O(gate195inter4));
  nand2 gate790(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate791(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate792(.a(G590), .O(gate195inter7));
  inv1  gate793(.a(G591), .O(gate195inter8));
  nand2 gate794(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate795(.a(s_35), .b(gate195inter3), .O(gate195inter10));
  nor2  gate796(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate797(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate798(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate911(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate912(.a(gate198inter0), .b(s_52), .O(gate198inter1));
  and2  gate913(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate914(.a(s_52), .O(gate198inter3));
  inv1  gate915(.a(s_53), .O(gate198inter4));
  nand2 gate916(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate917(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate918(.a(G596), .O(gate198inter7));
  inv1  gate919(.a(G597), .O(gate198inter8));
  nand2 gate920(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate921(.a(s_53), .b(gate198inter3), .O(gate198inter10));
  nor2  gate922(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate923(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate924(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1751(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1752(.a(gate200inter0), .b(s_172), .O(gate200inter1));
  and2  gate1753(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1754(.a(s_172), .O(gate200inter3));
  inv1  gate1755(.a(s_173), .O(gate200inter4));
  nand2 gate1756(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1757(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1758(.a(G600), .O(gate200inter7));
  inv1  gate1759(.a(G601), .O(gate200inter8));
  nand2 gate1760(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1761(.a(s_173), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1762(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1763(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1764(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1023(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1024(.a(gate212inter0), .b(s_68), .O(gate212inter1));
  and2  gate1025(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1026(.a(s_68), .O(gate212inter3));
  inv1  gate1027(.a(s_69), .O(gate212inter4));
  nand2 gate1028(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1029(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1030(.a(G617), .O(gate212inter7));
  inv1  gate1031(.a(G669), .O(gate212inter8));
  nand2 gate1032(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1033(.a(s_69), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1034(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1035(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1036(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1471(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1472(.a(gate213inter0), .b(s_132), .O(gate213inter1));
  and2  gate1473(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1474(.a(s_132), .O(gate213inter3));
  inv1  gate1475(.a(s_133), .O(gate213inter4));
  nand2 gate1476(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1477(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1478(.a(G602), .O(gate213inter7));
  inv1  gate1479(.a(G672), .O(gate213inter8));
  nand2 gate1480(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1481(.a(s_133), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1482(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1483(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1484(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1555(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1556(.a(gate214inter0), .b(s_144), .O(gate214inter1));
  and2  gate1557(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1558(.a(s_144), .O(gate214inter3));
  inv1  gate1559(.a(s_145), .O(gate214inter4));
  nand2 gate1560(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1561(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1562(.a(G612), .O(gate214inter7));
  inv1  gate1563(.a(G672), .O(gate214inter8));
  nand2 gate1564(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1565(.a(s_145), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1566(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1567(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1568(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1415(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1416(.a(gate215inter0), .b(s_124), .O(gate215inter1));
  and2  gate1417(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1418(.a(s_124), .O(gate215inter3));
  inv1  gate1419(.a(s_125), .O(gate215inter4));
  nand2 gate1420(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1421(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1422(.a(G607), .O(gate215inter7));
  inv1  gate1423(.a(G675), .O(gate215inter8));
  nand2 gate1424(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1425(.a(s_125), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1426(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1427(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1428(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1639(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1640(.a(gate218inter0), .b(s_156), .O(gate218inter1));
  and2  gate1641(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1642(.a(s_156), .O(gate218inter3));
  inv1  gate1643(.a(s_157), .O(gate218inter4));
  nand2 gate1644(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1645(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1646(.a(G627), .O(gate218inter7));
  inv1  gate1647(.a(G678), .O(gate218inter8));
  nand2 gate1648(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1649(.a(s_157), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1650(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1651(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1652(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1849(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1850(.a(gate222inter0), .b(s_186), .O(gate222inter1));
  and2  gate1851(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1852(.a(s_186), .O(gate222inter3));
  inv1  gate1853(.a(s_187), .O(gate222inter4));
  nand2 gate1854(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1855(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1856(.a(G632), .O(gate222inter7));
  inv1  gate1857(.a(G684), .O(gate222inter8));
  nand2 gate1858(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1859(.a(s_187), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1860(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1861(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1862(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1583(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1584(.a(gate227inter0), .b(s_148), .O(gate227inter1));
  and2  gate1585(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1586(.a(s_148), .O(gate227inter3));
  inv1  gate1587(.a(s_149), .O(gate227inter4));
  nand2 gate1588(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1589(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1590(.a(G694), .O(gate227inter7));
  inv1  gate1591(.a(G695), .O(gate227inter8));
  nand2 gate1592(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1593(.a(s_149), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1594(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1595(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1596(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1499(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1500(.a(gate230inter0), .b(s_136), .O(gate230inter1));
  and2  gate1501(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1502(.a(s_136), .O(gate230inter3));
  inv1  gate1503(.a(s_137), .O(gate230inter4));
  nand2 gate1504(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1505(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1506(.a(G700), .O(gate230inter7));
  inv1  gate1507(.a(G701), .O(gate230inter8));
  nand2 gate1508(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1509(.a(s_137), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1510(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1511(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1512(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate883(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate884(.a(gate233inter0), .b(s_48), .O(gate233inter1));
  and2  gate885(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate886(.a(s_48), .O(gate233inter3));
  inv1  gate887(.a(s_49), .O(gate233inter4));
  nand2 gate888(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate889(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate890(.a(G242), .O(gate233inter7));
  inv1  gate891(.a(G718), .O(gate233inter8));
  nand2 gate892(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate893(.a(s_49), .b(gate233inter3), .O(gate233inter10));
  nor2  gate894(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate895(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate896(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1541(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1542(.a(gate239inter0), .b(s_142), .O(gate239inter1));
  and2  gate1543(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1544(.a(s_142), .O(gate239inter3));
  inv1  gate1545(.a(s_143), .O(gate239inter4));
  nand2 gate1546(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1547(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1548(.a(G260), .O(gate239inter7));
  inv1  gate1549(.a(G712), .O(gate239inter8));
  nand2 gate1550(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1551(.a(s_143), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1552(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1553(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1554(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1275(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1276(.a(gate243inter0), .b(s_104), .O(gate243inter1));
  and2  gate1277(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1278(.a(s_104), .O(gate243inter3));
  inv1  gate1279(.a(s_105), .O(gate243inter4));
  nand2 gate1280(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1281(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1282(.a(G245), .O(gate243inter7));
  inv1  gate1283(.a(G733), .O(gate243inter8));
  nand2 gate1284(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1285(.a(s_105), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1286(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1287(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1288(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1905(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1906(.a(gate248inter0), .b(s_194), .O(gate248inter1));
  and2  gate1907(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1908(.a(s_194), .O(gate248inter3));
  inv1  gate1909(.a(s_195), .O(gate248inter4));
  nand2 gate1910(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1911(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1912(.a(G727), .O(gate248inter7));
  inv1  gate1913(.a(G739), .O(gate248inter8));
  nand2 gate1914(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1915(.a(s_195), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1916(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1917(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1918(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1261(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1262(.a(gate250inter0), .b(s_102), .O(gate250inter1));
  and2  gate1263(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1264(.a(s_102), .O(gate250inter3));
  inv1  gate1265(.a(s_103), .O(gate250inter4));
  nand2 gate1266(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1267(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1268(.a(G706), .O(gate250inter7));
  inv1  gate1269(.a(G742), .O(gate250inter8));
  nand2 gate1270(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1271(.a(s_103), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1272(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1273(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1274(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1303(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1304(.a(gate254inter0), .b(s_108), .O(gate254inter1));
  and2  gate1305(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1306(.a(s_108), .O(gate254inter3));
  inv1  gate1307(.a(s_109), .O(gate254inter4));
  nand2 gate1308(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1309(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1310(.a(G712), .O(gate254inter7));
  inv1  gate1311(.a(G748), .O(gate254inter8));
  nand2 gate1312(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1313(.a(s_109), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1314(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1315(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1316(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1485(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1486(.a(gate264inter0), .b(s_134), .O(gate264inter1));
  and2  gate1487(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1488(.a(s_134), .O(gate264inter3));
  inv1  gate1489(.a(s_135), .O(gate264inter4));
  nand2 gate1490(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1491(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1492(.a(G768), .O(gate264inter7));
  inv1  gate1493(.a(G769), .O(gate264inter8));
  nand2 gate1494(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1495(.a(s_135), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1496(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1497(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1498(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2017(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2018(.a(gate271inter0), .b(s_210), .O(gate271inter1));
  and2  gate2019(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2020(.a(s_210), .O(gate271inter3));
  inv1  gate2021(.a(s_211), .O(gate271inter4));
  nand2 gate2022(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2023(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2024(.a(G660), .O(gate271inter7));
  inv1  gate2025(.a(G788), .O(gate271inter8));
  nand2 gate2026(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2027(.a(s_211), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2028(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2029(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2030(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1135(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1136(.a(gate282inter0), .b(s_84), .O(gate282inter1));
  and2  gate1137(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1138(.a(s_84), .O(gate282inter3));
  inv1  gate1139(.a(s_85), .O(gate282inter4));
  nand2 gate1140(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1141(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1142(.a(G782), .O(gate282inter7));
  inv1  gate1143(.a(G806), .O(gate282inter8));
  nand2 gate1144(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1145(.a(s_85), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1146(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1147(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1148(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1625(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1626(.a(gate284inter0), .b(s_154), .O(gate284inter1));
  and2  gate1627(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1628(.a(s_154), .O(gate284inter3));
  inv1  gate1629(.a(s_155), .O(gate284inter4));
  nand2 gate1630(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1631(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1632(.a(G785), .O(gate284inter7));
  inv1  gate1633(.a(G809), .O(gate284inter8));
  nand2 gate1634(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1635(.a(s_155), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1636(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1637(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1638(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1835(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1836(.a(gate285inter0), .b(s_184), .O(gate285inter1));
  and2  gate1837(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1838(.a(s_184), .O(gate285inter3));
  inv1  gate1839(.a(s_185), .O(gate285inter4));
  nand2 gate1840(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1841(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1842(.a(G660), .O(gate285inter7));
  inv1  gate1843(.a(G812), .O(gate285inter8));
  nand2 gate1844(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1845(.a(s_185), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1846(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1847(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1848(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1737(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1738(.a(gate287inter0), .b(s_170), .O(gate287inter1));
  and2  gate1739(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1740(.a(s_170), .O(gate287inter3));
  inv1  gate1741(.a(s_171), .O(gate287inter4));
  nand2 gate1742(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1743(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1744(.a(G663), .O(gate287inter7));
  inv1  gate1745(.a(G815), .O(gate287inter8));
  nand2 gate1746(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1747(.a(s_171), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1748(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1749(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1750(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1401(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1402(.a(gate387inter0), .b(s_122), .O(gate387inter1));
  and2  gate1403(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1404(.a(s_122), .O(gate387inter3));
  inv1  gate1405(.a(s_123), .O(gate387inter4));
  nand2 gate1406(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1407(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1408(.a(G1), .O(gate387inter7));
  inv1  gate1409(.a(G1036), .O(gate387inter8));
  nand2 gate1410(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1411(.a(s_123), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1412(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1413(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1414(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1667(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1668(.a(gate394inter0), .b(s_160), .O(gate394inter1));
  and2  gate1669(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1670(.a(s_160), .O(gate394inter3));
  inv1  gate1671(.a(s_161), .O(gate394inter4));
  nand2 gate1672(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1673(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1674(.a(G8), .O(gate394inter7));
  inv1  gate1675(.a(G1057), .O(gate394inter8));
  nand2 gate1676(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1677(.a(s_161), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1678(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1679(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1680(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1933(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1934(.a(gate396inter0), .b(s_198), .O(gate396inter1));
  and2  gate1935(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1936(.a(s_198), .O(gate396inter3));
  inv1  gate1937(.a(s_199), .O(gate396inter4));
  nand2 gate1938(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1939(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1940(.a(G10), .O(gate396inter7));
  inv1  gate1941(.a(G1063), .O(gate396inter8));
  nand2 gate1942(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1943(.a(s_199), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1944(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1945(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1946(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate589(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate590(.a(gate399inter0), .b(s_6), .O(gate399inter1));
  and2  gate591(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate592(.a(s_6), .O(gate399inter3));
  inv1  gate593(.a(s_7), .O(gate399inter4));
  nand2 gate594(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate595(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate596(.a(G13), .O(gate399inter7));
  inv1  gate597(.a(G1072), .O(gate399inter8));
  nand2 gate598(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate599(.a(s_7), .b(gate399inter3), .O(gate399inter10));
  nor2  gate600(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate601(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate602(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1989(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1990(.a(gate402inter0), .b(s_206), .O(gate402inter1));
  and2  gate1991(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1992(.a(s_206), .O(gate402inter3));
  inv1  gate1993(.a(s_207), .O(gate402inter4));
  nand2 gate1994(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1995(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1996(.a(G16), .O(gate402inter7));
  inv1  gate1997(.a(G1081), .O(gate402inter8));
  nand2 gate1998(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1999(.a(s_207), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2000(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2001(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2002(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate701(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate702(.a(gate407inter0), .b(s_22), .O(gate407inter1));
  and2  gate703(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate704(.a(s_22), .O(gate407inter3));
  inv1  gate705(.a(s_23), .O(gate407inter4));
  nand2 gate706(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate707(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate708(.a(G21), .O(gate407inter7));
  inv1  gate709(.a(G1096), .O(gate407inter8));
  nand2 gate710(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate711(.a(s_23), .b(gate407inter3), .O(gate407inter10));
  nor2  gate712(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate713(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate714(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1513(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1514(.a(gate411inter0), .b(s_138), .O(gate411inter1));
  and2  gate1515(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1516(.a(s_138), .O(gate411inter3));
  inv1  gate1517(.a(s_139), .O(gate411inter4));
  nand2 gate1518(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1519(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1520(.a(G25), .O(gate411inter7));
  inv1  gate1521(.a(G1108), .O(gate411inter8));
  nand2 gate1522(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1523(.a(s_139), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1524(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1525(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1526(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate757(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate758(.a(gate415inter0), .b(s_30), .O(gate415inter1));
  and2  gate759(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate760(.a(s_30), .O(gate415inter3));
  inv1  gate761(.a(s_31), .O(gate415inter4));
  nand2 gate762(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate763(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate764(.a(G29), .O(gate415inter7));
  inv1  gate765(.a(G1120), .O(gate415inter8));
  nand2 gate766(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate767(.a(s_31), .b(gate415inter3), .O(gate415inter10));
  nor2  gate768(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate769(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate770(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate953(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate954(.a(gate428inter0), .b(s_58), .O(gate428inter1));
  and2  gate955(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate956(.a(s_58), .O(gate428inter3));
  inv1  gate957(.a(s_59), .O(gate428inter4));
  nand2 gate958(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate959(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate960(.a(G1048), .O(gate428inter7));
  inv1  gate961(.a(G1144), .O(gate428inter8));
  nand2 gate962(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate963(.a(s_59), .b(gate428inter3), .O(gate428inter10));
  nor2  gate964(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate965(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate966(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate729(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate730(.a(gate431inter0), .b(s_26), .O(gate431inter1));
  and2  gate731(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate732(.a(s_26), .O(gate431inter3));
  inv1  gate733(.a(s_27), .O(gate431inter4));
  nand2 gate734(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate735(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate736(.a(G7), .O(gate431inter7));
  inv1  gate737(.a(G1150), .O(gate431inter8));
  nand2 gate738(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate739(.a(s_27), .b(gate431inter3), .O(gate431inter10));
  nor2  gate740(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate741(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate742(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1765(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1766(.a(gate445inter0), .b(s_174), .O(gate445inter1));
  and2  gate1767(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1768(.a(s_174), .O(gate445inter3));
  inv1  gate1769(.a(s_175), .O(gate445inter4));
  nand2 gate1770(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1771(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1772(.a(G14), .O(gate445inter7));
  inv1  gate1773(.a(G1171), .O(gate445inter8));
  nand2 gate1774(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1775(.a(s_175), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1776(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1777(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1778(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1793(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1794(.a(gate455inter0), .b(s_178), .O(gate455inter1));
  and2  gate1795(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1796(.a(s_178), .O(gate455inter3));
  inv1  gate1797(.a(s_179), .O(gate455inter4));
  nand2 gate1798(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1799(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1800(.a(G19), .O(gate455inter7));
  inv1  gate1801(.a(G1186), .O(gate455inter8));
  nand2 gate1802(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1803(.a(s_179), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1804(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1805(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1806(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate645(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate646(.a(gate456inter0), .b(s_14), .O(gate456inter1));
  and2  gate647(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate648(.a(s_14), .O(gate456inter3));
  inv1  gate649(.a(s_15), .O(gate456inter4));
  nand2 gate650(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate651(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate652(.a(G1090), .O(gate456inter7));
  inv1  gate653(.a(G1186), .O(gate456inter8));
  nand2 gate654(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate655(.a(s_15), .b(gate456inter3), .O(gate456inter10));
  nor2  gate656(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate657(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate658(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1289(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1290(.a(gate457inter0), .b(s_106), .O(gate457inter1));
  and2  gate1291(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1292(.a(s_106), .O(gate457inter3));
  inv1  gate1293(.a(s_107), .O(gate457inter4));
  nand2 gate1294(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1295(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1296(.a(G20), .O(gate457inter7));
  inv1  gate1297(.a(G1189), .O(gate457inter8));
  nand2 gate1298(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1299(.a(s_107), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1300(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1301(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1302(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1919(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1920(.a(gate459inter0), .b(s_196), .O(gate459inter1));
  and2  gate1921(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1922(.a(s_196), .O(gate459inter3));
  inv1  gate1923(.a(s_197), .O(gate459inter4));
  nand2 gate1924(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1925(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1926(.a(G21), .O(gate459inter7));
  inv1  gate1927(.a(G1192), .O(gate459inter8));
  nand2 gate1928(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1929(.a(s_197), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1930(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1931(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1932(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate561(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate562(.a(gate464inter0), .b(s_2), .O(gate464inter1));
  and2  gate563(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate564(.a(s_2), .O(gate464inter3));
  inv1  gate565(.a(s_3), .O(gate464inter4));
  nand2 gate566(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate567(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate568(.a(G1102), .O(gate464inter7));
  inv1  gate569(.a(G1198), .O(gate464inter8));
  nand2 gate570(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate571(.a(s_3), .b(gate464inter3), .O(gate464inter10));
  nor2  gate572(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate573(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate574(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1345(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1346(.a(gate465inter0), .b(s_114), .O(gate465inter1));
  and2  gate1347(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1348(.a(s_114), .O(gate465inter3));
  inv1  gate1349(.a(s_115), .O(gate465inter4));
  nand2 gate1350(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1351(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1352(.a(G24), .O(gate465inter7));
  inv1  gate1353(.a(G1201), .O(gate465inter8));
  nand2 gate1354(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1355(.a(s_115), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1356(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1357(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1358(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1443(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1444(.a(gate467inter0), .b(s_128), .O(gate467inter1));
  and2  gate1445(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1446(.a(s_128), .O(gate467inter3));
  inv1  gate1447(.a(s_129), .O(gate467inter4));
  nand2 gate1448(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1449(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1450(.a(G25), .O(gate467inter7));
  inv1  gate1451(.a(G1204), .O(gate467inter8));
  nand2 gate1452(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1453(.a(s_129), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1454(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1455(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1456(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate925(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate926(.a(gate468inter0), .b(s_54), .O(gate468inter1));
  and2  gate927(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate928(.a(s_54), .O(gate468inter3));
  inv1  gate929(.a(s_55), .O(gate468inter4));
  nand2 gate930(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate931(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate932(.a(G1108), .O(gate468inter7));
  inv1  gate933(.a(G1204), .O(gate468inter8));
  nand2 gate934(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate935(.a(s_55), .b(gate468inter3), .O(gate468inter10));
  nor2  gate936(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate937(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate938(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate1877(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1878(.a(gate469inter0), .b(s_190), .O(gate469inter1));
  and2  gate1879(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1880(.a(s_190), .O(gate469inter3));
  inv1  gate1881(.a(s_191), .O(gate469inter4));
  nand2 gate1882(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1883(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1884(.a(G26), .O(gate469inter7));
  inv1  gate1885(.a(G1207), .O(gate469inter8));
  nand2 gate1886(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1887(.a(s_191), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1888(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1889(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1890(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate1807(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1808(.a(gate470inter0), .b(s_180), .O(gate470inter1));
  and2  gate1809(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1810(.a(s_180), .O(gate470inter3));
  inv1  gate1811(.a(s_181), .O(gate470inter4));
  nand2 gate1812(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1813(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1814(.a(G1111), .O(gate470inter7));
  inv1  gate1815(.a(G1207), .O(gate470inter8));
  nand2 gate1816(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1817(.a(s_181), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1818(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1819(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1820(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1065(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1066(.a(gate472inter0), .b(s_74), .O(gate472inter1));
  and2  gate1067(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1068(.a(s_74), .O(gate472inter3));
  inv1  gate1069(.a(s_75), .O(gate472inter4));
  nand2 gate1070(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1071(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1072(.a(G1114), .O(gate472inter7));
  inv1  gate1073(.a(G1210), .O(gate472inter8));
  nand2 gate1074(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1075(.a(s_75), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1076(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1077(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1078(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate939(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate940(.a(gate474inter0), .b(s_56), .O(gate474inter1));
  and2  gate941(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate942(.a(s_56), .O(gate474inter3));
  inv1  gate943(.a(s_57), .O(gate474inter4));
  nand2 gate944(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate945(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate946(.a(G1117), .O(gate474inter7));
  inv1  gate947(.a(G1213), .O(gate474inter8));
  nand2 gate948(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate949(.a(s_57), .b(gate474inter3), .O(gate474inter10));
  nor2  gate950(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate951(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate952(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1709(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1710(.a(gate478inter0), .b(s_166), .O(gate478inter1));
  and2  gate1711(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1712(.a(s_166), .O(gate478inter3));
  inv1  gate1713(.a(s_167), .O(gate478inter4));
  nand2 gate1714(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1715(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1716(.a(G1123), .O(gate478inter7));
  inv1  gate1717(.a(G1219), .O(gate478inter8));
  nand2 gate1718(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1719(.a(s_167), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1720(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1721(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1722(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate827(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate828(.a(gate490inter0), .b(s_40), .O(gate490inter1));
  and2  gate829(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate830(.a(s_40), .O(gate490inter3));
  inv1  gate831(.a(s_41), .O(gate490inter4));
  nand2 gate832(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate833(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate834(.a(G1242), .O(gate490inter7));
  inv1  gate835(.a(G1243), .O(gate490inter8));
  nand2 gate836(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate837(.a(s_41), .b(gate490inter3), .O(gate490inter10));
  nor2  gate838(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate839(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate840(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1177(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1178(.a(gate493inter0), .b(s_90), .O(gate493inter1));
  and2  gate1179(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1180(.a(s_90), .O(gate493inter3));
  inv1  gate1181(.a(s_91), .O(gate493inter4));
  nand2 gate1182(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1183(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1184(.a(G1248), .O(gate493inter7));
  inv1  gate1185(.a(G1249), .O(gate493inter8));
  nand2 gate1186(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1187(.a(s_91), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1188(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1189(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1190(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate617(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate618(.a(gate499inter0), .b(s_10), .O(gate499inter1));
  and2  gate619(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate620(.a(s_10), .O(gate499inter3));
  inv1  gate621(.a(s_11), .O(gate499inter4));
  nand2 gate622(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate623(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate624(.a(G1260), .O(gate499inter7));
  inv1  gate625(.a(G1261), .O(gate499inter8));
  nand2 gate626(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate627(.a(s_11), .b(gate499inter3), .O(gate499inter10));
  nor2  gate628(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate629(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate630(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1695(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1696(.a(gate503inter0), .b(s_164), .O(gate503inter1));
  and2  gate1697(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1698(.a(s_164), .O(gate503inter3));
  inv1  gate1699(.a(s_165), .O(gate503inter4));
  nand2 gate1700(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1701(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1702(.a(G1268), .O(gate503inter7));
  inv1  gate1703(.a(G1269), .O(gate503inter8));
  nand2 gate1704(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1705(.a(s_165), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1706(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1707(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1708(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate673(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate674(.a(gate504inter0), .b(s_18), .O(gate504inter1));
  and2  gate675(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate676(.a(s_18), .O(gate504inter3));
  inv1  gate677(.a(s_19), .O(gate504inter4));
  nand2 gate678(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate679(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate680(.a(G1270), .O(gate504inter7));
  inv1  gate681(.a(G1271), .O(gate504inter8));
  nand2 gate682(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate683(.a(s_19), .b(gate504inter3), .O(gate504inter10));
  nor2  gate684(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate685(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate686(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1219(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1220(.a(gate511inter0), .b(s_96), .O(gate511inter1));
  and2  gate1221(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1222(.a(s_96), .O(gate511inter3));
  inv1  gate1223(.a(s_97), .O(gate511inter4));
  nand2 gate1224(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1225(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1226(.a(G1284), .O(gate511inter7));
  inv1  gate1227(.a(G1285), .O(gate511inter8));
  nand2 gate1228(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1229(.a(s_97), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1230(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1231(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1232(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1681(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1682(.a(gate513inter0), .b(s_162), .O(gate513inter1));
  and2  gate1683(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1684(.a(s_162), .O(gate513inter3));
  inv1  gate1685(.a(s_163), .O(gate513inter4));
  nand2 gate1686(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1687(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1688(.a(G1288), .O(gate513inter7));
  inv1  gate1689(.a(G1289), .O(gate513inter8));
  nand2 gate1690(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1691(.a(s_163), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1692(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1693(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1694(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate967(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate968(.a(gate514inter0), .b(s_60), .O(gate514inter1));
  and2  gate969(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate970(.a(s_60), .O(gate514inter3));
  inv1  gate971(.a(s_61), .O(gate514inter4));
  nand2 gate972(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate973(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate974(.a(G1290), .O(gate514inter7));
  inv1  gate975(.a(G1291), .O(gate514inter8));
  nand2 gate976(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate977(.a(s_61), .b(gate514inter3), .O(gate514inter10));
  nor2  gate978(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate979(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate980(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule