module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1555(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1556(.a(gate12inter0), .b(s_144), .O(gate12inter1));
  and2  gate1557(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1558(.a(s_144), .O(gate12inter3));
  inv1  gate1559(.a(s_145), .O(gate12inter4));
  nand2 gate1560(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1561(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1562(.a(G7), .O(gate12inter7));
  inv1  gate1563(.a(G8), .O(gate12inter8));
  nand2 gate1564(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1565(.a(s_145), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1566(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1567(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1568(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1009(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1010(.a(gate15inter0), .b(s_66), .O(gate15inter1));
  and2  gate1011(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1012(.a(s_66), .O(gate15inter3));
  inv1  gate1013(.a(s_67), .O(gate15inter4));
  nand2 gate1014(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1015(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1016(.a(G13), .O(gate15inter7));
  inv1  gate1017(.a(G14), .O(gate15inter8));
  nand2 gate1018(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1019(.a(s_67), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1020(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1021(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1022(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1345(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1346(.a(gate18inter0), .b(s_114), .O(gate18inter1));
  and2  gate1347(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1348(.a(s_114), .O(gate18inter3));
  inv1  gate1349(.a(s_115), .O(gate18inter4));
  nand2 gate1350(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1351(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1352(.a(G19), .O(gate18inter7));
  inv1  gate1353(.a(G20), .O(gate18inter8));
  nand2 gate1354(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1355(.a(s_115), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1356(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1357(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1358(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate939(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate940(.a(gate21inter0), .b(s_56), .O(gate21inter1));
  and2  gate941(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate942(.a(s_56), .O(gate21inter3));
  inv1  gate943(.a(s_57), .O(gate21inter4));
  nand2 gate944(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate945(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate946(.a(G25), .O(gate21inter7));
  inv1  gate947(.a(G26), .O(gate21inter8));
  nand2 gate948(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate949(.a(s_57), .b(gate21inter3), .O(gate21inter10));
  nor2  gate950(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate951(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate952(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2507(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2508(.a(gate23inter0), .b(s_280), .O(gate23inter1));
  and2  gate2509(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2510(.a(s_280), .O(gate23inter3));
  inv1  gate2511(.a(s_281), .O(gate23inter4));
  nand2 gate2512(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2513(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2514(.a(G29), .O(gate23inter7));
  inv1  gate2515(.a(G30), .O(gate23inter8));
  nand2 gate2516(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2517(.a(s_281), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2518(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2519(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2520(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2045(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2046(.a(gate25inter0), .b(s_214), .O(gate25inter1));
  and2  gate2047(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2048(.a(s_214), .O(gate25inter3));
  inv1  gate2049(.a(s_215), .O(gate25inter4));
  nand2 gate2050(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2051(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2052(.a(G1), .O(gate25inter7));
  inv1  gate2053(.a(G5), .O(gate25inter8));
  nand2 gate2054(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2055(.a(s_215), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2056(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2057(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2058(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1135(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1136(.a(gate26inter0), .b(s_84), .O(gate26inter1));
  and2  gate1137(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1138(.a(s_84), .O(gate26inter3));
  inv1  gate1139(.a(s_85), .O(gate26inter4));
  nand2 gate1140(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1141(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1142(.a(G9), .O(gate26inter7));
  inv1  gate1143(.a(G13), .O(gate26inter8));
  nand2 gate1144(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1145(.a(s_85), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1146(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1147(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1148(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2409(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2410(.a(gate35inter0), .b(s_266), .O(gate35inter1));
  and2  gate2411(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2412(.a(s_266), .O(gate35inter3));
  inv1  gate2413(.a(s_267), .O(gate35inter4));
  nand2 gate2414(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2415(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2416(.a(G18), .O(gate35inter7));
  inv1  gate2417(.a(G22), .O(gate35inter8));
  nand2 gate2418(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2419(.a(s_267), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2420(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2421(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2422(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1191(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1192(.a(gate39inter0), .b(s_92), .O(gate39inter1));
  and2  gate1193(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1194(.a(s_92), .O(gate39inter3));
  inv1  gate1195(.a(s_93), .O(gate39inter4));
  nand2 gate1196(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1197(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1198(.a(G20), .O(gate39inter7));
  inv1  gate1199(.a(G24), .O(gate39inter8));
  nand2 gate1200(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1201(.a(s_93), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1202(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1203(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1204(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1835(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1836(.a(gate42inter0), .b(s_184), .O(gate42inter1));
  and2  gate1837(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1838(.a(s_184), .O(gate42inter3));
  inv1  gate1839(.a(s_185), .O(gate42inter4));
  nand2 gate1840(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1841(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1842(.a(G2), .O(gate42inter7));
  inv1  gate1843(.a(G266), .O(gate42inter8));
  nand2 gate1844(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1845(.a(s_185), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1846(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1847(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1848(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate981(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate982(.a(gate44inter0), .b(s_62), .O(gate44inter1));
  and2  gate983(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate984(.a(s_62), .O(gate44inter3));
  inv1  gate985(.a(s_63), .O(gate44inter4));
  nand2 gate986(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate987(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate988(.a(G4), .O(gate44inter7));
  inv1  gate989(.a(G269), .O(gate44inter8));
  nand2 gate990(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate991(.a(s_63), .b(gate44inter3), .O(gate44inter10));
  nor2  gate992(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate993(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate994(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1667(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1668(.a(gate48inter0), .b(s_160), .O(gate48inter1));
  and2  gate1669(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1670(.a(s_160), .O(gate48inter3));
  inv1  gate1671(.a(s_161), .O(gate48inter4));
  nand2 gate1672(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1673(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1674(.a(G8), .O(gate48inter7));
  inv1  gate1675(.a(G275), .O(gate48inter8));
  nand2 gate1676(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1677(.a(s_161), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1678(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1679(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1680(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1919(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1920(.a(gate54inter0), .b(s_196), .O(gate54inter1));
  and2  gate1921(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1922(.a(s_196), .O(gate54inter3));
  inv1  gate1923(.a(s_197), .O(gate54inter4));
  nand2 gate1924(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1925(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1926(.a(G14), .O(gate54inter7));
  inv1  gate1927(.a(G284), .O(gate54inter8));
  nand2 gate1928(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1929(.a(s_197), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1930(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1931(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1932(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1233(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1234(.a(gate55inter0), .b(s_98), .O(gate55inter1));
  and2  gate1235(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1236(.a(s_98), .O(gate55inter3));
  inv1  gate1237(.a(s_99), .O(gate55inter4));
  nand2 gate1238(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1239(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1240(.a(G15), .O(gate55inter7));
  inv1  gate1241(.a(G287), .O(gate55inter8));
  nand2 gate1242(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1243(.a(s_99), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1244(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1245(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1246(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate897(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate898(.a(gate56inter0), .b(s_50), .O(gate56inter1));
  and2  gate899(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate900(.a(s_50), .O(gate56inter3));
  inv1  gate901(.a(s_51), .O(gate56inter4));
  nand2 gate902(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate903(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate904(.a(G16), .O(gate56inter7));
  inv1  gate905(.a(G287), .O(gate56inter8));
  nand2 gate906(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate907(.a(s_51), .b(gate56inter3), .O(gate56inter10));
  nor2  gate908(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate909(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate910(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1751(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1752(.a(gate58inter0), .b(s_172), .O(gate58inter1));
  and2  gate1753(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1754(.a(s_172), .O(gate58inter3));
  inv1  gate1755(.a(s_173), .O(gate58inter4));
  nand2 gate1756(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1757(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1758(.a(G18), .O(gate58inter7));
  inv1  gate1759(.a(G290), .O(gate58inter8));
  nand2 gate1760(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1761(.a(s_173), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1762(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1763(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1764(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2493(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2494(.a(gate60inter0), .b(s_278), .O(gate60inter1));
  and2  gate2495(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2496(.a(s_278), .O(gate60inter3));
  inv1  gate2497(.a(s_279), .O(gate60inter4));
  nand2 gate2498(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2499(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2500(.a(G20), .O(gate60inter7));
  inv1  gate2501(.a(G293), .O(gate60inter8));
  nand2 gate2502(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2503(.a(s_279), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2504(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2505(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2506(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2129(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2130(.a(gate61inter0), .b(s_226), .O(gate61inter1));
  and2  gate2131(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2132(.a(s_226), .O(gate61inter3));
  inv1  gate2133(.a(s_227), .O(gate61inter4));
  nand2 gate2134(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2135(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2136(.a(G21), .O(gate61inter7));
  inv1  gate2137(.a(G296), .O(gate61inter8));
  nand2 gate2138(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2139(.a(s_227), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2140(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2141(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2142(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2381(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2382(.a(gate62inter0), .b(s_262), .O(gate62inter1));
  and2  gate2383(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2384(.a(s_262), .O(gate62inter3));
  inv1  gate2385(.a(s_263), .O(gate62inter4));
  nand2 gate2386(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2387(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2388(.a(G22), .O(gate62inter7));
  inv1  gate2389(.a(G296), .O(gate62inter8));
  nand2 gate2390(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2391(.a(s_263), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2392(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2393(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2394(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate603(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate604(.a(gate67inter0), .b(s_8), .O(gate67inter1));
  and2  gate605(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate606(.a(s_8), .O(gate67inter3));
  inv1  gate607(.a(s_9), .O(gate67inter4));
  nand2 gate608(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate609(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate610(.a(G27), .O(gate67inter7));
  inv1  gate611(.a(G305), .O(gate67inter8));
  nand2 gate612(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate613(.a(s_9), .b(gate67inter3), .O(gate67inter10));
  nor2  gate614(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate615(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate616(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1709(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1710(.a(gate68inter0), .b(s_166), .O(gate68inter1));
  and2  gate1711(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1712(.a(s_166), .O(gate68inter3));
  inv1  gate1713(.a(s_167), .O(gate68inter4));
  nand2 gate1714(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1715(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1716(.a(G28), .O(gate68inter7));
  inv1  gate1717(.a(G305), .O(gate68inter8));
  nand2 gate1718(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1719(.a(s_167), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1720(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1721(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1722(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate715(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate716(.a(gate70inter0), .b(s_24), .O(gate70inter1));
  and2  gate717(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate718(.a(s_24), .O(gate70inter3));
  inv1  gate719(.a(s_25), .O(gate70inter4));
  nand2 gate720(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate721(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate722(.a(G30), .O(gate70inter7));
  inv1  gate723(.a(G308), .O(gate70inter8));
  nand2 gate724(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate725(.a(s_25), .b(gate70inter3), .O(gate70inter10));
  nor2  gate726(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate727(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate728(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1737(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1738(.a(gate77inter0), .b(s_170), .O(gate77inter1));
  and2  gate1739(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1740(.a(s_170), .O(gate77inter3));
  inv1  gate1741(.a(s_171), .O(gate77inter4));
  nand2 gate1742(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1743(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1744(.a(G2), .O(gate77inter7));
  inv1  gate1745(.a(G320), .O(gate77inter8));
  nand2 gate1746(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1747(.a(s_171), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1748(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1749(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1750(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1863(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1864(.a(gate78inter0), .b(s_188), .O(gate78inter1));
  and2  gate1865(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1866(.a(s_188), .O(gate78inter3));
  inv1  gate1867(.a(s_189), .O(gate78inter4));
  nand2 gate1868(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1869(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1870(.a(G6), .O(gate78inter7));
  inv1  gate1871(.a(G320), .O(gate78inter8));
  nand2 gate1872(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1873(.a(s_189), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1874(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1875(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1876(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1415(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1416(.a(gate79inter0), .b(s_124), .O(gate79inter1));
  and2  gate1417(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1418(.a(s_124), .O(gate79inter3));
  inv1  gate1419(.a(s_125), .O(gate79inter4));
  nand2 gate1420(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1421(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1422(.a(G10), .O(gate79inter7));
  inv1  gate1423(.a(G323), .O(gate79inter8));
  nand2 gate1424(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1425(.a(s_125), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1426(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1427(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1428(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate883(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate884(.a(gate80inter0), .b(s_48), .O(gate80inter1));
  and2  gate885(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate886(.a(s_48), .O(gate80inter3));
  inv1  gate887(.a(s_49), .O(gate80inter4));
  nand2 gate888(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate889(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate890(.a(G14), .O(gate80inter7));
  inv1  gate891(.a(G323), .O(gate80inter8));
  nand2 gate892(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate893(.a(s_49), .b(gate80inter3), .O(gate80inter10));
  nor2  gate894(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate895(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate896(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2549(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2550(.a(gate84inter0), .b(s_286), .O(gate84inter1));
  and2  gate2551(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2552(.a(s_286), .O(gate84inter3));
  inv1  gate2553(.a(s_287), .O(gate84inter4));
  nand2 gate2554(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2555(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2556(.a(G15), .O(gate84inter7));
  inv1  gate2557(.a(G329), .O(gate84inter8));
  nand2 gate2558(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2559(.a(s_287), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2560(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2561(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2562(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1625(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1626(.a(gate85inter0), .b(s_154), .O(gate85inter1));
  and2  gate1627(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1628(.a(s_154), .O(gate85inter3));
  inv1  gate1629(.a(s_155), .O(gate85inter4));
  nand2 gate1630(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1631(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1632(.a(G4), .O(gate85inter7));
  inv1  gate1633(.a(G332), .O(gate85inter8));
  nand2 gate1634(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1635(.a(s_155), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1636(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1637(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1638(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate673(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate674(.a(gate86inter0), .b(s_18), .O(gate86inter1));
  and2  gate675(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate676(.a(s_18), .O(gate86inter3));
  inv1  gate677(.a(s_19), .O(gate86inter4));
  nand2 gate678(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate679(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate680(.a(G8), .O(gate86inter7));
  inv1  gate681(.a(G332), .O(gate86inter8));
  nand2 gate682(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate683(.a(s_19), .b(gate86inter3), .O(gate86inter10));
  nor2  gate684(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate685(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate686(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2577(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2578(.a(gate87inter0), .b(s_290), .O(gate87inter1));
  and2  gate2579(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2580(.a(s_290), .O(gate87inter3));
  inv1  gate2581(.a(s_291), .O(gate87inter4));
  nand2 gate2582(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2583(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2584(.a(G12), .O(gate87inter7));
  inv1  gate2585(.a(G335), .O(gate87inter8));
  nand2 gate2586(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2587(.a(s_291), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2588(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2589(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2590(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1275(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1276(.a(gate89inter0), .b(s_104), .O(gate89inter1));
  and2  gate1277(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1278(.a(s_104), .O(gate89inter3));
  inv1  gate1279(.a(s_105), .O(gate89inter4));
  nand2 gate1280(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1281(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1282(.a(G17), .O(gate89inter7));
  inv1  gate1283(.a(G338), .O(gate89inter8));
  nand2 gate1284(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1285(.a(s_105), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1286(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1287(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1288(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1177(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1178(.a(gate91inter0), .b(s_90), .O(gate91inter1));
  and2  gate1179(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1180(.a(s_90), .O(gate91inter3));
  inv1  gate1181(.a(s_91), .O(gate91inter4));
  nand2 gate1182(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1183(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1184(.a(G25), .O(gate91inter7));
  inv1  gate1185(.a(G341), .O(gate91inter8));
  nand2 gate1186(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1187(.a(s_91), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1188(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1189(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1190(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1289(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1290(.a(gate97inter0), .b(s_106), .O(gate97inter1));
  and2  gate1291(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1292(.a(s_106), .O(gate97inter3));
  inv1  gate1293(.a(s_107), .O(gate97inter4));
  nand2 gate1294(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1295(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1296(.a(G19), .O(gate97inter7));
  inv1  gate1297(.a(G350), .O(gate97inter8));
  nand2 gate1298(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1299(.a(s_107), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1300(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1301(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1302(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1317(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1318(.a(gate106inter0), .b(s_110), .O(gate106inter1));
  and2  gate1319(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1320(.a(s_110), .O(gate106inter3));
  inv1  gate1321(.a(s_111), .O(gate106inter4));
  nand2 gate1322(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1323(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1324(.a(G364), .O(gate106inter7));
  inv1  gate1325(.a(G365), .O(gate106inter8));
  nand2 gate1326(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1327(.a(s_111), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1328(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1329(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1330(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2451(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2452(.a(gate107inter0), .b(s_272), .O(gate107inter1));
  and2  gate2453(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2454(.a(s_272), .O(gate107inter3));
  inv1  gate2455(.a(s_273), .O(gate107inter4));
  nand2 gate2456(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2457(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2458(.a(G366), .O(gate107inter7));
  inv1  gate2459(.a(G367), .O(gate107inter8));
  nand2 gate2460(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2461(.a(s_273), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2462(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2463(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2464(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1583(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1584(.a(gate109inter0), .b(s_148), .O(gate109inter1));
  and2  gate1585(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1586(.a(s_148), .O(gate109inter3));
  inv1  gate1587(.a(s_149), .O(gate109inter4));
  nand2 gate1588(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1589(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1590(.a(G370), .O(gate109inter7));
  inv1  gate1591(.a(G371), .O(gate109inter8));
  nand2 gate1592(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1593(.a(s_149), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1594(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1595(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1596(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate2535(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2536(.a(gate110inter0), .b(s_284), .O(gate110inter1));
  and2  gate2537(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2538(.a(s_284), .O(gate110inter3));
  inv1  gate2539(.a(s_285), .O(gate110inter4));
  nand2 gate2540(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2541(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2542(.a(G372), .O(gate110inter7));
  inv1  gate2543(.a(G373), .O(gate110inter8));
  nand2 gate2544(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2545(.a(s_285), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2546(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2547(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2548(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2591(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2592(.a(gate112inter0), .b(s_292), .O(gate112inter1));
  and2  gate2593(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2594(.a(s_292), .O(gate112inter3));
  inv1  gate2595(.a(s_293), .O(gate112inter4));
  nand2 gate2596(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2597(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2598(.a(G376), .O(gate112inter7));
  inv1  gate2599(.a(G377), .O(gate112inter8));
  nand2 gate2600(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2601(.a(s_293), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2602(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2603(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2604(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate925(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate926(.a(gate113inter0), .b(s_54), .O(gate113inter1));
  and2  gate927(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate928(.a(s_54), .O(gate113inter3));
  inv1  gate929(.a(s_55), .O(gate113inter4));
  nand2 gate930(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate931(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate932(.a(G378), .O(gate113inter7));
  inv1  gate933(.a(G379), .O(gate113inter8));
  nand2 gate934(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate935(.a(s_55), .b(gate113inter3), .O(gate113inter10));
  nor2  gate936(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate937(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate938(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2787(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2788(.a(gate117inter0), .b(s_320), .O(gate117inter1));
  and2  gate2789(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2790(.a(s_320), .O(gate117inter3));
  inv1  gate2791(.a(s_321), .O(gate117inter4));
  nand2 gate2792(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2793(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2794(.a(G386), .O(gate117inter7));
  inv1  gate2795(.a(G387), .O(gate117inter8));
  nand2 gate2796(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2797(.a(s_321), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2798(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2799(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2800(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2367(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2368(.a(gate124inter0), .b(s_260), .O(gate124inter1));
  and2  gate2369(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2370(.a(s_260), .O(gate124inter3));
  inv1  gate2371(.a(s_261), .O(gate124inter4));
  nand2 gate2372(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2373(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2374(.a(G400), .O(gate124inter7));
  inv1  gate2375(.a(G401), .O(gate124inter8));
  nand2 gate2376(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2377(.a(s_261), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2378(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2379(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2380(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate855(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate856(.a(gate126inter0), .b(s_44), .O(gate126inter1));
  and2  gate857(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate858(.a(s_44), .O(gate126inter3));
  inv1  gate859(.a(s_45), .O(gate126inter4));
  nand2 gate860(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate861(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate862(.a(G404), .O(gate126inter7));
  inv1  gate863(.a(G405), .O(gate126inter8));
  nand2 gate864(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate865(.a(s_45), .b(gate126inter3), .O(gate126inter10));
  nor2  gate866(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate867(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate868(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2185(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2186(.a(gate135inter0), .b(s_234), .O(gate135inter1));
  and2  gate2187(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2188(.a(s_234), .O(gate135inter3));
  inv1  gate2189(.a(s_235), .O(gate135inter4));
  nand2 gate2190(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2191(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2192(.a(G422), .O(gate135inter7));
  inv1  gate2193(.a(G423), .O(gate135inter8));
  nand2 gate2194(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2195(.a(s_235), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2196(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2197(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2198(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2241(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2242(.a(gate137inter0), .b(s_242), .O(gate137inter1));
  and2  gate2243(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2244(.a(s_242), .O(gate137inter3));
  inv1  gate2245(.a(s_243), .O(gate137inter4));
  nand2 gate2246(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2247(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2248(.a(G426), .O(gate137inter7));
  inv1  gate2249(.a(G429), .O(gate137inter8));
  nand2 gate2250(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2251(.a(s_243), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2252(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2253(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2254(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1093(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1094(.a(gate139inter0), .b(s_78), .O(gate139inter1));
  and2  gate1095(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1096(.a(s_78), .O(gate139inter3));
  inv1  gate1097(.a(s_79), .O(gate139inter4));
  nand2 gate1098(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1099(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1100(.a(G438), .O(gate139inter7));
  inv1  gate1101(.a(G441), .O(gate139inter8));
  nand2 gate1102(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1103(.a(s_79), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1104(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1105(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1106(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1457(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1458(.a(gate143inter0), .b(s_130), .O(gate143inter1));
  and2  gate1459(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1460(.a(s_130), .O(gate143inter3));
  inv1  gate1461(.a(s_131), .O(gate143inter4));
  nand2 gate1462(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1463(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1464(.a(G462), .O(gate143inter7));
  inv1  gate1465(.a(G465), .O(gate143inter8));
  nand2 gate1466(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1467(.a(s_131), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1468(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1469(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1470(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1359(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1360(.a(gate144inter0), .b(s_116), .O(gate144inter1));
  and2  gate1361(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1362(.a(s_116), .O(gate144inter3));
  inv1  gate1363(.a(s_117), .O(gate144inter4));
  nand2 gate1364(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1365(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1366(.a(G468), .O(gate144inter7));
  inv1  gate1367(.a(G471), .O(gate144inter8));
  nand2 gate1368(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1369(.a(s_117), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1370(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1371(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1372(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1933(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1934(.a(gate145inter0), .b(s_198), .O(gate145inter1));
  and2  gate1935(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1936(.a(s_198), .O(gate145inter3));
  inv1  gate1937(.a(s_199), .O(gate145inter4));
  nand2 gate1938(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1939(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1940(.a(G474), .O(gate145inter7));
  inv1  gate1941(.a(G477), .O(gate145inter8));
  nand2 gate1942(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1943(.a(s_199), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1944(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1945(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1946(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate617(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate618(.a(gate150inter0), .b(s_10), .O(gate150inter1));
  and2  gate619(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate620(.a(s_10), .O(gate150inter3));
  inv1  gate621(.a(s_11), .O(gate150inter4));
  nand2 gate622(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate623(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate624(.a(G504), .O(gate150inter7));
  inv1  gate625(.a(G507), .O(gate150inter8));
  nand2 gate626(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate627(.a(s_11), .b(gate150inter3), .O(gate150inter10));
  nor2  gate628(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate629(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate630(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1639(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1640(.a(gate153inter0), .b(s_156), .O(gate153inter1));
  and2  gate1641(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1642(.a(s_156), .O(gate153inter3));
  inv1  gate1643(.a(s_157), .O(gate153inter4));
  nand2 gate1644(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1645(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1646(.a(G426), .O(gate153inter7));
  inv1  gate1647(.a(G522), .O(gate153inter8));
  nand2 gate1648(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1649(.a(s_157), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1650(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1651(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1652(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1513(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1514(.a(gate154inter0), .b(s_138), .O(gate154inter1));
  and2  gate1515(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1516(.a(s_138), .O(gate154inter3));
  inv1  gate1517(.a(s_139), .O(gate154inter4));
  nand2 gate1518(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1519(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1520(.a(G429), .O(gate154inter7));
  inv1  gate1521(.a(G522), .O(gate154inter8));
  nand2 gate1522(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1523(.a(s_139), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1524(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1525(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1526(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2479(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2480(.a(gate155inter0), .b(s_276), .O(gate155inter1));
  and2  gate2481(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2482(.a(s_276), .O(gate155inter3));
  inv1  gate2483(.a(s_277), .O(gate155inter4));
  nand2 gate2484(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2485(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2486(.a(G432), .O(gate155inter7));
  inv1  gate2487(.a(G525), .O(gate155inter8));
  nand2 gate2488(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2489(.a(s_277), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2490(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2491(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2492(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2759(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2760(.a(gate157inter0), .b(s_316), .O(gate157inter1));
  and2  gate2761(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2762(.a(s_316), .O(gate157inter3));
  inv1  gate2763(.a(s_317), .O(gate157inter4));
  nand2 gate2764(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2765(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2766(.a(G438), .O(gate157inter7));
  inv1  gate2767(.a(G528), .O(gate157inter8));
  nand2 gate2768(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2769(.a(s_317), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2770(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2771(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2772(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2059(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2060(.a(gate159inter0), .b(s_216), .O(gate159inter1));
  and2  gate2061(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2062(.a(s_216), .O(gate159inter3));
  inv1  gate2063(.a(s_217), .O(gate159inter4));
  nand2 gate2064(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2065(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2066(.a(G444), .O(gate159inter7));
  inv1  gate2067(.a(G531), .O(gate159inter8));
  nand2 gate2068(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2069(.a(s_217), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2070(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2071(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2072(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2465(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2466(.a(gate161inter0), .b(s_274), .O(gate161inter1));
  and2  gate2467(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2468(.a(s_274), .O(gate161inter3));
  inv1  gate2469(.a(s_275), .O(gate161inter4));
  nand2 gate2470(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2471(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2472(.a(G450), .O(gate161inter7));
  inv1  gate2473(.a(G534), .O(gate161inter8));
  nand2 gate2474(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2475(.a(s_275), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2476(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2477(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2478(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1569(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1570(.a(gate163inter0), .b(s_146), .O(gate163inter1));
  and2  gate1571(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1572(.a(s_146), .O(gate163inter3));
  inv1  gate1573(.a(s_147), .O(gate163inter4));
  nand2 gate1574(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1575(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1576(.a(G456), .O(gate163inter7));
  inv1  gate1577(.a(G537), .O(gate163inter8));
  nand2 gate1578(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1579(.a(s_147), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1580(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1581(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1582(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1989(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1990(.a(gate165inter0), .b(s_206), .O(gate165inter1));
  and2  gate1991(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1992(.a(s_206), .O(gate165inter3));
  inv1  gate1993(.a(s_207), .O(gate165inter4));
  nand2 gate1994(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1995(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1996(.a(G462), .O(gate165inter7));
  inv1  gate1997(.a(G540), .O(gate165inter8));
  nand2 gate1998(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1999(.a(s_207), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2000(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2001(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2002(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate645(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate646(.a(gate166inter0), .b(s_14), .O(gate166inter1));
  and2  gate647(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate648(.a(s_14), .O(gate166inter3));
  inv1  gate649(.a(s_15), .O(gate166inter4));
  nand2 gate650(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate651(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate652(.a(G465), .O(gate166inter7));
  inv1  gate653(.a(G540), .O(gate166inter8));
  nand2 gate654(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate655(.a(s_15), .b(gate166inter3), .O(gate166inter10));
  nor2  gate656(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate657(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate658(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate967(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate968(.a(gate170inter0), .b(s_60), .O(gate170inter1));
  and2  gate969(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate970(.a(s_60), .O(gate170inter3));
  inv1  gate971(.a(s_61), .O(gate170inter4));
  nand2 gate972(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate973(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate974(.a(G477), .O(gate170inter7));
  inv1  gate975(.a(G546), .O(gate170inter8));
  nand2 gate976(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate977(.a(s_61), .b(gate170inter3), .O(gate170inter10));
  nor2  gate978(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate979(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate980(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1961(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1962(.a(gate175inter0), .b(s_202), .O(gate175inter1));
  and2  gate1963(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1964(.a(s_202), .O(gate175inter3));
  inv1  gate1965(.a(s_203), .O(gate175inter4));
  nand2 gate1966(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1967(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1968(.a(G492), .O(gate175inter7));
  inv1  gate1969(.a(G555), .O(gate175inter8));
  nand2 gate1970(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1971(.a(s_203), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1972(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1973(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1974(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate2773(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2774(.a(gate177inter0), .b(s_318), .O(gate177inter1));
  and2  gate2775(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2776(.a(s_318), .O(gate177inter3));
  inv1  gate2777(.a(s_319), .O(gate177inter4));
  nand2 gate2778(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2779(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2780(.a(G498), .O(gate177inter7));
  inv1  gate2781(.a(G558), .O(gate177inter8));
  nand2 gate2782(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2783(.a(s_319), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2784(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2785(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2786(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2213(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2214(.a(gate180inter0), .b(s_238), .O(gate180inter1));
  and2  gate2215(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2216(.a(s_238), .O(gate180inter3));
  inv1  gate2217(.a(s_239), .O(gate180inter4));
  nand2 gate2218(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2219(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2220(.a(G507), .O(gate180inter7));
  inv1  gate2221(.a(G561), .O(gate180inter8));
  nand2 gate2222(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2223(.a(s_239), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2224(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2225(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2226(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2437(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2438(.a(gate185inter0), .b(s_270), .O(gate185inter1));
  and2  gate2439(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2440(.a(s_270), .O(gate185inter3));
  inv1  gate2441(.a(s_271), .O(gate185inter4));
  nand2 gate2442(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2443(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2444(.a(G570), .O(gate185inter7));
  inv1  gate2445(.a(G571), .O(gate185inter8));
  nand2 gate2446(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2447(.a(s_271), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2448(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2449(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2450(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2339(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2340(.a(gate186inter0), .b(s_256), .O(gate186inter1));
  and2  gate2341(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2342(.a(s_256), .O(gate186inter3));
  inv1  gate2343(.a(s_257), .O(gate186inter4));
  nand2 gate2344(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2345(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2346(.a(G572), .O(gate186inter7));
  inv1  gate2347(.a(G573), .O(gate186inter8));
  nand2 gate2348(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2349(.a(s_257), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2350(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2351(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2352(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1121(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1122(.a(gate187inter0), .b(s_82), .O(gate187inter1));
  and2  gate1123(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1124(.a(s_82), .O(gate187inter3));
  inv1  gate1125(.a(s_83), .O(gate187inter4));
  nand2 gate1126(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1127(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1128(.a(G574), .O(gate187inter7));
  inv1  gate1129(.a(G575), .O(gate187inter8));
  nand2 gate1130(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1131(.a(s_83), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1132(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1133(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1134(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1611(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1612(.a(gate188inter0), .b(s_152), .O(gate188inter1));
  and2  gate1613(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1614(.a(s_152), .O(gate188inter3));
  inv1  gate1615(.a(s_153), .O(gate188inter4));
  nand2 gate1616(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1617(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1618(.a(G576), .O(gate188inter7));
  inv1  gate1619(.a(G577), .O(gate188inter8));
  nand2 gate1620(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1621(.a(s_153), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1622(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1623(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1624(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2563(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2564(.a(gate194inter0), .b(s_288), .O(gate194inter1));
  and2  gate2565(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2566(.a(s_288), .O(gate194inter3));
  inv1  gate2567(.a(s_289), .O(gate194inter4));
  nand2 gate2568(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2569(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2570(.a(G588), .O(gate194inter7));
  inv1  gate2571(.a(G589), .O(gate194inter8));
  nand2 gate2572(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2573(.a(s_289), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2574(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2575(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2576(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate2087(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2088(.a(gate196inter0), .b(s_220), .O(gate196inter1));
  and2  gate2089(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2090(.a(s_220), .O(gate196inter3));
  inv1  gate2091(.a(s_221), .O(gate196inter4));
  nand2 gate2092(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2093(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2094(.a(G592), .O(gate196inter7));
  inv1  gate2095(.a(G593), .O(gate196inter8));
  nand2 gate2096(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2097(.a(s_221), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2098(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2099(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2100(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1247(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1248(.a(gate198inter0), .b(s_100), .O(gate198inter1));
  and2  gate1249(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1250(.a(s_100), .O(gate198inter3));
  inv1  gate1251(.a(s_101), .O(gate198inter4));
  nand2 gate1252(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1253(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1254(.a(G596), .O(gate198inter7));
  inv1  gate1255(.a(G597), .O(gate198inter8));
  nand2 gate1256(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1257(.a(s_101), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1258(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1259(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1260(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1681(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1682(.a(gate201inter0), .b(s_162), .O(gate201inter1));
  and2  gate1683(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1684(.a(s_162), .O(gate201inter3));
  inv1  gate1685(.a(s_163), .O(gate201inter4));
  nand2 gate1686(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1687(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1688(.a(G602), .O(gate201inter7));
  inv1  gate1689(.a(G607), .O(gate201inter8));
  nand2 gate1690(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1691(.a(s_163), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1692(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1693(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1694(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1695(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1696(.a(gate204inter0), .b(s_164), .O(gate204inter1));
  and2  gate1697(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1698(.a(s_164), .O(gate204inter3));
  inv1  gate1699(.a(s_165), .O(gate204inter4));
  nand2 gate1700(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1701(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1702(.a(G607), .O(gate204inter7));
  inv1  gate1703(.a(G617), .O(gate204inter8));
  nand2 gate1704(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1705(.a(s_165), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1706(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1707(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1708(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate841(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate842(.a(gate210inter0), .b(s_42), .O(gate210inter1));
  and2  gate843(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate844(.a(s_42), .O(gate210inter3));
  inv1  gate845(.a(s_43), .O(gate210inter4));
  nand2 gate846(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate847(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate848(.a(G607), .O(gate210inter7));
  inv1  gate849(.a(G666), .O(gate210inter8));
  nand2 gate850(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate851(.a(s_43), .b(gate210inter3), .O(gate210inter10));
  nor2  gate852(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate853(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate854(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1485(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1486(.a(gate212inter0), .b(s_134), .O(gate212inter1));
  and2  gate1487(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1488(.a(s_134), .O(gate212inter3));
  inv1  gate1489(.a(s_135), .O(gate212inter4));
  nand2 gate1490(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1491(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1492(.a(G617), .O(gate212inter7));
  inv1  gate1493(.a(G669), .O(gate212inter8));
  nand2 gate1494(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1495(.a(s_135), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1496(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1497(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1498(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1079(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1080(.a(gate214inter0), .b(s_76), .O(gate214inter1));
  and2  gate1081(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1082(.a(s_76), .O(gate214inter3));
  inv1  gate1083(.a(s_77), .O(gate214inter4));
  nand2 gate1084(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1085(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1086(.a(G612), .O(gate214inter7));
  inv1  gate1087(.a(G672), .O(gate214inter8));
  nand2 gate1088(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1089(.a(s_77), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1090(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1091(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1092(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1429(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1430(.a(gate215inter0), .b(s_126), .O(gate215inter1));
  and2  gate1431(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1432(.a(s_126), .O(gate215inter3));
  inv1  gate1433(.a(s_127), .O(gate215inter4));
  nand2 gate1434(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1435(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1436(.a(G607), .O(gate215inter7));
  inv1  gate1437(.a(G675), .O(gate215inter8));
  nand2 gate1438(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1439(.a(s_127), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1440(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1441(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1442(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate813(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate814(.a(gate221inter0), .b(s_38), .O(gate221inter1));
  and2  gate815(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate816(.a(s_38), .O(gate221inter3));
  inv1  gate817(.a(s_39), .O(gate221inter4));
  nand2 gate818(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate819(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate820(.a(G622), .O(gate221inter7));
  inv1  gate821(.a(G684), .O(gate221inter8));
  nand2 gate822(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate823(.a(s_39), .b(gate221inter3), .O(gate221inter10));
  nor2  gate824(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate825(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate826(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2633(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2634(.a(gate225inter0), .b(s_298), .O(gate225inter1));
  and2  gate2635(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2636(.a(s_298), .O(gate225inter3));
  inv1  gate2637(.a(s_299), .O(gate225inter4));
  nand2 gate2638(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2639(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2640(.a(G690), .O(gate225inter7));
  inv1  gate2641(.a(G691), .O(gate225inter8));
  nand2 gate2642(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2643(.a(s_299), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2644(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2645(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2646(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate659(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate660(.a(gate226inter0), .b(s_16), .O(gate226inter1));
  and2  gate661(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate662(.a(s_16), .O(gate226inter3));
  inv1  gate663(.a(s_17), .O(gate226inter4));
  nand2 gate664(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate665(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate666(.a(G692), .O(gate226inter7));
  inv1  gate667(.a(G693), .O(gate226inter8));
  nand2 gate668(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate669(.a(s_17), .b(gate226inter3), .O(gate226inter10));
  nor2  gate670(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate671(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate672(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate631(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate632(.a(gate232inter0), .b(s_12), .O(gate232inter1));
  and2  gate633(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate634(.a(s_12), .O(gate232inter3));
  inv1  gate635(.a(s_13), .O(gate232inter4));
  nand2 gate636(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate637(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate638(.a(G704), .O(gate232inter7));
  inv1  gate639(.a(G705), .O(gate232inter8));
  nand2 gate640(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate641(.a(s_13), .b(gate232inter3), .O(gate232inter10));
  nor2  gate642(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate643(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate644(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1723(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1724(.a(gate236inter0), .b(s_168), .O(gate236inter1));
  and2  gate1725(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1726(.a(s_168), .O(gate236inter3));
  inv1  gate1727(.a(s_169), .O(gate236inter4));
  nand2 gate1728(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1729(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1730(.a(G251), .O(gate236inter7));
  inv1  gate1731(.a(G727), .O(gate236inter8));
  nand2 gate1732(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1733(.a(s_169), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1734(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1735(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1736(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1261(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1262(.a(gate239inter0), .b(s_102), .O(gate239inter1));
  and2  gate1263(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1264(.a(s_102), .O(gate239inter3));
  inv1  gate1265(.a(s_103), .O(gate239inter4));
  nand2 gate1266(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1267(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1268(.a(G260), .O(gate239inter7));
  inv1  gate1269(.a(G712), .O(gate239inter8));
  nand2 gate1270(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1271(.a(s_103), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1272(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1273(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1274(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2157(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2158(.a(gate244inter0), .b(s_230), .O(gate244inter1));
  and2  gate2159(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2160(.a(s_230), .O(gate244inter3));
  inv1  gate2161(.a(s_231), .O(gate244inter4));
  nand2 gate2162(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2163(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2164(.a(G721), .O(gate244inter7));
  inv1  gate2165(.a(G733), .O(gate244inter8));
  nand2 gate2166(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2167(.a(s_231), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2168(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2169(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2170(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2269(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2270(.a(gate246inter0), .b(s_246), .O(gate246inter1));
  and2  gate2271(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2272(.a(s_246), .O(gate246inter3));
  inv1  gate2273(.a(s_247), .O(gate246inter4));
  nand2 gate2274(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2275(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2276(.a(G724), .O(gate246inter7));
  inv1  gate2277(.a(G736), .O(gate246inter8));
  nand2 gate2278(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2279(.a(s_247), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2280(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2281(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2282(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1877(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1878(.a(gate247inter0), .b(s_190), .O(gate247inter1));
  and2  gate1879(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1880(.a(s_190), .O(gate247inter3));
  inv1  gate1881(.a(s_191), .O(gate247inter4));
  nand2 gate1882(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1883(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1884(.a(G251), .O(gate247inter7));
  inv1  gate1885(.a(G739), .O(gate247inter8));
  nand2 gate1886(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1887(.a(s_191), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1888(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1889(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1890(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2717(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2718(.a(gate248inter0), .b(s_310), .O(gate248inter1));
  and2  gate2719(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2720(.a(s_310), .O(gate248inter3));
  inv1  gate2721(.a(s_311), .O(gate248inter4));
  nand2 gate2722(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2723(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2724(.a(G727), .O(gate248inter7));
  inv1  gate2725(.a(G739), .O(gate248inter8));
  nand2 gate2726(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2727(.a(s_311), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2728(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2729(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2730(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2143(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2144(.a(gate249inter0), .b(s_228), .O(gate249inter1));
  and2  gate2145(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2146(.a(s_228), .O(gate249inter3));
  inv1  gate2147(.a(s_229), .O(gate249inter4));
  nand2 gate2148(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2149(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2150(.a(G254), .O(gate249inter7));
  inv1  gate2151(.a(G742), .O(gate249inter8));
  nand2 gate2152(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2153(.a(s_229), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2154(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2155(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2156(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1205(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1206(.a(gate251inter0), .b(s_94), .O(gate251inter1));
  and2  gate1207(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1208(.a(s_94), .O(gate251inter3));
  inv1  gate1209(.a(s_95), .O(gate251inter4));
  nand2 gate1210(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1211(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1212(.a(G257), .O(gate251inter7));
  inv1  gate1213(.a(G745), .O(gate251inter8));
  nand2 gate1214(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1215(.a(s_95), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1216(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1217(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1218(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2115(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2116(.a(gate254inter0), .b(s_224), .O(gate254inter1));
  and2  gate2117(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2118(.a(s_224), .O(gate254inter3));
  inv1  gate2119(.a(s_225), .O(gate254inter4));
  nand2 gate2120(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2121(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2122(.a(G712), .O(gate254inter7));
  inv1  gate2123(.a(G748), .O(gate254inter8));
  nand2 gate2124(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2125(.a(s_225), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2126(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2127(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2128(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1373(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1374(.a(gate256inter0), .b(s_118), .O(gate256inter1));
  and2  gate1375(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1376(.a(s_118), .O(gate256inter3));
  inv1  gate1377(.a(s_119), .O(gate256inter4));
  nand2 gate1378(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1379(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1380(.a(G715), .O(gate256inter7));
  inv1  gate1381(.a(G751), .O(gate256inter8));
  nand2 gate1382(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1383(.a(s_119), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1384(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1385(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1386(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate743(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate744(.a(gate261inter0), .b(s_28), .O(gate261inter1));
  and2  gate745(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate746(.a(s_28), .O(gate261inter3));
  inv1  gate747(.a(s_29), .O(gate261inter4));
  nand2 gate748(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate749(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate750(.a(G762), .O(gate261inter7));
  inv1  gate751(.a(G763), .O(gate261inter8));
  nand2 gate752(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate753(.a(s_29), .b(gate261inter3), .O(gate261inter10));
  nor2  gate754(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate755(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate756(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate575(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate576(.a(gate265inter0), .b(s_4), .O(gate265inter1));
  and2  gate577(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate578(.a(s_4), .O(gate265inter3));
  inv1  gate579(.a(s_5), .O(gate265inter4));
  nand2 gate580(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate581(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate582(.a(G642), .O(gate265inter7));
  inv1  gate583(.a(G770), .O(gate265inter8));
  nand2 gate584(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate585(.a(s_5), .b(gate265inter3), .O(gate265inter10));
  nor2  gate586(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate587(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate588(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1107(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1108(.a(gate266inter0), .b(s_80), .O(gate266inter1));
  and2  gate1109(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1110(.a(s_80), .O(gate266inter3));
  inv1  gate1111(.a(s_81), .O(gate266inter4));
  nand2 gate1112(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1113(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1114(.a(G645), .O(gate266inter7));
  inv1  gate1115(.a(G773), .O(gate266inter8));
  nand2 gate1116(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1117(.a(s_81), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1118(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1119(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1120(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1947(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1948(.a(gate270inter0), .b(s_200), .O(gate270inter1));
  and2  gate1949(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1950(.a(s_200), .O(gate270inter3));
  inv1  gate1951(.a(s_201), .O(gate270inter4));
  nand2 gate1952(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1953(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1954(.a(G657), .O(gate270inter7));
  inv1  gate1955(.a(G785), .O(gate270inter8));
  nand2 gate1956(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1957(.a(s_201), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1958(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1959(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1960(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2619(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2620(.a(gate272inter0), .b(s_296), .O(gate272inter1));
  and2  gate2621(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2622(.a(s_296), .O(gate272inter3));
  inv1  gate2623(.a(s_297), .O(gate272inter4));
  nand2 gate2624(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2625(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2626(.a(G663), .O(gate272inter7));
  inv1  gate2627(.a(G791), .O(gate272inter8));
  nand2 gate2628(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2629(.a(s_297), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2630(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2631(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2632(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2731(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2732(.a(gate277inter0), .b(s_312), .O(gate277inter1));
  and2  gate2733(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2734(.a(s_312), .O(gate277inter3));
  inv1  gate2735(.a(s_313), .O(gate277inter4));
  nand2 gate2736(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2737(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2738(.a(G648), .O(gate277inter7));
  inv1  gate2739(.a(G800), .O(gate277inter8));
  nand2 gate2740(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2741(.a(s_313), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2742(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2743(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2744(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2395(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2396(.a(gate280inter0), .b(s_264), .O(gate280inter1));
  and2  gate2397(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2398(.a(s_264), .O(gate280inter3));
  inv1  gate2399(.a(s_265), .O(gate280inter4));
  nand2 gate2400(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2401(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2402(.a(G779), .O(gate280inter7));
  inv1  gate2403(.a(G803), .O(gate280inter8));
  nand2 gate2404(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2405(.a(s_265), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2406(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2407(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2408(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2017(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2018(.a(gate282inter0), .b(s_210), .O(gate282inter1));
  and2  gate2019(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2020(.a(s_210), .O(gate282inter3));
  inv1  gate2021(.a(s_211), .O(gate282inter4));
  nand2 gate2022(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2023(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2024(.a(G782), .O(gate282inter7));
  inv1  gate2025(.a(G806), .O(gate282inter8));
  nand2 gate2026(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2027(.a(s_211), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2028(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2029(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2030(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2675(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2676(.a(gate283inter0), .b(s_304), .O(gate283inter1));
  and2  gate2677(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2678(.a(s_304), .O(gate283inter3));
  inv1  gate2679(.a(s_305), .O(gate283inter4));
  nand2 gate2680(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2681(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2682(.a(G657), .O(gate283inter7));
  inv1  gate2683(.a(G809), .O(gate283inter8));
  nand2 gate2684(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2685(.a(s_305), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2686(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2687(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2688(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate589(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate590(.a(gate284inter0), .b(s_6), .O(gate284inter1));
  and2  gate591(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate592(.a(s_6), .O(gate284inter3));
  inv1  gate593(.a(s_7), .O(gate284inter4));
  nand2 gate594(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate595(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate596(.a(G785), .O(gate284inter7));
  inv1  gate597(.a(G809), .O(gate284inter8));
  nand2 gate598(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate599(.a(s_7), .b(gate284inter3), .O(gate284inter10));
  nor2  gate600(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate601(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate602(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1765(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1766(.a(gate285inter0), .b(s_174), .O(gate285inter1));
  and2  gate1767(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1768(.a(s_174), .O(gate285inter3));
  inv1  gate1769(.a(s_175), .O(gate285inter4));
  nand2 gate1770(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1771(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1772(.a(G660), .O(gate285inter7));
  inv1  gate1773(.a(G812), .O(gate285inter8));
  nand2 gate1774(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1775(.a(s_175), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1776(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1777(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1778(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate827(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate828(.a(gate289inter0), .b(s_40), .O(gate289inter1));
  and2  gate829(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate830(.a(s_40), .O(gate289inter3));
  inv1  gate831(.a(s_41), .O(gate289inter4));
  nand2 gate832(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate833(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate834(.a(G818), .O(gate289inter7));
  inv1  gate835(.a(G819), .O(gate289inter8));
  nand2 gate836(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate837(.a(s_41), .b(gate289inter3), .O(gate289inter10));
  nor2  gate838(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate839(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate840(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate2745(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2746(.a(gate290inter0), .b(s_314), .O(gate290inter1));
  and2  gate2747(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2748(.a(s_314), .O(gate290inter3));
  inv1  gate2749(.a(s_315), .O(gate290inter4));
  nand2 gate2750(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2751(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2752(.a(G820), .O(gate290inter7));
  inv1  gate2753(.a(G821), .O(gate290inter8));
  nand2 gate2754(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2755(.a(s_315), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2756(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2757(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2758(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2073(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2074(.a(gate291inter0), .b(s_218), .O(gate291inter1));
  and2  gate2075(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2076(.a(s_218), .O(gate291inter3));
  inv1  gate2077(.a(s_219), .O(gate291inter4));
  nand2 gate2078(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2079(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2080(.a(G822), .O(gate291inter7));
  inv1  gate2081(.a(G823), .O(gate291inter8));
  nand2 gate2082(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2083(.a(s_219), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2084(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2085(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2086(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2283(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2284(.a(gate294inter0), .b(s_248), .O(gate294inter1));
  and2  gate2285(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2286(.a(s_248), .O(gate294inter3));
  inv1  gate2287(.a(s_249), .O(gate294inter4));
  nand2 gate2288(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2289(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2290(.a(G832), .O(gate294inter7));
  inv1  gate2291(.a(G833), .O(gate294inter8));
  nand2 gate2292(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2293(.a(s_249), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2294(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2295(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2296(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1037(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1038(.a(gate295inter0), .b(s_70), .O(gate295inter1));
  and2  gate1039(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1040(.a(s_70), .O(gate295inter3));
  inv1  gate1041(.a(s_71), .O(gate295inter4));
  nand2 gate1042(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1043(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1044(.a(G830), .O(gate295inter7));
  inv1  gate1045(.a(G831), .O(gate295inter8));
  nand2 gate1046(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1047(.a(s_71), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1048(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1049(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1050(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1849(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1850(.a(gate296inter0), .b(s_186), .O(gate296inter1));
  and2  gate1851(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1852(.a(s_186), .O(gate296inter3));
  inv1  gate1853(.a(s_187), .O(gate296inter4));
  nand2 gate1854(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1855(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1856(.a(G826), .O(gate296inter7));
  inv1  gate1857(.a(G827), .O(gate296inter8));
  nand2 gate1858(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1859(.a(s_187), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1860(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1861(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1862(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate785(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate786(.a(gate387inter0), .b(s_34), .O(gate387inter1));
  and2  gate787(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate788(.a(s_34), .O(gate387inter3));
  inv1  gate789(.a(s_35), .O(gate387inter4));
  nand2 gate790(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate791(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate792(.a(G1), .O(gate387inter7));
  inv1  gate793(.a(G1036), .O(gate387inter8));
  nand2 gate794(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate795(.a(s_35), .b(gate387inter3), .O(gate387inter10));
  nor2  gate796(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate797(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate798(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate2605(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2606(.a(gate388inter0), .b(s_294), .O(gate388inter1));
  and2  gate2607(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2608(.a(s_294), .O(gate388inter3));
  inv1  gate2609(.a(s_295), .O(gate388inter4));
  nand2 gate2610(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2611(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2612(.a(G2), .O(gate388inter7));
  inv1  gate2613(.a(G1039), .O(gate388inter8));
  nand2 gate2614(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2615(.a(s_295), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2616(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2617(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2618(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1387(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1388(.a(gate391inter0), .b(s_120), .O(gate391inter1));
  and2  gate1389(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1390(.a(s_120), .O(gate391inter3));
  inv1  gate1391(.a(s_121), .O(gate391inter4));
  nand2 gate1392(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1393(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1394(.a(G5), .O(gate391inter7));
  inv1  gate1395(.a(G1048), .O(gate391inter8));
  nand2 gate1396(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1397(.a(s_121), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1398(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1399(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1400(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate2353(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2354(.a(gate392inter0), .b(s_258), .O(gate392inter1));
  and2  gate2355(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2356(.a(s_258), .O(gate392inter3));
  inv1  gate2357(.a(s_259), .O(gate392inter4));
  nand2 gate2358(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2359(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2360(.a(G6), .O(gate392inter7));
  inv1  gate2361(.a(G1051), .O(gate392inter8));
  nand2 gate2362(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2363(.a(s_259), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2364(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2365(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2366(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1653(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1654(.a(gate394inter0), .b(s_158), .O(gate394inter1));
  and2  gate1655(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1656(.a(s_158), .O(gate394inter3));
  inv1  gate1657(.a(s_159), .O(gate394inter4));
  nand2 gate1658(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1659(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1660(.a(G8), .O(gate394inter7));
  inv1  gate1661(.a(G1057), .O(gate394inter8));
  nand2 gate1662(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1663(.a(s_159), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1664(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1665(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1666(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2423(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2424(.a(gate396inter0), .b(s_268), .O(gate396inter1));
  and2  gate2425(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2426(.a(s_268), .O(gate396inter3));
  inv1  gate2427(.a(s_269), .O(gate396inter4));
  nand2 gate2428(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2429(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2430(.a(G10), .O(gate396inter7));
  inv1  gate2431(.a(G1063), .O(gate396inter8));
  nand2 gate2432(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2433(.a(s_269), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2434(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2435(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2436(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1303(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1304(.a(gate399inter0), .b(s_108), .O(gate399inter1));
  and2  gate1305(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1306(.a(s_108), .O(gate399inter3));
  inv1  gate1307(.a(s_109), .O(gate399inter4));
  nand2 gate1308(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1309(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1310(.a(G13), .O(gate399inter7));
  inv1  gate1311(.a(G1072), .O(gate399inter8));
  nand2 gate1312(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1313(.a(s_109), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1314(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1315(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1316(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1541(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1542(.a(gate407inter0), .b(s_142), .O(gate407inter1));
  and2  gate1543(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1544(.a(s_142), .O(gate407inter3));
  inv1  gate1545(.a(s_143), .O(gate407inter4));
  nand2 gate1546(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1547(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1548(.a(G21), .O(gate407inter7));
  inv1  gate1549(.a(G1096), .O(gate407inter8));
  nand2 gate1550(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1551(.a(s_143), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1552(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1553(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1554(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1471(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1472(.a(gate409inter0), .b(s_132), .O(gate409inter1));
  and2  gate1473(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1474(.a(s_132), .O(gate409inter3));
  inv1  gate1475(.a(s_133), .O(gate409inter4));
  nand2 gate1476(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1477(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1478(.a(G23), .O(gate409inter7));
  inv1  gate1479(.a(G1102), .O(gate409inter8));
  nand2 gate1480(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1481(.a(s_133), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1482(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1483(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1484(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate995(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate996(.a(gate410inter0), .b(s_64), .O(gate410inter1));
  and2  gate997(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate998(.a(s_64), .O(gate410inter3));
  inv1  gate999(.a(s_65), .O(gate410inter4));
  nand2 gate1000(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1001(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1002(.a(G24), .O(gate410inter7));
  inv1  gate1003(.a(G1105), .O(gate410inter8));
  nand2 gate1004(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1005(.a(s_65), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1006(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1007(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1008(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1975(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1976(.a(gate411inter0), .b(s_204), .O(gate411inter1));
  and2  gate1977(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1978(.a(s_204), .O(gate411inter3));
  inv1  gate1979(.a(s_205), .O(gate411inter4));
  nand2 gate1980(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1981(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1982(.a(G25), .O(gate411inter7));
  inv1  gate1983(.a(G1108), .O(gate411inter8));
  nand2 gate1984(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1985(.a(s_205), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1986(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1987(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1988(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1443(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1444(.a(gate412inter0), .b(s_128), .O(gate412inter1));
  and2  gate1445(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1446(.a(s_128), .O(gate412inter3));
  inv1  gate1447(.a(s_129), .O(gate412inter4));
  nand2 gate1448(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1449(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1450(.a(G26), .O(gate412inter7));
  inv1  gate1451(.a(G1111), .O(gate412inter8));
  nand2 gate1452(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1453(.a(s_129), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1454(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1455(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1456(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate771(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate772(.a(gate416inter0), .b(s_32), .O(gate416inter1));
  and2  gate773(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate774(.a(s_32), .O(gate416inter3));
  inv1  gate775(.a(s_33), .O(gate416inter4));
  nand2 gate776(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate777(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate778(.a(G30), .O(gate416inter7));
  inv1  gate779(.a(G1123), .O(gate416inter8));
  nand2 gate780(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate781(.a(s_33), .b(gate416inter3), .O(gate416inter10));
  nor2  gate782(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate783(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate784(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate757(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate758(.a(gate420inter0), .b(s_30), .O(gate420inter1));
  and2  gate759(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate760(.a(s_30), .O(gate420inter3));
  inv1  gate761(.a(s_31), .O(gate420inter4));
  nand2 gate762(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate763(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate764(.a(G1036), .O(gate420inter7));
  inv1  gate765(.a(G1132), .O(gate420inter8));
  nand2 gate766(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate767(.a(s_31), .b(gate420inter3), .O(gate420inter10));
  nor2  gate768(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate769(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate770(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate547(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate548(.a(gate421inter0), .b(s_0), .O(gate421inter1));
  and2  gate549(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate550(.a(s_0), .O(gate421inter3));
  inv1  gate551(.a(s_1), .O(gate421inter4));
  nand2 gate552(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate553(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate554(.a(G2), .O(gate421inter7));
  inv1  gate555(.a(G1135), .O(gate421inter8));
  nand2 gate556(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate557(.a(s_1), .b(gate421inter3), .O(gate421inter10));
  nor2  gate558(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate559(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate560(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2311(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2312(.a(gate423inter0), .b(s_252), .O(gate423inter1));
  and2  gate2313(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2314(.a(s_252), .O(gate423inter3));
  inv1  gate2315(.a(s_253), .O(gate423inter4));
  nand2 gate2316(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2317(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2318(.a(G3), .O(gate423inter7));
  inv1  gate2319(.a(G1138), .O(gate423inter8));
  nand2 gate2320(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2321(.a(s_253), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2322(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2323(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2324(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1401(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1402(.a(gate426inter0), .b(s_122), .O(gate426inter1));
  and2  gate1403(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1404(.a(s_122), .O(gate426inter3));
  inv1  gate1405(.a(s_123), .O(gate426inter4));
  nand2 gate1406(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1407(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1408(.a(G1045), .O(gate426inter7));
  inv1  gate1409(.a(G1141), .O(gate426inter8));
  nand2 gate1410(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1411(.a(s_123), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1412(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1413(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1414(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate953(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate954(.a(gate428inter0), .b(s_58), .O(gate428inter1));
  and2  gate955(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate956(.a(s_58), .O(gate428inter3));
  inv1  gate957(.a(s_59), .O(gate428inter4));
  nand2 gate958(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate959(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate960(.a(G1048), .O(gate428inter7));
  inv1  gate961(.a(G1144), .O(gate428inter8));
  nand2 gate962(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate963(.a(s_59), .b(gate428inter3), .O(gate428inter10));
  nor2  gate964(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate965(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate966(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate561(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate562(.a(gate432inter0), .b(s_2), .O(gate432inter1));
  and2  gate563(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate564(.a(s_2), .O(gate432inter3));
  inv1  gate565(.a(s_3), .O(gate432inter4));
  nand2 gate566(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate567(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate568(.a(G1054), .O(gate432inter7));
  inv1  gate569(.a(G1150), .O(gate432inter8));
  nand2 gate570(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate571(.a(s_3), .b(gate432inter3), .O(gate432inter10));
  nor2  gate572(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate573(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate574(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1499(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1500(.a(gate434inter0), .b(s_136), .O(gate434inter1));
  and2  gate1501(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1502(.a(s_136), .O(gate434inter3));
  inv1  gate1503(.a(s_137), .O(gate434inter4));
  nand2 gate1504(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1505(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1506(.a(G1057), .O(gate434inter7));
  inv1  gate1507(.a(G1153), .O(gate434inter8));
  nand2 gate1508(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1509(.a(s_137), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1510(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1511(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1512(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1331(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1332(.a(gate435inter0), .b(s_112), .O(gate435inter1));
  and2  gate1333(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1334(.a(s_112), .O(gate435inter3));
  inv1  gate1335(.a(s_113), .O(gate435inter4));
  nand2 gate1336(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1337(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1338(.a(G9), .O(gate435inter7));
  inv1  gate1339(.a(G1156), .O(gate435inter8));
  nand2 gate1340(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1341(.a(s_113), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1342(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1343(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1344(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1149(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1150(.a(gate437inter0), .b(s_86), .O(gate437inter1));
  and2  gate1151(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1152(.a(s_86), .O(gate437inter3));
  inv1  gate1153(.a(s_87), .O(gate437inter4));
  nand2 gate1154(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1155(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1156(.a(G10), .O(gate437inter7));
  inv1  gate1157(.a(G1159), .O(gate437inter8));
  nand2 gate1158(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1159(.a(s_87), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1160(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1161(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1162(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2647(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2648(.a(gate440inter0), .b(s_300), .O(gate440inter1));
  and2  gate2649(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2650(.a(s_300), .O(gate440inter3));
  inv1  gate2651(.a(s_301), .O(gate440inter4));
  nand2 gate2652(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2653(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2654(.a(G1066), .O(gate440inter7));
  inv1  gate2655(.a(G1162), .O(gate440inter8));
  nand2 gate2656(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2657(.a(s_301), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2658(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2659(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2660(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1023(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1024(.a(gate442inter0), .b(s_68), .O(gate442inter1));
  and2  gate1025(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1026(.a(s_68), .O(gate442inter3));
  inv1  gate1027(.a(s_69), .O(gate442inter4));
  nand2 gate1028(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1029(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1030(.a(G1069), .O(gate442inter7));
  inv1  gate1031(.a(G1165), .O(gate442inter8));
  nand2 gate1032(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1033(.a(s_69), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1034(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1035(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1036(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate2101(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2102(.a(gate443inter0), .b(s_222), .O(gate443inter1));
  and2  gate2103(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2104(.a(s_222), .O(gate443inter3));
  inv1  gate2105(.a(s_223), .O(gate443inter4));
  nand2 gate2106(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2107(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2108(.a(G13), .O(gate443inter7));
  inv1  gate2109(.a(G1168), .O(gate443inter8));
  nand2 gate2110(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2111(.a(s_223), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2112(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2113(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2114(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate911(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate912(.a(gate444inter0), .b(s_52), .O(gate444inter1));
  and2  gate913(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate914(.a(s_52), .O(gate444inter3));
  inv1  gate915(.a(s_53), .O(gate444inter4));
  nand2 gate916(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate917(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate918(.a(G1072), .O(gate444inter7));
  inv1  gate919(.a(G1168), .O(gate444inter8));
  nand2 gate920(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate921(.a(s_53), .b(gate444inter3), .O(gate444inter10));
  nor2  gate922(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate923(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate924(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate2003(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2004(.a(gate445inter0), .b(s_208), .O(gate445inter1));
  and2  gate2005(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2006(.a(s_208), .O(gate445inter3));
  inv1  gate2007(.a(s_209), .O(gate445inter4));
  nand2 gate2008(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2009(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2010(.a(G14), .O(gate445inter7));
  inv1  gate2011(.a(G1171), .O(gate445inter8));
  nand2 gate2012(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2013(.a(s_209), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2014(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2015(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2016(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1905(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1906(.a(gate448inter0), .b(s_194), .O(gate448inter1));
  and2  gate1907(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1908(.a(s_194), .O(gate448inter3));
  inv1  gate1909(.a(s_195), .O(gate448inter4));
  nand2 gate1910(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1911(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1912(.a(G1078), .O(gate448inter7));
  inv1  gate1913(.a(G1174), .O(gate448inter8));
  nand2 gate1914(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1915(.a(s_195), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1916(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1917(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1918(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate799(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate800(.a(gate449inter0), .b(s_36), .O(gate449inter1));
  and2  gate801(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate802(.a(s_36), .O(gate449inter3));
  inv1  gate803(.a(s_37), .O(gate449inter4));
  nand2 gate804(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate805(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate806(.a(G16), .O(gate449inter7));
  inv1  gate807(.a(G1177), .O(gate449inter8));
  nand2 gate808(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate809(.a(s_37), .b(gate449inter3), .O(gate449inter10));
  nor2  gate810(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate811(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate812(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate2255(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2256(.a(gate450inter0), .b(s_244), .O(gate450inter1));
  and2  gate2257(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2258(.a(s_244), .O(gate450inter3));
  inv1  gate2259(.a(s_245), .O(gate450inter4));
  nand2 gate2260(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2261(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2262(.a(G1081), .O(gate450inter7));
  inv1  gate2263(.a(G1177), .O(gate450inter8));
  nand2 gate2264(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2265(.a(s_245), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2266(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2267(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2268(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2661(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2662(.a(gate451inter0), .b(s_302), .O(gate451inter1));
  and2  gate2663(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2664(.a(s_302), .O(gate451inter3));
  inv1  gate2665(.a(s_303), .O(gate451inter4));
  nand2 gate2666(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2667(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2668(.a(G17), .O(gate451inter7));
  inv1  gate2669(.a(G1180), .O(gate451inter8));
  nand2 gate2670(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2671(.a(s_303), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2672(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2673(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2674(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate2521(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2522(.a(gate452inter0), .b(s_282), .O(gate452inter1));
  and2  gate2523(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2524(.a(s_282), .O(gate452inter3));
  inv1  gate2525(.a(s_283), .O(gate452inter4));
  nand2 gate2526(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2527(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2528(.a(G1084), .O(gate452inter7));
  inv1  gate2529(.a(G1180), .O(gate452inter8));
  nand2 gate2530(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2531(.a(s_283), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2532(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2533(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2534(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate729(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate730(.a(gate453inter0), .b(s_26), .O(gate453inter1));
  and2  gate731(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate732(.a(s_26), .O(gate453inter3));
  inv1  gate733(.a(s_27), .O(gate453inter4));
  nand2 gate734(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate735(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate736(.a(G18), .O(gate453inter7));
  inv1  gate737(.a(G1183), .O(gate453inter8));
  nand2 gate738(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate739(.a(s_27), .b(gate453inter3), .O(gate453inter10));
  nor2  gate740(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate741(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate742(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1597(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1598(.a(gate454inter0), .b(s_150), .O(gate454inter1));
  and2  gate1599(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1600(.a(s_150), .O(gate454inter3));
  inv1  gate1601(.a(s_151), .O(gate454inter4));
  nand2 gate1602(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1603(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1604(.a(G1087), .O(gate454inter7));
  inv1  gate1605(.a(G1183), .O(gate454inter8));
  nand2 gate1606(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1607(.a(s_151), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1608(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1609(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1610(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2297(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2298(.a(gate457inter0), .b(s_250), .O(gate457inter1));
  and2  gate2299(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2300(.a(s_250), .O(gate457inter3));
  inv1  gate2301(.a(s_251), .O(gate457inter4));
  nand2 gate2302(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2303(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2304(.a(G20), .O(gate457inter7));
  inv1  gate2305(.a(G1189), .O(gate457inter8));
  nand2 gate2306(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2307(.a(s_251), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2308(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2309(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2310(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1821(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1822(.a(gate458inter0), .b(s_182), .O(gate458inter1));
  and2  gate1823(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1824(.a(s_182), .O(gate458inter3));
  inv1  gate1825(.a(s_183), .O(gate458inter4));
  nand2 gate1826(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1827(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1828(.a(G1093), .O(gate458inter7));
  inv1  gate1829(.a(G1189), .O(gate458inter8));
  nand2 gate1830(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1831(.a(s_183), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1832(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1833(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1834(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1807(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1808(.a(gate461inter0), .b(s_180), .O(gate461inter1));
  and2  gate1809(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1810(.a(s_180), .O(gate461inter3));
  inv1  gate1811(.a(s_181), .O(gate461inter4));
  nand2 gate1812(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1813(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1814(.a(G22), .O(gate461inter7));
  inv1  gate1815(.a(G1195), .O(gate461inter8));
  nand2 gate1816(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1817(.a(s_181), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1818(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1819(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1820(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2227(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2228(.a(gate463inter0), .b(s_240), .O(gate463inter1));
  and2  gate2229(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2230(.a(s_240), .O(gate463inter3));
  inv1  gate2231(.a(s_241), .O(gate463inter4));
  nand2 gate2232(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2233(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2234(.a(G23), .O(gate463inter7));
  inv1  gate2235(.a(G1198), .O(gate463inter8));
  nand2 gate2236(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2237(.a(s_241), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2238(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2239(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2240(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2325(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2326(.a(gate465inter0), .b(s_254), .O(gate465inter1));
  and2  gate2327(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2328(.a(s_254), .O(gate465inter3));
  inv1  gate2329(.a(s_255), .O(gate465inter4));
  nand2 gate2330(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2331(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2332(.a(G24), .O(gate465inter7));
  inv1  gate2333(.a(G1201), .O(gate465inter8));
  nand2 gate2334(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2335(.a(s_255), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2336(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2337(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2338(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2703(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2704(.a(gate466inter0), .b(s_308), .O(gate466inter1));
  and2  gate2705(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2706(.a(s_308), .O(gate466inter3));
  inv1  gate2707(.a(s_309), .O(gate466inter4));
  nand2 gate2708(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2709(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2710(.a(G1105), .O(gate466inter7));
  inv1  gate2711(.a(G1201), .O(gate466inter8));
  nand2 gate2712(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2713(.a(s_309), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2714(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2715(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2716(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2689(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2690(.a(gate469inter0), .b(s_306), .O(gate469inter1));
  and2  gate2691(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2692(.a(s_306), .O(gate469inter3));
  inv1  gate2693(.a(s_307), .O(gate469inter4));
  nand2 gate2694(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2695(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2696(.a(G26), .O(gate469inter7));
  inv1  gate2697(.a(G1207), .O(gate469inter8));
  nand2 gate2698(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2699(.a(s_307), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2700(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2701(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2702(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1891(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1892(.a(gate471inter0), .b(s_192), .O(gate471inter1));
  and2  gate1893(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1894(.a(s_192), .O(gate471inter3));
  inv1  gate1895(.a(s_193), .O(gate471inter4));
  nand2 gate1896(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1897(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1898(.a(G27), .O(gate471inter7));
  inv1  gate1899(.a(G1210), .O(gate471inter8));
  nand2 gate1900(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1901(.a(s_193), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1902(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1903(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1904(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1051(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1052(.a(gate474inter0), .b(s_72), .O(gate474inter1));
  and2  gate1053(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1054(.a(s_72), .O(gate474inter3));
  inv1  gate1055(.a(s_73), .O(gate474inter4));
  nand2 gate1056(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1057(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1058(.a(G1117), .O(gate474inter7));
  inv1  gate1059(.a(G1213), .O(gate474inter8));
  nand2 gate1060(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1061(.a(s_73), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1062(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1063(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1064(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1527(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1528(.a(gate476inter0), .b(s_140), .O(gate476inter1));
  and2  gate1529(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1530(.a(s_140), .O(gate476inter3));
  inv1  gate1531(.a(s_141), .O(gate476inter4));
  nand2 gate1532(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1533(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1534(.a(G1120), .O(gate476inter7));
  inv1  gate1535(.a(G1216), .O(gate476inter8));
  nand2 gate1536(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1537(.a(s_141), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1538(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1539(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1540(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate869(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate870(.a(gate479inter0), .b(s_46), .O(gate479inter1));
  and2  gate871(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate872(.a(s_46), .O(gate479inter3));
  inv1  gate873(.a(s_47), .O(gate479inter4));
  nand2 gate874(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate875(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate876(.a(G31), .O(gate479inter7));
  inv1  gate877(.a(G1222), .O(gate479inter8));
  nand2 gate878(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate879(.a(s_47), .b(gate479inter3), .O(gate479inter10));
  nor2  gate880(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate881(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate882(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1779(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1780(.a(gate480inter0), .b(s_176), .O(gate480inter1));
  and2  gate1781(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1782(.a(s_176), .O(gate480inter3));
  inv1  gate1783(.a(s_177), .O(gate480inter4));
  nand2 gate1784(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1785(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1786(.a(G1126), .O(gate480inter7));
  inv1  gate1787(.a(G1222), .O(gate480inter8));
  nand2 gate1788(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1789(.a(s_177), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1790(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1791(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1792(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1793(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1794(.a(gate481inter0), .b(s_178), .O(gate481inter1));
  and2  gate1795(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1796(.a(s_178), .O(gate481inter3));
  inv1  gate1797(.a(s_179), .O(gate481inter4));
  nand2 gate1798(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1799(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1800(.a(G32), .O(gate481inter7));
  inv1  gate1801(.a(G1225), .O(gate481inter8));
  nand2 gate1802(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1803(.a(s_179), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1804(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1805(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1806(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2171(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2172(.a(gate483inter0), .b(s_232), .O(gate483inter1));
  and2  gate2173(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2174(.a(s_232), .O(gate483inter3));
  inv1  gate2175(.a(s_233), .O(gate483inter4));
  nand2 gate2176(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2177(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2178(.a(G1228), .O(gate483inter7));
  inv1  gate2179(.a(G1229), .O(gate483inter8));
  nand2 gate2180(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2181(.a(s_233), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2182(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2183(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2184(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1065(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1066(.a(gate487inter0), .b(s_74), .O(gate487inter1));
  and2  gate1067(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1068(.a(s_74), .O(gate487inter3));
  inv1  gate1069(.a(s_75), .O(gate487inter4));
  nand2 gate1070(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1071(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1072(.a(G1236), .O(gate487inter7));
  inv1  gate1073(.a(G1237), .O(gate487inter8));
  nand2 gate1074(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1075(.a(s_75), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1076(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1077(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1078(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate701(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate702(.a(gate499inter0), .b(s_22), .O(gate499inter1));
  and2  gate703(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate704(.a(s_22), .O(gate499inter3));
  inv1  gate705(.a(s_23), .O(gate499inter4));
  nand2 gate706(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate707(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate708(.a(G1260), .O(gate499inter7));
  inv1  gate709(.a(G1261), .O(gate499inter8));
  nand2 gate710(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate711(.a(s_23), .b(gate499inter3), .O(gate499inter10));
  nor2  gate712(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate713(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate714(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1219(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1220(.a(gate502inter0), .b(s_96), .O(gate502inter1));
  and2  gate1221(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1222(.a(s_96), .O(gate502inter3));
  inv1  gate1223(.a(s_97), .O(gate502inter4));
  nand2 gate1224(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1225(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1226(.a(G1266), .O(gate502inter7));
  inv1  gate1227(.a(G1267), .O(gate502inter8));
  nand2 gate1228(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1229(.a(s_97), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1230(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1231(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1232(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate687(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate688(.a(gate504inter0), .b(s_20), .O(gate504inter1));
  and2  gate689(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate690(.a(s_20), .O(gate504inter3));
  inv1  gate691(.a(s_21), .O(gate504inter4));
  nand2 gate692(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate693(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate694(.a(G1270), .O(gate504inter7));
  inv1  gate695(.a(G1271), .O(gate504inter8));
  nand2 gate696(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate697(.a(s_21), .b(gate504inter3), .O(gate504inter10));
  nor2  gate698(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate699(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate700(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2031(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2032(.a(gate508inter0), .b(s_212), .O(gate508inter1));
  and2  gate2033(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2034(.a(s_212), .O(gate508inter3));
  inv1  gate2035(.a(s_213), .O(gate508inter4));
  nand2 gate2036(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2037(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2038(.a(G1278), .O(gate508inter7));
  inv1  gate2039(.a(G1279), .O(gate508inter8));
  nand2 gate2040(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2041(.a(s_213), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2042(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2043(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2044(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2199(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2200(.a(gate510inter0), .b(s_236), .O(gate510inter1));
  and2  gate2201(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2202(.a(s_236), .O(gate510inter3));
  inv1  gate2203(.a(s_237), .O(gate510inter4));
  nand2 gate2204(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2205(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2206(.a(G1282), .O(gate510inter7));
  inv1  gate2207(.a(G1283), .O(gate510inter8));
  nand2 gate2208(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2209(.a(s_237), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2210(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2211(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2212(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1163(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1164(.a(gate513inter0), .b(s_88), .O(gate513inter1));
  and2  gate1165(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1166(.a(s_88), .O(gate513inter3));
  inv1  gate1167(.a(s_89), .O(gate513inter4));
  nand2 gate1168(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1169(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1170(.a(G1288), .O(gate513inter7));
  inv1  gate1171(.a(G1289), .O(gate513inter8));
  nand2 gate1172(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1173(.a(s_89), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1174(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1175(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1176(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule