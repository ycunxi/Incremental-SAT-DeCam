module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate855(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate856(.a(gate9inter0), .b(s_44), .O(gate9inter1));
  and2  gate857(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate858(.a(s_44), .O(gate9inter3));
  inv1  gate859(.a(s_45), .O(gate9inter4));
  nand2 gate860(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate861(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate862(.a(G1), .O(gate9inter7));
  inv1  gate863(.a(G2), .O(gate9inter8));
  nand2 gate864(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate865(.a(s_45), .b(gate9inter3), .O(gate9inter10));
  nor2  gate866(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate867(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate868(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2353(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2354(.a(gate10inter0), .b(s_258), .O(gate10inter1));
  and2  gate2355(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2356(.a(s_258), .O(gate10inter3));
  inv1  gate2357(.a(s_259), .O(gate10inter4));
  nand2 gate2358(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2359(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2360(.a(G3), .O(gate10inter7));
  inv1  gate2361(.a(G4), .O(gate10inter8));
  nand2 gate2362(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2363(.a(s_259), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2364(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2365(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2366(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1149(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1150(.a(gate13inter0), .b(s_86), .O(gate13inter1));
  and2  gate1151(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1152(.a(s_86), .O(gate13inter3));
  inv1  gate1153(.a(s_87), .O(gate13inter4));
  nand2 gate1154(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1155(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1156(.a(G9), .O(gate13inter7));
  inv1  gate1157(.a(G10), .O(gate13inter8));
  nand2 gate1158(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1159(.a(s_87), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1160(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1161(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1162(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2087(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2088(.a(gate17inter0), .b(s_220), .O(gate17inter1));
  and2  gate2089(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2090(.a(s_220), .O(gate17inter3));
  inv1  gate2091(.a(s_221), .O(gate17inter4));
  nand2 gate2092(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2093(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2094(.a(G17), .O(gate17inter7));
  inv1  gate2095(.a(G18), .O(gate17inter8));
  nand2 gate2096(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2097(.a(s_221), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2098(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2099(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2100(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1177(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1178(.a(gate19inter0), .b(s_90), .O(gate19inter1));
  and2  gate1179(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1180(.a(s_90), .O(gate19inter3));
  inv1  gate1181(.a(s_91), .O(gate19inter4));
  nand2 gate1182(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1183(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1184(.a(G21), .O(gate19inter7));
  inv1  gate1185(.a(G22), .O(gate19inter8));
  nand2 gate1186(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1187(.a(s_91), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1188(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1189(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1190(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2017(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2018(.a(gate22inter0), .b(s_210), .O(gate22inter1));
  and2  gate2019(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2020(.a(s_210), .O(gate22inter3));
  inv1  gate2021(.a(s_211), .O(gate22inter4));
  nand2 gate2022(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2023(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2024(.a(G27), .O(gate22inter7));
  inv1  gate2025(.a(G28), .O(gate22inter8));
  nand2 gate2026(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2027(.a(s_211), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2028(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2029(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2030(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1121(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1122(.a(gate25inter0), .b(s_82), .O(gate25inter1));
  and2  gate1123(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1124(.a(s_82), .O(gate25inter3));
  inv1  gate1125(.a(s_83), .O(gate25inter4));
  nand2 gate1126(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1127(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1128(.a(G1), .O(gate25inter7));
  inv1  gate1129(.a(G5), .O(gate25inter8));
  nand2 gate1130(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1131(.a(s_83), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1132(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1133(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1134(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate841(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate842(.a(gate31inter0), .b(s_42), .O(gate31inter1));
  and2  gate843(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate844(.a(s_42), .O(gate31inter3));
  inv1  gate845(.a(s_43), .O(gate31inter4));
  nand2 gate846(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate847(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate848(.a(G4), .O(gate31inter7));
  inv1  gate849(.a(G8), .O(gate31inter8));
  nand2 gate850(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate851(.a(s_43), .b(gate31inter3), .O(gate31inter10));
  nor2  gate852(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate853(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate854(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate981(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate982(.a(gate32inter0), .b(s_62), .O(gate32inter1));
  and2  gate983(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate984(.a(s_62), .O(gate32inter3));
  inv1  gate985(.a(s_63), .O(gate32inter4));
  nand2 gate986(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate987(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate988(.a(G12), .O(gate32inter7));
  inv1  gate989(.a(G16), .O(gate32inter8));
  nand2 gate990(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate991(.a(s_63), .b(gate32inter3), .O(gate32inter10));
  nor2  gate992(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate993(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate994(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate2241(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2242(.a(gate33inter0), .b(s_242), .O(gate33inter1));
  and2  gate2243(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2244(.a(s_242), .O(gate33inter3));
  inv1  gate2245(.a(s_243), .O(gate33inter4));
  nand2 gate2246(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2247(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2248(.a(G17), .O(gate33inter7));
  inv1  gate2249(.a(G21), .O(gate33inter8));
  nand2 gate2250(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2251(.a(s_243), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2252(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2253(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2254(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1387(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1388(.a(gate34inter0), .b(s_120), .O(gate34inter1));
  and2  gate1389(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1390(.a(s_120), .O(gate34inter3));
  inv1  gate1391(.a(s_121), .O(gate34inter4));
  nand2 gate1392(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1393(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1394(.a(G25), .O(gate34inter7));
  inv1  gate1395(.a(G29), .O(gate34inter8));
  nand2 gate1396(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1397(.a(s_121), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1398(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1399(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1400(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate799(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate800(.a(gate41inter0), .b(s_36), .O(gate41inter1));
  and2  gate801(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate802(.a(s_36), .O(gate41inter3));
  inv1  gate803(.a(s_37), .O(gate41inter4));
  nand2 gate804(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate805(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate806(.a(G1), .O(gate41inter7));
  inv1  gate807(.a(G266), .O(gate41inter8));
  nand2 gate808(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate809(.a(s_37), .b(gate41inter3), .O(gate41inter10));
  nor2  gate810(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate811(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate812(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1373(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1374(.a(gate42inter0), .b(s_118), .O(gate42inter1));
  and2  gate1375(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1376(.a(s_118), .O(gate42inter3));
  inv1  gate1377(.a(s_119), .O(gate42inter4));
  nand2 gate1378(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1379(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1380(.a(G2), .O(gate42inter7));
  inv1  gate1381(.a(G266), .O(gate42inter8));
  nand2 gate1382(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1383(.a(s_119), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1384(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1385(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1386(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1247(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1248(.a(gate44inter0), .b(s_100), .O(gate44inter1));
  and2  gate1249(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1250(.a(s_100), .O(gate44inter3));
  inv1  gate1251(.a(s_101), .O(gate44inter4));
  nand2 gate1252(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1253(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1254(.a(G4), .O(gate44inter7));
  inv1  gate1255(.a(G269), .O(gate44inter8));
  nand2 gate1256(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1257(.a(s_101), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1258(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1259(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1260(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1303(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1304(.a(gate45inter0), .b(s_108), .O(gate45inter1));
  and2  gate1305(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1306(.a(s_108), .O(gate45inter3));
  inv1  gate1307(.a(s_109), .O(gate45inter4));
  nand2 gate1308(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1309(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1310(.a(G5), .O(gate45inter7));
  inv1  gate1311(.a(G272), .O(gate45inter8));
  nand2 gate1312(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1313(.a(s_109), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1314(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1315(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1316(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate547(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate548(.a(gate57inter0), .b(s_0), .O(gate57inter1));
  and2  gate549(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate550(.a(s_0), .O(gate57inter3));
  inv1  gate551(.a(s_1), .O(gate57inter4));
  nand2 gate552(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate553(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate554(.a(G17), .O(gate57inter7));
  inv1  gate555(.a(G290), .O(gate57inter8));
  nand2 gate556(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate557(.a(s_1), .b(gate57inter3), .O(gate57inter10));
  nor2  gate558(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate559(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate560(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate645(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate646(.a(gate58inter0), .b(s_14), .O(gate58inter1));
  and2  gate647(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate648(.a(s_14), .O(gate58inter3));
  inv1  gate649(.a(s_15), .O(gate58inter4));
  nand2 gate650(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate651(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate652(.a(G18), .O(gate58inter7));
  inv1  gate653(.a(G290), .O(gate58inter8));
  nand2 gate654(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate655(.a(s_15), .b(gate58inter3), .O(gate58inter10));
  nor2  gate656(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate657(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate658(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2171(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2172(.a(gate60inter0), .b(s_232), .O(gate60inter1));
  and2  gate2173(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2174(.a(s_232), .O(gate60inter3));
  inv1  gate2175(.a(s_233), .O(gate60inter4));
  nand2 gate2176(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2177(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2178(.a(G20), .O(gate60inter7));
  inv1  gate2179(.a(G293), .O(gate60inter8));
  nand2 gate2180(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2181(.a(s_233), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2182(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2183(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2184(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1765(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1766(.a(gate64inter0), .b(s_174), .O(gate64inter1));
  and2  gate1767(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1768(.a(s_174), .O(gate64inter3));
  inv1  gate1769(.a(s_175), .O(gate64inter4));
  nand2 gate1770(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1771(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1772(.a(G24), .O(gate64inter7));
  inv1  gate1773(.a(G299), .O(gate64inter8));
  nand2 gate1774(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1775(.a(s_175), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1776(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1777(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1778(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2535(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2536(.a(gate70inter0), .b(s_284), .O(gate70inter1));
  and2  gate2537(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2538(.a(s_284), .O(gate70inter3));
  inv1  gate2539(.a(s_285), .O(gate70inter4));
  nand2 gate2540(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2541(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2542(.a(G30), .O(gate70inter7));
  inv1  gate2543(.a(G308), .O(gate70inter8));
  nand2 gate2544(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2545(.a(s_285), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2546(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2547(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2548(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1513(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1514(.a(gate75inter0), .b(s_138), .O(gate75inter1));
  and2  gate1515(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1516(.a(s_138), .O(gate75inter3));
  inv1  gate1517(.a(s_139), .O(gate75inter4));
  nand2 gate1518(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1519(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1520(.a(G9), .O(gate75inter7));
  inv1  gate1521(.a(G317), .O(gate75inter8));
  nand2 gate1522(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1523(.a(s_139), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1524(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1525(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1526(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2381(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2382(.a(gate78inter0), .b(s_262), .O(gate78inter1));
  and2  gate2383(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2384(.a(s_262), .O(gate78inter3));
  inv1  gate2385(.a(s_263), .O(gate78inter4));
  nand2 gate2386(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2387(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2388(.a(G6), .O(gate78inter7));
  inv1  gate2389(.a(G320), .O(gate78inter8));
  nand2 gate2390(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2391(.a(s_263), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2392(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2393(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2394(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1961(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1962(.a(gate81inter0), .b(s_202), .O(gate81inter1));
  and2  gate1963(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1964(.a(s_202), .O(gate81inter3));
  inv1  gate1965(.a(s_203), .O(gate81inter4));
  nand2 gate1966(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1967(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1968(.a(G3), .O(gate81inter7));
  inv1  gate1969(.a(G326), .O(gate81inter8));
  nand2 gate1970(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1971(.a(s_203), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1972(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1973(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1974(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate771(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate772(.a(gate82inter0), .b(s_32), .O(gate82inter1));
  and2  gate773(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate774(.a(s_32), .O(gate82inter3));
  inv1  gate775(.a(s_33), .O(gate82inter4));
  nand2 gate776(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate777(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate778(.a(G7), .O(gate82inter7));
  inv1  gate779(.a(G326), .O(gate82inter8));
  nand2 gate780(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate781(.a(s_33), .b(gate82inter3), .O(gate82inter10));
  nor2  gate782(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate783(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate784(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1975(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1976(.a(gate87inter0), .b(s_204), .O(gate87inter1));
  and2  gate1977(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1978(.a(s_204), .O(gate87inter3));
  inv1  gate1979(.a(s_205), .O(gate87inter4));
  nand2 gate1980(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1981(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1982(.a(G12), .O(gate87inter7));
  inv1  gate1983(.a(G335), .O(gate87inter8));
  nand2 gate1984(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1985(.a(s_205), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1986(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1987(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1988(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate2563(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2564(.a(gate88inter0), .b(s_288), .O(gate88inter1));
  and2  gate2565(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2566(.a(s_288), .O(gate88inter3));
  inv1  gate2567(.a(s_289), .O(gate88inter4));
  nand2 gate2568(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2569(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2570(.a(G16), .O(gate88inter7));
  inv1  gate2571(.a(G335), .O(gate88inter8));
  nand2 gate2572(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2573(.a(s_289), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2574(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2575(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2576(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2255(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2256(.a(gate90inter0), .b(s_244), .O(gate90inter1));
  and2  gate2257(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2258(.a(s_244), .O(gate90inter3));
  inv1  gate2259(.a(s_245), .O(gate90inter4));
  nand2 gate2260(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2261(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2262(.a(G21), .O(gate90inter7));
  inv1  gate2263(.a(G338), .O(gate90inter8));
  nand2 gate2264(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2265(.a(s_245), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2266(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2267(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2268(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2003(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2004(.a(gate91inter0), .b(s_208), .O(gate91inter1));
  and2  gate2005(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2006(.a(s_208), .O(gate91inter3));
  inv1  gate2007(.a(s_209), .O(gate91inter4));
  nand2 gate2008(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2009(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2010(.a(G25), .O(gate91inter7));
  inv1  gate2011(.a(G341), .O(gate91inter8));
  nand2 gate2012(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2013(.a(s_209), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2014(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2015(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2016(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2521(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2522(.a(gate94inter0), .b(s_282), .O(gate94inter1));
  and2  gate2523(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2524(.a(s_282), .O(gate94inter3));
  inv1  gate2525(.a(s_283), .O(gate94inter4));
  nand2 gate2526(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2527(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2528(.a(G22), .O(gate94inter7));
  inv1  gate2529(.a(G344), .O(gate94inter8));
  nand2 gate2530(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2531(.a(s_283), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2532(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2533(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2534(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1275(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1276(.a(gate96inter0), .b(s_104), .O(gate96inter1));
  and2  gate1277(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1278(.a(s_104), .O(gate96inter3));
  inv1  gate1279(.a(s_105), .O(gate96inter4));
  nand2 gate1280(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1281(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1282(.a(G30), .O(gate96inter7));
  inv1  gate1283(.a(G347), .O(gate96inter8));
  nand2 gate1284(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1285(.a(s_105), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1286(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1287(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1288(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2199(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2200(.a(gate97inter0), .b(s_236), .O(gate97inter1));
  and2  gate2201(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2202(.a(s_236), .O(gate97inter3));
  inv1  gate2203(.a(s_237), .O(gate97inter4));
  nand2 gate2204(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2205(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2206(.a(G19), .O(gate97inter7));
  inv1  gate2207(.a(G350), .O(gate97inter8));
  nand2 gate2208(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2209(.a(s_237), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2210(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2211(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2212(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1947(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1948(.a(gate100inter0), .b(s_200), .O(gate100inter1));
  and2  gate1949(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1950(.a(s_200), .O(gate100inter3));
  inv1  gate1951(.a(s_201), .O(gate100inter4));
  nand2 gate1952(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1953(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1954(.a(G31), .O(gate100inter7));
  inv1  gate1955(.a(G353), .O(gate100inter8));
  nand2 gate1956(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1957(.a(s_201), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1958(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1959(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1960(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1807(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1808(.a(gate105inter0), .b(s_180), .O(gate105inter1));
  and2  gate1809(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1810(.a(s_180), .O(gate105inter3));
  inv1  gate1811(.a(s_181), .O(gate105inter4));
  nand2 gate1812(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1813(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1814(.a(G362), .O(gate105inter7));
  inv1  gate1815(.a(G363), .O(gate105inter8));
  nand2 gate1816(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1817(.a(s_181), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1818(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1819(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1820(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1527(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1528(.a(gate110inter0), .b(s_140), .O(gate110inter1));
  and2  gate1529(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1530(.a(s_140), .O(gate110inter3));
  inv1  gate1531(.a(s_141), .O(gate110inter4));
  nand2 gate1532(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1533(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1534(.a(G372), .O(gate110inter7));
  inv1  gate1535(.a(G373), .O(gate110inter8));
  nand2 gate1536(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1537(.a(s_141), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1538(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1539(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1540(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1849(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1850(.a(gate112inter0), .b(s_186), .O(gate112inter1));
  and2  gate1851(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1852(.a(s_186), .O(gate112inter3));
  inv1  gate1853(.a(s_187), .O(gate112inter4));
  nand2 gate1854(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1855(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1856(.a(G376), .O(gate112inter7));
  inv1  gate1857(.a(G377), .O(gate112inter8));
  nand2 gate1858(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1859(.a(s_187), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1860(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1861(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1862(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1933(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1934(.a(gate113inter0), .b(s_198), .O(gate113inter1));
  and2  gate1935(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1936(.a(s_198), .O(gate113inter3));
  inv1  gate1937(.a(s_199), .O(gate113inter4));
  nand2 gate1938(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1939(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1940(.a(G378), .O(gate113inter7));
  inv1  gate1941(.a(G379), .O(gate113inter8));
  nand2 gate1942(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1943(.a(s_199), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1944(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1945(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1946(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate659(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate660(.a(gate114inter0), .b(s_16), .O(gate114inter1));
  and2  gate661(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate662(.a(s_16), .O(gate114inter3));
  inv1  gate663(.a(s_17), .O(gate114inter4));
  nand2 gate664(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate665(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate666(.a(G380), .O(gate114inter7));
  inv1  gate667(.a(G381), .O(gate114inter8));
  nand2 gate668(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate669(.a(s_17), .b(gate114inter3), .O(gate114inter10));
  nor2  gate670(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate671(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate672(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2297(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2298(.a(gate116inter0), .b(s_250), .O(gate116inter1));
  and2  gate2299(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2300(.a(s_250), .O(gate116inter3));
  inv1  gate2301(.a(s_251), .O(gate116inter4));
  nand2 gate2302(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2303(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2304(.a(G384), .O(gate116inter7));
  inv1  gate2305(.a(G385), .O(gate116inter8));
  nand2 gate2306(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2307(.a(s_251), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2308(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2309(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2310(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1905(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1906(.a(gate121inter0), .b(s_194), .O(gate121inter1));
  and2  gate1907(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1908(.a(s_194), .O(gate121inter3));
  inv1  gate1909(.a(s_195), .O(gate121inter4));
  nand2 gate1910(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1911(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1912(.a(G394), .O(gate121inter7));
  inv1  gate1913(.a(G395), .O(gate121inter8));
  nand2 gate1914(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1915(.a(s_195), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1916(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1917(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1918(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2395(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2396(.a(gate122inter0), .b(s_264), .O(gate122inter1));
  and2  gate2397(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2398(.a(s_264), .O(gate122inter3));
  inv1  gate2399(.a(s_265), .O(gate122inter4));
  nand2 gate2400(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2401(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2402(.a(G396), .O(gate122inter7));
  inv1  gate2403(.a(G397), .O(gate122inter8));
  nand2 gate2404(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2405(.a(s_265), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2406(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2407(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2408(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1331(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1332(.a(gate125inter0), .b(s_112), .O(gate125inter1));
  and2  gate1333(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1334(.a(s_112), .O(gate125inter3));
  inv1  gate1335(.a(s_113), .O(gate125inter4));
  nand2 gate1336(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1337(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1338(.a(G402), .O(gate125inter7));
  inv1  gate1339(.a(G403), .O(gate125inter8));
  nand2 gate1340(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1341(.a(s_113), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1342(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1343(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1344(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1219(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1220(.a(gate128inter0), .b(s_96), .O(gate128inter1));
  and2  gate1221(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1222(.a(s_96), .O(gate128inter3));
  inv1  gate1223(.a(s_97), .O(gate128inter4));
  nand2 gate1224(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1225(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1226(.a(G408), .O(gate128inter7));
  inv1  gate1227(.a(G409), .O(gate128inter8));
  nand2 gate1228(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1229(.a(s_97), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1230(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1231(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1232(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2423(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2424(.a(gate131inter0), .b(s_268), .O(gate131inter1));
  and2  gate2425(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2426(.a(s_268), .O(gate131inter3));
  inv1  gate2427(.a(s_269), .O(gate131inter4));
  nand2 gate2428(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2429(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2430(.a(G414), .O(gate131inter7));
  inv1  gate2431(.a(G415), .O(gate131inter8));
  nand2 gate2432(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2433(.a(s_269), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2434(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2435(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2436(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1051(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1052(.a(gate132inter0), .b(s_72), .O(gate132inter1));
  and2  gate1053(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1054(.a(s_72), .O(gate132inter3));
  inv1  gate1055(.a(s_73), .O(gate132inter4));
  nand2 gate1056(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1057(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1058(.a(G416), .O(gate132inter7));
  inv1  gate1059(.a(G417), .O(gate132inter8));
  nand2 gate1060(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1061(.a(s_73), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1062(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1063(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1064(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1499(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1500(.a(gate140inter0), .b(s_136), .O(gate140inter1));
  and2  gate1501(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1502(.a(s_136), .O(gate140inter3));
  inv1  gate1503(.a(s_137), .O(gate140inter4));
  nand2 gate1504(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1505(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1506(.a(G444), .O(gate140inter7));
  inv1  gate1507(.a(G447), .O(gate140inter8));
  nand2 gate1508(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1509(.a(s_137), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1510(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1511(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1512(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1863(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1864(.a(gate141inter0), .b(s_188), .O(gate141inter1));
  and2  gate1865(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1866(.a(s_188), .O(gate141inter3));
  inv1  gate1867(.a(s_189), .O(gate141inter4));
  nand2 gate1868(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1869(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1870(.a(G450), .O(gate141inter7));
  inv1  gate1871(.a(G453), .O(gate141inter8));
  nand2 gate1872(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1873(.a(s_189), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1874(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1875(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1876(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate701(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate702(.a(gate142inter0), .b(s_22), .O(gate142inter1));
  and2  gate703(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate704(.a(s_22), .O(gate142inter3));
  inv1  gate705(.a(s_23), .O(gate142inter4));
  nand2 gate706(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate707(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate708(.a(G456), .O(gate142inter7));
  inv1  gate709(.a(G459), .O(gate142inter8));
  nand2 gate710(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate711(.a(s_23), .b(gate142inter3), .O(gate142inter10));
  nor2  gate712(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate713(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate714(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate715(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate716(.a(gate143inter0), .b(s_24), .O(gate143inter1));
  and2  gate717(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate718(.a(s_24), .O(gate143inter3));
  inv1  gate719(.a(s_25), .O(gate143inter4));
  nand2 gate720(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate721(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate722(.a(G462), .O(gate143inter7));
  inv1  gate723(.a(G465), .O(gate143inter8));
  nand2 gate724(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate725(.a(s_25), .b(gate143inter3), .O(gate143inter10));
  nor2  gate726(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate727(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate728(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate589(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate590(.a(gate144inter0), .b(s_6), .O(gate144inter1));
  and2  gate591(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate592(.a(s_6), .O(gate144inter3));
  inv1  gate593(.a(s_7), .O(gate144inter4));
  nand2 gate594(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate595(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate596(.a(G468), .O(gate144inter7));
  inv1  gate597(.a(G471), .O(gate144inter8));
  nand2 gate598(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate599(.a(s_7), .b(gate144inter3), .O(gate144inter10));
  nor2  gate600(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate601(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate602(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate743(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate744(.a(gate145inter0), .b(s_28), .O(gate145inter1));
  and2  gate745(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate746(.a(s_28), .O(gate145inter3));
  inv1  gate747(.a(s_29), .O(gate145inter4));
  nand2 gate748(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate749(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate750(.a(G474), .O(gate145inter7));
  inv1  gate751(.a(G477), .O(gate145inter8));
  nand2 gate752(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate753(.a(s_29), .b(gate145inter3), .O(gate145inter10));
  nor2  gate754(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate755(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate756(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1191(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1192(.a(gate147inter0), .b(s_92), .O(gate147inter1));
  and2  gate1193(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1194(.a(s_92), .O(gate147inter3));
  inv1  gate1195(.a(s_93), .O(gate147inter4));
  nand2 gate1196(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1197(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1198(.a(G486), .O(gate147inter7));
  inv1  gate1199(.a(G489), .O(gate147inter8));
  nand2 gate1200(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1201(.a(s_93), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1202(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1203(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1204(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1555(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1556(.a(gate151inter0), .b(s_144), .O(gate151inter1));
  and2  gate1557(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1558(.a(s_144), .O(gate151inter3));
  inv1  gate1559(.a(s_145), .O(gate151inter4));
  nand2 gate1560(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1561(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1562(.a(G510), .O(gate151inter7));
  inv1  gate1563(.a(G513), .O(gate151inter8));
  nand2 gate1564(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1565(.a(s_145), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1566(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1567(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1568(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2143(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2144(.a(gate152inter0), .b(s_228), .O(gate152inter1));
  and2  gate2145(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2146(.a(s_228), .O(gate152inter3));
  inv1  gate2147(.a(s_229), .O(gate152inter4));
  nand2 gate2148(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2149(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2150(.a(G516), .O(gate152inter7));
  inv1  gate2151(.a(G519), .O(gate152inter8));
  nand2 gate2152(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2153(.a(s_229), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2154(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2155(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2156(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate1737(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1738(.a(gate153inter0), .b(s_170), .O(gate153inter1));
  and2  gate1739(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1740(.a(s_170), .O(gate153inter3));
  inv1  gate1741(.a(s_171), .O(gate153inter4));
  nand2 gate1742(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1743(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1744(.a(G426), .O(gate153inter7));
  inv1  gate1745(.a(G522), .O(gate153inter8));
  nand2 gate1746(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1747(.a(s_171), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1748(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1749(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1750(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2269(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2270(.a(gate157inter0), .b(s_246), .O(gate157inter1));
  and2  gate2271(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2272(.a(s_246), .O(gate157inter3));
  inv1  gate2273(.a(s_247), .O(gate157inter4));
  nand2 gate2274(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2275(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2276(.a(G438), .O(gate157inter7));
  inv1  gate2277(.a(G528), .O(gate157inter8));
  nand2 gate2278(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2279(.a(s_247), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2280(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2281(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2282(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1037(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1038(.a(gate158inter0), .b(s_70), .O(gate158inter1));
  and2  gate1039(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1040(.a(s_70), .O(gate158inter3));
  inv1  gate1041(.a(s_71), .O(gate158inter4));
  nand2 gate1042(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1043(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1044(.a(G441), .O(gate158inter7));
  inv1  gate1045(.a(G528), .O(gate158inter8));
  nand2 gate1046(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1047(.a(s_71), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1048(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1049(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1050(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1415(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1416(.a(gate162inter0), .b(s_124), .O(gate162inter1));
  and2  gate1417(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1418(.a(s_124), .O(gate162inter3));
  inv1  gate1419(.a(s_125), .O(gate162inter4));
  nand2 gate1420(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1421(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1422(.a(G453), .O(gate162inter7));
  inv1  gate1423(.a(G534), .O(gate162inter8));
  nand2 gate1424(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1425(.a(s_125), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1426(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1427(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1428(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate911(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate912(.a(gate164inter0), .b(s_52), .O(gate164inter1));
  and2  gate913(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate914(.a(s_52), .O(gate164inter3));
  inv1  gate915(.a(s_53), .O(gate164inter4));
  nand2 gate916(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate917(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate918(.a(G459), .O(gate164inter7));
  inv1  gate919(.a(G537), .O(gate164inter8));
  nand2 gate920(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate921(.a(s_53), .b(gate164inter3), .O(gate164inter10));
  nor2  gate922(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate923(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate924(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate897(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate898(.a(gate168inter0), .b(s_50), .O(gate168inter1));
  and2  gate899(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate900(.a(s_50), .O(gate168inter3));
  inv1  gate901(.a(s_51), .O(gate168inter4));
  nand2 gate902(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate903(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate904(.a(G471), .O(gate168inter7));
  inv1  gate905(.a(G543), .O(gate168inter8));
  nand2 gate906(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate907(.a(s_51), .b(gate168inter3), .O(gate168inter10));
  nor2  gate908(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate909(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate910(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1429(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1430(.a(gate169inter0), .b(s_126), .O(gate169inter1));
  and2  gate1431(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1432(.a(s_126), .O(gate169inter3));
  inv1  gate1433(.a(s_127), .O(gate169inter4));
  nand2 gate1434(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1435(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1436(.a(G474), .O(gate169inter7));
  inv1  gate1437(.a(G546), .O(gate169inter8));
  nand2 gate1438(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1439(.a(s_127), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1440(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1441(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1442(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1709(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1710(.a(gate173inter0), .b(s_166), .O(gate173inter1));
  and2  gate1711(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1712(.a(s_166), .O(gate173inter3));
  inv1  gate1713(.a(s_167), .O(gate173inter4));
  nand2 gate1714(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1715(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1716(.a(G486), .O(gate173inter7));
  inv1  gate1717(.a(G552), .O(gate173inter8));
  nand2 gate1718(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1719(.a(s_167), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1720(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1721(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1722(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1093(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1094(.a(gate175inter0), .b(s_78), .O(gate175inter1));
  and2  gate1095(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1096(.a(s_78), .O(gate175inter3));
  inv1  gate1097(.a(s_79), .O(gate175inter4));
  nand2 gate1098(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1099(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1100(.a(G492), .O(gate175inter7));
  inv1  gate1101(.a(G555), .O(gate175inter8));
  nand2 gate1102(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1103(.a(s_79), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1104(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1105(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1106(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate673(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate674(.a(gate183inter0), .b(s_18), .O(gate183inter1));
  and2  gate675(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate676(.a(s_18), .O(gate183inter3));
  inv1  gate677(.a(s_19), .O(gate183inter4));
  nand2 gate678(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate679(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate680(.a(G516), .O(gate183inter7));
  inv1  gate681(.a(G567), .O(gate183inter8));
  nand2 gate682(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate683(.a(s_19), .b(gate183inter3), .O(gate183inter10));
  nor2  gate684(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate685(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate686(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2507(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2508(.a(gate188inter0), .b(s_280), .O(gate188inter1));
  and2  gate2509(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2510(.a(s_280), .O(gate188inter3));
  inv1  gate2511(.a(s_281), .O(gate188inter4));
  nand2 gate2512(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2513(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2514(.a(G576), .O(gate188inter7));
  inv1  gate2515(.a(G577), .O(gate188inter8));
  nand2 gate2516(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2517(.a(s_281), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2518(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2519(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2520(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1695(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1696(.a(gate189inter0), .b(s_164), .O(gate189inter1));
  and2  gate1697(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1698(.a(s_164), .O(gate189inter3));
  inv1  gate1699(.a(s_165), .O(gate189inter4));
  nand2 gate1700(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1701(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1702(.a(G578), .O(gate189inter7));
  inv1  gate1703(.a(G579), .O(gate189inter8));
  nand2 gate1704(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1705(.a(s_165), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1706(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1707(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1708(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate953(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate954(.a(gate192inter0), .b(s_58), .O(gate192inter1));
  and2  gate955(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate956(.a(s_58), .O(gate192inter3));
  inv1  gate957(.a(s_59), .O(gate192inter4));
  nand2 gate958(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate959(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate960(.a(G584), .O(gate192inter7));
  inv1  gate961(.a(G585), .O(gate192inter8));
  nand2 gate962(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate963(.a(s_59), .b(gate192inter3), .O(gate192inter10));
  nor2  gate964(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate965(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate966(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1611(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1612(.a(gate195inter0), .b(s_152), .O(gate195inter1));
  and2  gate1613(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1614(.a(s_152), .O(gate195inter3));
  inv1  gate1615(.a(s_153), .O(gate195inter4));
  nand2 gate1616(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1617(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1618(.a(G590), .O(gate195inter7));
  inv1  gate1619(.a(G591), .O(gate195inter8));
  nand2 gate1620(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1621(.a(s_153), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1622(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1623(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1624(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1541(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1542(.a(gate202inter0), .b(s_142), .O(gate202inter1));
  and2  gate1543(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1544(.a(s_142), .O(gate202inter3));
  inv1  gate1545(.a(s_143), .O(gate202inter4));
  nand2 gate1546(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1547(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1548(.a(G612), .O(gate202inter7));
  inv1  gate1549(.a(G617), .O(gate202inter8));
  nand2 gate1550(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1551(.a(s_143), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1552(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1553(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1554(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate2437(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2438(.a(gate203inter0), .b(s_270), .O(gate203inter1));
  and2  gate2439(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2440(.a(s_270), .O(gate203inter3));
  inv1  gate2441(.a(s_271), .O(gate203inter4));
  nand2 gate2442(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2443(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2444(.a(G602), .O(gate203inter7));
  inv1  gate2445(.a(G612), .O(gate203inter8));
  nand2 gate2446(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2447(.a(s_271), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2448(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2449(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2450(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2493(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2494(.a(gate208inter0), .b(s_278), .O(gate208inter1));
  and2  gate2495(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2496(.a(s_278), .O(gate208inter3));
  inv1  gate2497(.a(s_279), .O(gate208inter4));
  nand2 gate2498(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2499(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2500(.a(G627), .O(gate208inter7));
  inv1  gate2501(.a(G637), .O(gate208inter8));
  nand2 gate2502(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2503(.a(s_279), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2504(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2505(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2506(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1443(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1444(.a(gate213inter0), .b(s_128), .O(gate213inter1));
  and2  gate1445(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1446(.a(s_128), .O(gate213inter3));
  inv1  gate1447(.a(s_129), .O(gate213inter4));
  nand2 gate1448(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1449(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1450(.a(G602), .O(gate213inter7));
  inv1  gate1451(.a(G672), .O(gate213inter8));
  nand2 gate1452(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1453(.a(s_129), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1454(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1455(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1456(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1793(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1794(.a(gate215inter0), .b(s_178), .O(gate215inter1));
  and2  gate1795(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1796(.a(s_178), .O(gate215inter3));
  inv1  gate1797(.a(s_179), .O(gate215inter4));
  nand2 gate1798(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1799(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1800(.a(G607), .O(gate215inter7));
  inv1  gate1801(.a(G675), .O(gate215inter8));
  nand2 gate1802(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1803(.a(s_179), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1804(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1805(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1806(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1583(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1584(.a(gate216inter0), .b(s_148), .O(gate216inter1));
  and2  gate1585(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1586(.a(s_148), .O(gate216inter3));
  inv1  gate1587(.a(s_149), .O(gate216inter4));
  nand2 gate1588(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1589(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1590(.a(G617), .O(gate216inter7));
  inv1  gate1591(.a(G675), .O(gate216inter8));
  nand2 gate1592(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1593(.a(s_149), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1594(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1595(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1596(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1653(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1654(.a(gate218inter0), .b(s_158), .O(gate218inter1));
  and2  gate1655(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1656(.a(s_158), .O(gate218inter3));
  inv1  gate1657(.a(s_159), .O(gate218inter4));
  nand2 gate1658(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1659(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1660(.a(G627), .O(gate218inter7));
  inv1  gate1661(.a(G678), .O(gate218inter8));
  nand2 gate1662(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1663(.a(s_159), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1664(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1665(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1666(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate2367(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2368(.a(gate221inter0), .b(s_260), .O(gate221inter1));
  and2  gate2369(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2370(.a(s_260), .O(gate221inter3));
  inv1  gate2371(.a(s_261), .O(gate221inter4));
  nand2 gate2372(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2373(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2374(.a(G622), .O(gate221inter7));
  inv1  gate2375(.a(G684), .O(gate221inter8));
  nand2 gate2376(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2377(.a(s_261), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2378(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2379(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2380(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate687(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate688(.a(gate229inter0), .b(s_20), .O(gate229inter1));
  and2  gate689(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate690(.a(s_20), .O(gate229inter3));
  inv1  gate691(.a(s_21), .O(gate229inter4));
  nand2 gate692(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate693(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate694(.a(G698), .O(gate229inter7));
  inv1  gate695(.a(G699), .O(gate229inter8));
  nand2 gate696(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate697(.a(s_21), .b(gate229inter3), .O(gate229inter10));
  nor2  gate698(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate699(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate700(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate883(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate884(.a(gate232inter0), .b(s_48), .O(gate232inter1));
  and2  gate885(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate886(.a(s_48), .O(gate232inter3));
  inv1  gate887(.a(s_49), .O(gate232inter4));
  nand2 gate888(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate889(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate890(.a(G704), .O(gate232inter7));
  inv1  gate891(.a(G705), .O(gate232inter8));
  nand2 gate892(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate893(.a(s_49), .b(gate232inter3), .O(gate232inter10));
  nor2  gate894(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate895(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate896(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1877(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1878(.a(gate235inter0), .b(s_190), .O(gate235inter1));
  and2  gate1879(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1880(.a(s_190), .O(gate235inter3));
  inv1  gate1881(.a(s_191), .O(gate235inter4));
  nand2 gate1882(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1883(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1884(.a(G248), .O(gate235inter7));
  inv1  gate1885(.a(G724), .O(gate235inter8));
  nand2 gate1886(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1887(.a(s_191), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1888(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1889(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1890(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1835(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1836(.a(gate237inter0), .b(s_184), .O(gate237inter1));
  and2  gate1837(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1838(.a(s_184), .O(gate237inter3));
  inv1  gate1839(.a(s_185), .O(gate237inter4));
  nand2 gate1840(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1841(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1842(.a(G254), .O(gate237inter7));
  inv1  gate1843(.a(G706), .O(gate237inter8));
  nand2 gate1844(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1845(.a(s_185), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1846(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1847(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1848(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate603(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate604(.a(gate243inter0), .b(s_8), .O(gate243inter1));
  and2  gate605(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate606(.a(s_8), .O(gate243inter3));
  inv1  gate607(.a(s_9), .O(gate243inter4));
  nand2 gate608(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate609(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate610(.a(G245), .O(gate243inter7));
  inv1  gate611(.a(G733), .O(gate243inter8));
  nand2 gate612(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate613(.a(s_9), .b(gate243inter3), .O(gate243inter10));
  nor2  gate614(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate615(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate616(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1009(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1010(.a(gate245inter0), .b(s_66), .O(gate245inter1));
  and2  gate1011(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1012(.a(s_66), .O(gate245inter3));
  inv1  gate1013(.a(s_67), .O(gate245inter4));
  nand2 gate1014(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1015(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1016(.a(G248), .O(gate245inter7));
  inv1  gate1017(.a(G736), .O(gate245inter8));
  nand2 gate1018(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1019(.a(s_67), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1020(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1021(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1022(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate785(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate786(.a(gate248inter0), .b(s_34), .O(gate248inter1));
  and2  gate787(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate788(.a(s_34), .O(gate248inter3));
  inv1  gate789(.a(s_35), .O(gate248inter4));
  nand2 gate790(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate791(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate792(.a(G727), .O(gate248inter7));
  inv1  gate793(.a(G739), .O(gate248inter8));
  nand2 gate794(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate795(.a(s_35), .b(gate248inter3), .O(gate248inter10));
  nor2  gate796(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate797(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate798(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate575(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate576(.a(gate249inter0), .b(s_4), .O(gate249inter1));
  and2  gate577(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate578(.a(s_4), .O(gate249inter3));
  inv1  gate579(.a(s_5), .O(gate249inter4));
  nand2 gate580(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate581(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate582(.a(G254), .O(gate249inter7));
  inv1  gate583(.a(G742), .O(gate249inter8));
  nand2 gate584(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate585(.a(s_5), .b(gate249inter3), .O(gate249inter10));
  nor2  gate586(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate587(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate588(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate995(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate996(.a(gate252inter0), .b(s_64), .O(gate252inter1));
  and2  gate997(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate998(.a(s_64), .O(gate252inter3));
  inv1  gate999(.a(s_65), .O(gate252inter4));
  nand2 gate1000(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1001(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1002(.a(G709), .O(gate252inter7));
  inv1  gate1003(.a(G745), .O(gate252inter8));
  nand2 gate1004(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1005(.a(s_65), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1006(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1007(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1008(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate2479(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2480(.a(gate253inter0), .b(s_276), .O(gate253inter1));
  and2  gate2481(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2482(.a(s_276), .O(gate253inter3));
  inv1  gate2483(.a(s_277), .O(gate253inter4));
  nand2 gate2484(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2485(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2486(.a(G260), .O(gate253inter7));
  inv1  gate2487(.a(G748), .O(gate253inter8));
  nand2 gate2488(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2489(.a(s_277), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2490(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2491(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2492(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate2185(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2186(.a(gate254inter0), .b(s_234), .O(gate254inter1));
  and2  gate2187(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2188(.a(s_234), .O(gate254inter3));
  inv1  gate2189(.a(s_235), .O(gate254inter4));
  nand2 gate2190(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2191(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2192(.a(G712), .O(gate254inter7));
  inv1  gate2193(.a(G748), .O(gate254inter8));
  nand2 gate2194(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2195(.a(s_235), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2196(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2197(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2198(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate2031(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2032(.a(gate255inter0), .b(s_212), .O(gate255inter1));
  and2  gate2033(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2034(.a(s_212), .O(gate255inter3));
  inv1  gate2035(.a(s_213), .O(gate255inter4));
  nand2 gate2036(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2037(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2038(.a(G263), .O(gate255inter7));
  inv1  gate2039(.a(G751), .O(gate255inter8));
  nand2 gate2040(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2041(.a(s_213), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2042(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2043(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2044(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2073(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2074(.a(gate258inter0), .b(s_218), .O(gate258inter1));
  and2  gate2075(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2076(.a(s_218), .O(gate258inter3));
  inv1  gate2077(.a(s_219), .O(gate258inter4));
  nand2 gate2078(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2079(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2080(.a(G756), .O(gate258inter7));
  inv1  gate2081(.a(G757), .O(gate258inter8));
  nand2 gate2082(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2083(.a(s_219), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2084(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2085(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2086(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1261(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1262(.a(gate259inter0), .b(s_102), .O(gate259inter1));
  and2  gate1263(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1264(.a(s_102), .O(gate259inter3));
  inv1  gate1265(.a(s_103), .O(gate259inter4));
  nand2 gate1266(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1267(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1268(.a(G758), .O(gate259inter7));
  inv1  gate1269(.a(G759), .O(gate259inter8));
  nand2 gate1270(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1271(.a(s_103), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1272(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1273(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1274(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1079(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1080(.a(gate261inter0), .b(s_76), .O(gate261inter1));
  and2  gate1081(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1082(.a(s_76), .O(gate261inter3));
  inv1  gate1083(.a(s_77), .O(gate261inter4));
  nand2 gate1084(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1085(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1086(.a(G762), .O(gate261inter7));
  inv1  gate1087(.a(G763), .O(gate261inter8));
  nand2 gate1088(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1089(.a(s_77), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1090(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1091(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1092(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate925(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate926(.a(gate266inter0), .b(s_54), .O(gate266inter1));
  and2  gate927(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate928(.a(s_54), .O(gate266inter3));
  inv1  gate929(.a(s_55), .O(gate266inter4));
  nand2 gate930(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate931(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate932(.a(G645), .O(gate266inter7));
  inv1  gate933(.a(G773), .O(gate266inter8));
  nand2 gate934(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate935(.a(s_55), .b(gate266inter3), .O(gate266inter10));
  nor2  gate936(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate937(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate938(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate561(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate562(.a(gate270inter0), .b(s_2), .O(gate270inter1));
  and2  gate563(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate564(.a(s_2), .O(gate270inter3));
  inv1  gate565(.a(s_3), .O(gate270inter4));
  nand2 gate566(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate567(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate568(.a(G657), .O(gate270inter7));
  inv1  gate569(.a(G785), .O(gate270inter8));
  nand2 gate570(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate571(.a(s_3), .b(gate270inter3), .O(gate270inter10));
  nor2  gate572(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate573(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate574(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2325(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2326(.a(gate271inter0), .b(s_254), .O(gate271inter1));
  and2  gate2327(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2328(.a(s_254), .O(gate271inter3));
  inv1  gate2329(.a(s_255), .O(gate271inter4));
  nand2 gate2330(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2331(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2332(.a(G660), .O(gate271inter7));
  inv1  gate2333(.a(G788), .O(gate271inter8));
  nand2 gate2334(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2335(.a(s_255), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2336(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2337(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2338(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2283(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2284(.a(gate272inter0), .b(s_248), .O(gate272inter1));
  and2  gate2285(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2286(.a(s_248), .O(gate272inter3));
  inv1  gate2287(.a(s_249), .O(gate272inter4));
  nand2 gate2288(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2289(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2290(.a(G663), .O(gate272inter7));
  inv1  gate2291(.a(G791), .O(gate272inter8));
  nand2 gate2292(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2293(.a(s_249), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2294(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2295(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2296(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1205(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1206(.a(gate273inter0), .b(s_94), .O(gate273inter1));
  and2  gate1207(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1208(.a(s_94), .O(gate273inter3));
  inv1  gate1209(.a(s_95), .O(gate273inter4));
  nand2 gate1210(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1211(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1212(.a(G642), .O(gate273inter7));
  inv1  gate1213(.a(G794), .O(gate273inter8));
  nand2 gate1214(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1215(.a(s_95), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1216(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1217(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1218(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1471(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1472(.a(gate274inter0), .b(s_132), .O(gate274inter1));
  and2  gate1473(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1474(.a(s_132), .O(gate274inter3));
  inv1  gate1475(.a(s_133), .O(gate274inter4));
  nand2 gate1476(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1477(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1478(.a(G770), .O(gate274inter7));
  inv1  gate1479(.a(G794), .O(gate274inter8));
  nand2 gate1480(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1481(.a(s_133), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1482(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1483(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1484(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1821(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1822(.a(gate277inter0), .b(s_182), .O(gate277inter1));
  and2  gate1823(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1824(.a(s_182), .O(gate277inter3));
  inv1  gate1825(.a(s_183), .O(gate277inter4));
  nand2 gate1826(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1827(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1828(.a(G648), .O(gate277inter7));
  inv1  gate1829(.a(G800), .O(gate277inter8));
  nand2 gate1830(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1831(.a(s_183), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1832(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1833(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1834(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1569(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1570(.a(gate285inter0), .b(s_146), .O(gate285inter1));
  and2  gate1571(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1572(.a(s_146), .O(gate285inter3));
  inv1  gate1573(.a(s_147), .O(gate285inter4));
  nand2 gate1574(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1575(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1576(.a(G660), .O(gate285inter7));
  inv1  gate1577(.a(G812), .O(gate285inter8));
  nand2 gate1578(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1579(.a(s_147), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1580(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1581(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1582(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1345(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1346(.a(gate294inter0), .b(s_114), .O(gate294inter1));
  and2  gate1347(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1348(.a(s_114), .O(gate294inter3));
  inv1  gate1349(.a(s_115), .O(gate294inter4));
  nand2 gate1350(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1351(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1352(.a(G832), .O(gate294inter7));
  inv1  gate1353(.a(G833), .O(gate294inter8));
  nand2 gate1354(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1355(.a(s_115), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1356(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1357(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1358(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1751(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1752(.a(gate389inter0), .b(s_172), .O(gate389inter1));
  and2  gate1753(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1754(.a(s_172), .O(gate389inter3));
  inv1  gate1755(.a(s_173), .O(gate389inter4));
  nand2 gate1756(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1757(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1758(.a(G3), .O(gate389inter7));
  inv1  gate1759(.a(G1042), .O(gate389inter8));
  nand2 gate1760(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1761(.a(s_173), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1762(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1763(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1764(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1163(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1164(.a(gate390inter0), .b(s_88), .O(gate390inter1));
  and2  gate1165(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1166(.a(s_88), .O(gate390inter3));
  inv1  gate1167(.a(s_89), .O(gate390inter4));
  nand2 gate1168(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1169(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1170(.a(G4), .O(gate390inter7));
  inv1  gate1171(.a(G1045), .O(gate390inter8));
  nand2 gate1172(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1173(.a(s_89), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1174(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1175(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1176(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1107(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1108(.a(gate394inter0), .b(s_80), .O(gate394inter1));
  and2  gate1109(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1110(.a(s_80), .O(gate394inter3));
  inv1  gate1111(.a(s_81), .O(gate394inter4));
  nand2 gate1112(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1113(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1114(.a(G8), .O(gate394inter7));
  inv1  gate1115(.a(G1057), .O(gate394inter8));
  nand2 gate1116(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1117(.a(s_81), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1118(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1119(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1120(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2465(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2466(.a(gate396inter0), .b(s_274), .O(gate396inter1));
  and2  gate2467(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2468(.a(s_274), .O(gate396inter3));
  inv1  gate2469(.a(s_275), .O(gate396inter4));
  nand2 gate2470(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2471(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2472(.a(G10), .O(gate396inter7));
  inv1  gate2473(.a(G1063), .O(gate396inter8));
  nand2 gate2474(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2475(.a(s_275), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2476(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2477(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2478(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2451(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2452(.a(gate398inter0), .b(s_272), .O(gate398inter1));
  and2  gate2453(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2454(.a(s_272), .O(gate398inter3));
  inv1  gate2455(.a(s_273), .O(gate398inter4));
  nand2 gate2456(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2457(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2458(.a(G12), .O(gate398inter7));
  inv1  gate2459(.a(G1069), .O(gate398inter8));
  nand2 gate2460(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2461(.a(s_273), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2462(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2463(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2464(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2577(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2578(.a(gate400inter0), .b(s_290), .O(gate400inter1));
  and2  gate2579(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2580(.a(s_290), .O(gate400inter3));
  inv1  gate2581(.a(s_291), .O(gate400inter4));
  nand2 gate2582(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2583(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2584(.a(G14), .O(gate400inter7));
  inv1  gate2585(.a(G1075), .O(gate400inter8));
  nand2 gate2586(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2587(.a(s_291), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2588(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2589(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2590(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2549(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2550(.a(gate401inter0), .b(s_286), .O(gate401inter1));
  and2  gate2551(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2552(.a(s_286), .O(gate401inter3));
  inv1  gate2553(.a(s_287), .O(gate401inter4));
  nand2 gate2554(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2555(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2556(.a(G15), .O(gate401inter7));
  inv1  gate2557(.a(G1078), .O(gate401inter8));
  nand2 gate2558(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2559(.a(s_287), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2560(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2561(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2562(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate729(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate730(.a(gate404inter0), .b(s_26), .O(gate404inter1));
  and2  gate731(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate732(.a(s_26), .O(gate404inter3));
  inv1  gate733(.a(s_27), .O(gate404inter4));
  nand2 gate734(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate735(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate736(.a(G18), .O(gate404inter7));
  inv1  gate737(.a(G1087), .O(gate404inter8));
  nand2 gate738(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate739(.a(s_27), .b(gate404inter3), .O(gate404inter10));
  nor2  gate740(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate741(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate742(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2213(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2214(.a(gate409inter0), .b(s_238), .O(gate409inter1));
  and2  gate2215(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2216(.a(s_238), .O(gate409inter3));
  inv1  gate2217(.a(s_239), .O(gate409inter4));
  nand2 gate2218(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2219(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2220(.a(G23), .O(gate409inter7));
  inv1  gate2221(.a(G1102), .O(gate409inter8));
  nand2 gate2222(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2223(.a(s_239), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2224(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2225(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2226(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2115(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2116(.a(gate410inter0), .b(s_224), .O(gate410inter1));
  and2  gate2117(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2118(.a(s_224), .O(gate410inter3));
  inv1  gate2119(.a(s_225), .O(gate410inter4));
  nand2 gate2120(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2121(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2122(.a(G24), .O(gate410inter7));
  inv1  gate2123(.a(G1105), .O(gate410inter8));
  nand2 gate2124(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2125(.a(s_225), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2126(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2127(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2128(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2129(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2130(.a(gate416inter0), .b(s_226), .O(gate416inter1));
  and2  gate2131(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2132(.a(s_226), .O(gate416inter3));
  inv1  gate2133(.a(s_227), .O(gate416inter4));
  nand2 gate2134(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2135(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2136(.a(G30), .O(gate416inter7));
  inv1  gate2137(.a(G1123), .O(gate416inter8));
  nand2 gate2138(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2139(.a(s_227), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2140(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2141(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2142(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1485(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1486(.a(gate417inter0), .b(s_134), .O(gate417inter1));
  and2  gate1487(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1488(.a(s_134), .O(gate417inter3));
  inv1  gate1489(.a(s_135), .O(gate417inter4));
  nand2 gate1490(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1491(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1492(.a(G31), .O(gate417inter7));
  inv1  gate1493(.a(G1126), .O(gate417inter8));
  nand2 gate1494(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1495(.a(s_135), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1496(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1497(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1498(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1023(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1024(.a(gate418inter0), .b(s_68), .O(gate418inter1));
  and2  gate1025(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1026(.a(s_68), .O(gate418inter3));
  inv1  gate1027(.a(s_69), .O(gate418inter4));
  nand2 gate1028(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1029(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1030(.a(G32), .O(gate418inter7));
  inv1  gate1031(.a(G1129), .O(gate418inter8));
  nand2 gate1032(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1033(.a(s_69), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1034(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1035(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1036(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate827(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate828(.a(gate430inter0), .b(s_40), .O(gate430inter1));
  and2  gate829(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate830(.a(s_40), .O(gate430inter3));
  inv1  gate831(.a(s_41), .O(gate430inter4));
  nand2 gate832(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate833(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate834(.a(G1051), .O(gate430inter7));
  inv1  gate835(.a(G1147), .O(gate430inter8));
  nand2 gate836(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate837(.a(s_41), .b(gate430inter3), .O(gate430inter10));
  nor2  gate838(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate839(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate840(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate631(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate632(.a(gate436inter0), .b(s_12), .O(gate436inter1));
  and2  gate633(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate634(.a(s_12), .O(gate436inter3));
  inv1  gate635(.a(s_13), .O(gate436inter4));
  nand2 gate636(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate637(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate638(.a(G1060), .O(gate436inter7));
  inv1  gate639(.a(G1156), .O(gate436inter8));
  nand2 gate640(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate641(.a(s_13), .b(gate436inter3), .O(gate436inter10));
  nor2  gate642(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate643(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate644(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1233(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1234(.a(gate440inter0), .b(s_98), .O(gate440inter1));
  and2  gate1235(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1236(.a(s_98), .O(gate440inter3));
  inv1  gate1237(.a(s_99), .O(gate440inter4));
  nand2 gate1238(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1239(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1240(.a(G1066), .O(gate440inter7));
  inv1  gate1241(.a(G1162), .O(gate440inter8));
  nand2 gate1242(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1243(.a(s_99), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1244(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1245(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1246(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate869(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate870(.a(gate444inter0), .b(s_46), .O(gate444inter1));
  and2  gate871(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate872(.a(s_46), .O(gate444inter3));
  inv1  gate873(.a(s_47), .O(gate444inter4));
  nand2 gate874(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate875(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate876(.a(G1072), .O(gate444inter7));
  inv1  gate877(.a(G1168), .O(gate444inter8));
  nand2 gate878(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate879(.a(s_47), .b(gate444inter3), .O(gate444inter10));
  nor2  gate880(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate881(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate882(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1919(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1920(.a(gate446inter0), .b(s_196), .O(gate446inter1));
  and2  gate1921(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1922(.a(s_196), .O(gate446inter3));
  inv1  gate1923(.a(s_197), .O(gate446inter4));
  nand2 gate1924(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1925(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1926(.a(G1075), .O(gate446inter7));
  inv1  gate1927(.a(G1171), .O(gate446inter8));
  nand2 gate1928(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1929(.a(s_197), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1930(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1931(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1932(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1135(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1136(.a(gate448inter0), .b(s_84), .O(gate448inter1));
  and2  gate1137(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1138(.a(s_84), .O(gate448inter3));
  inv1  gate1139(.a(s_85), .O(gate448inter4));
  nand2 gate1140(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1141(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1142(.a(G1078), .O(gate448inter7));
  inv1  gate1143(.a(G1174), .O(gate448inter8));
  nand2 gate1144(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1145(.a(s_85), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1146(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1147(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1148(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2045(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2046(.a(gate451inter0), .b(s_214), .O(gate451inter1));
  and2  gate2047(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2048(.a(s_214), .O(gate451inter3));
  inv1  gate2049(.a(s_215), .O(gate451inter4));
  nand2 gate2050(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2051(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2052(.a(G17), .O(gate451inter7));
  inv1  gate2053(.a(G1180), .O(gate451inter8));
  nand2 gate2054(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2055(.a(s_215), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2056(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2057(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2058(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1989(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1990(.a(gate455inter0), .b(s_206), .O(gate455inter1));
  and2  gate1991(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1992(.a(s_206), .O(gate455inter3));
  inv1  gate1993(.a(s_207), .O(gate455inter4));
  nand2 gate1994(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1995(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1996(.a(G19), .O(gate455inter7));
  inv1  gate1997(.a(G1186), .O(gate455inter8));
  nand2 gate1998(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1999(.a(s_207), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2000(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2001(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2002(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1457(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1458(.a(gate456inter0), .b(s_130), .O(gate456inter1));
  and2  gate1459(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1460(.a(s_130), .O(gate456inter3));
  inv1  gate1461(.a(s_131), .O(gate456inter4));
  nand2 gate1462(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1463(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1464(.a(G1090), .O(gate456inter7));
  inv1  gate1465(.a(G1186), .O(gate456inter8));
  nand2 gate1466(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1467(.a(s_131), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1468(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1469(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1470(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1317(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1318(.a(gate457inter0), .b(s_110), .O(gate457inter1));
  and2  gate1319(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1320(.a(s_110), .O(gate457inter3));
  inv1  gate1321(.a(s_111), .O(gate457inter4));
  nand2 gate1322(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1323(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1324(.a(G20), .O(gate457inter7));
  inv1  gate1325(.a(G1189), .O(gate457inter8));
  nand2 gate1326(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1327(.a(s_111), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1328(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1329(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1330(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate939(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate940(.a(gate459inter0), .b(s_56), .O(gate459inter1));
  and2  gate941(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate942(.a(s_56), .O(gate459inter3));
  inv1  gate943(.a(s_57), .O(gate459inter4));
  nand2 gate944(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate945(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate946(.a(G21), .O(gate459inter7));
  inv1  gate947(.a(G1192), .O(gate459inter8));
  nand2 gate948(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate949(.a(s_57), .b(gate459inter3), .O(gate459inter10));
  nor2  gate950(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate951(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate952(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1597(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1598(.a(gate461inter0), .b(s_150), .O(gate461inter1));
  and2  gate1599(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1600(.a(s_150), .O(gate461inter3));
  inv1  gate1601(.a(s_151), .O(gate461inter4));
  nand2 gate1602(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1603(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1604(.a(G22), .O(gate461inter7));
  inv1  gate1605(.a(G1195), .O(gate461inter8));
  nand2 gate1606(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1607(.a(s_151), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1608(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1609(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1610(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2059(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2060(.a(gate462inter0), .b(s_216), .O(gate462inter1));
  and2  gate2061(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2062(.a(s_216), .O(gate462inter3));
  inv1  gate2063(.a(s_217), .O(gate462inter4));
  nand2 gate2064(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2065(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2066(.a(G1099), .O(gate462inter7));
  inv1  gate2067(.a(G1195), .O(gate462inter8));
  nand2 gate2068(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2069(.a(s_217), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2070(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2071(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2072(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1625(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1626(.a(gate464inter0), .b(s_154), .O(gate464inter1));
  and2  gate1627(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1628(.a(s_154), .O(gate464inter3));
  inv1  gate1629(.a(s_155), .O(gate464inter4));
  nand2 gate1630(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1631(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1632(.a(G1102), .O(gate464inter7));
  inv1  gate1633(.a(G1198), .O(gate464inter8));
  nand2 gate1634(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1635(.a(s_155), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1636(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1637(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1638(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2409(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2410(.a(gate469inter0), .b(s_266), .O(gate469inter1));
  and2  gate2411(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2412(.a(s_266), .O(gate469inter3));
  inv1  gate2413(.a(s_267), .O(gate469inter4));
  nand2 gate2414(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2415(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2416(.a(G26), .O(gate469inter7));
  inv1  gate2417(.a(G1207), .O(gate469inter8));
  nand2 gate2418(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2419(.a(s_267), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2420(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2421(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2422(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1891(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1892(.a(gate471inter0), .b(s_192), .O(gate471inter1));
  and2  gate1893(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1894(.a(s_192), .O(gate471inter3));
  inv1  gate1895(.a(s_193), .O(gate471inter4));
  nand2 gate1896(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1897(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1898(.a(G27), .O(gate471inter7));
  inv1  gate1899(.a(G1210), .O(gate471inter8));
  nand2 gate1900(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1901(.a(s_193), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1902(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1903(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1904(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1667(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1668(.a(gate473inter0), .b(s_160), .O(gate473inter1));
  and2  gate1669(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1670(.a(s_160), .O(gate473inter3));
  inv1  gate1671(.a(s_161), .O(gate473inter4));
  nand2 gate1672(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1673(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1674(.a(G28), .O(gate473inter7));
  inv1  gate1675(.a(G1213), .O(gate473inter8));
  nand2 gate1676(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1677(.a(s_161), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1678(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1679(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1680(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate813(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate814(.a(gate475inter0), .b(s_38), .O(gate475inter1));
  and2  gate815(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate816(.a(s_38), .O(gate475inter3));
  inv1  gate817(.a(s_39), .O(gate475inter4));
  nand2 gate818(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate819(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate820(.a(G29), .O(gate475inter7));
  inv1  gate821(.a(G1216), .O(gate475inter8));
  nand2 gate822(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate823(.a(s_39), .b(gate475inter3), .O(gate475inter10));
  nor2  gate824(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate825(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate826(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2227(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2228(.a(gate476inter0), .b(s_240), .O(gate476inter1));
  and2  gate2229(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2230(.a(s_240), .O(gate476inter3));
  inv1  gate2231(.a(s_241), .O(gate476inter4));
  nand2 gate2232(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2233(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2234(.a(G1120), .O(gate476inter7));
  inv1  gate2235(.a(G1216), .O(gate476inter8));
  nand2 gate2236(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2237(.a(s_241), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2238(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2239(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2240(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1401(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1402(.a(gate480inter0), .b(s_122), .O(gate480inter1));
  and2  gate1403(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1404(.a(s_122), .O(gate480inter3));
  inv1  gate1405(.a(s_123), .O(gate480inter4));
  nand2 gate1406(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1407(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1408(.a(G1126), .O(gate480inter7));
  inv1  gate1409(.a(G1222), .O(gate480inter8));
  nand2 gate1410(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1411(.a(s_123), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1412(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1413(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1414(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1289(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1290(.a(gate484inter0), .b(s_106), .O(gate484inter1));
  and2  gate1291(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1292(.a(s_106), .O(gate484inter3));
  inv1  gate1293(.a(s_107), .O(gate484inter4));
  nand2 gate1294(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1295(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1296(.a(G1230), .O(gate484inter7));
  inv1  gate1297(.a(G1231), .O(gate484inter8));
  nand2 gate1298(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1299(.a(s_107), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1300(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1301(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1302(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1723(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1724(.a(gate486inter0), .b(s_168), .O(gate486inter1));
  and2  gate1725(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1726(.a(s_168), .O(gate486inter3));
  inv1  gate1727(.a(s_169), .O(gate486inter4));
  nand2 gate1728(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1729(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1730(.a(G1234), .O(gate486inter7));
  inv1  gate1731(.a(G1235), .O(gate486inter8));
  nand2 gate1732(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1733(.a(s_169), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1734(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1735(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1736(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2339(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2340(.a(gate487inter0), .b(s_256), .O(gate487inter1));
  and2  gate2341(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2342(.a(s_256), .O(gate487inter3));
  inv1  gate2343(.a(s_257), .O(gate487inter4));
  nand2 gate2344(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2345(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2346(.a(G1236), .O(gate487inter7));
  inv1  gate2347(.a(G1237), .O(gate487inter8));
  nand2 gate2348(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2349(.a(s_257), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2350(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2351(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2352(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1639(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1640(.a(gate489inter0), .b(s_156), .O(gate489inter1));
  and2  gate1641(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1642(.a(s_156), .O(gate489inter3));
  inv1  gate1643(.a(s_157), .O(gate489inter4));
  nand2 gate1644(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1645(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1646(.a(G1240), .O(gate489inter7));
  inv1  gate1647(.a(G1241), .O(gate489inter8));
  nand2 gate1648(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1649(.a(s_157), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1650(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1651(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1652(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2157(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2158(.a(gate493inter0), .b(s_230), .O(gate493inter1));
  and2  gate2159(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2160(.a(s_230), .O(gate493inter3));
  inv1  gate2161(.a(s_231), .O(gate493inter4));
  nand2 gate2162(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2163(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2164(.a(G1248), .O(gate493inter7));
  inv1  gate2165(.a(G1249), .O(gate493inter8));
  nand2 gate2166(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2167(.a(s_231), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2168(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2169(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2170(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate617(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate618(.a(gate494inter0), .b(s_10), .O(gate494inter1));
  and2  gate619(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate620(.a(s_10), .O(gate494inter3));
  inv1  gate621(.a(s_11), .O(gate494inter4));
  nand2 gate622(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate623(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate624(.a(G1250), .O(gate494inter7));
  inv1  gate625(.a(G1251), .O(gate494inter8));
  nand2 gate626(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate627(.a(s_11), .b(gate494inter3), .O(gate494inter10));
  nor2  gate628(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate629(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate630(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate967(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate968(.a(gate498inter0), .b(s_60), .O(gate498inter1));
  and2  gate969(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate970(.a(s_60), .O(gate498inter3));
  inv1  gate971(.a(s_61), .O(gate498inter4));
  nand2 gate972(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate973(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate974(.a(G1258), .O(gate498inter7));
  inv1  gate975(.a(G1259), .O(gate498inter8));
  nand2 gate976(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate977(.a(s_61), .b(gate498inter3), .O(gate498inter10));
  nor2  gate978(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate979(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate980(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate757(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate758(.a(gate500inter0), .b(s_30), .O(gate500inter1));
  and2  gate759(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate760(.a(s_30), .O(gate500inter3));
  inv1  gate761(.a(s_31), .O(gate500inter4));
  nand2 gate762(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate763(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate764(.a(G1262), .O(gate500inter7));
  inv1  gate765(.a(G1263), .O(gate500inter8));
  nand2 gate766(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate767(.a(s_31), .b(gate500inter3), .O(gate500inter10));
  nor2  gate768(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate769(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate770(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1779(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1780(.a(gate504inter0), .b(s_176), .O(gate504inter1));
  and2  gate1781(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1782(.a(s_176), .O(gate504inter3));
  inv1  gate1783(.a(s_177), .O(gate504inter4));
  nand2 gate1784(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1785(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1786(.a(G1270), .O(gate504inter7));
  inv1  gate1787(.a(G1271), .O(gate504inter8));
  nand2 gate1788(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1789(.a(s_177), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1790(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1791(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1792(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1065(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1066(.a(gate505inter0), .b(s_74), .O(gate505inter1));
  and2  gate1067(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1068(.a(s_74), .O(gate505inter3));
  inv1  gate1069(.a(s_75), .O(gate505inter4));
  nand2 gate1070(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1071(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1072(.a(G1272), .O(gate505inter7));
  inv1  gate1073(.a(G1273), .O(gate505inter8));
  nand2 gate1074(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1075(.a(s_75), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1076(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1077(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1078(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1681(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1682(.a(gate506inter0), .b(s_162), .O(gate506inter1));
  and2  gate1683(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1684(.a(s_162), .O(gate506inter3));
  inv1  gate1685(.a(s_163), .O(gate506inter4));
  nand2 gate1686(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1687(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1688(.a(G1274), .O(gate506inter7));
  inv1  gate1689(.a(G1275), .O(gate506inter8));
  nand2 gate1690(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1691(.a(s_163), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1692(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1693(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1694(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate2101(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2102(.a(gate507inter0), .b(s_222), .O(gate507inter1));
  and2  gate2103(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2104(.a(s_222), .O(gate507inter3));
  inv1  gate2105(.a(s_223), .O(gate507inter4));
  nand2 gate2106(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2107(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2108(.a(G1276), .O(gate507inter7));
  inv1  gate2109(.a(G1277), .O(gate507inter8));
  nand2 gate2110(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2111(.a(s_223), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2112(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2113(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2114(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1359(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1360(.a(gate511inter0), .b(s_116), .O(gate511inter1));
  and2  gate1361(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1362(.a(s_116), .O(gate511inter3));
  inv1  gate1363(.a(s_117), .O(gate511inter4));
  nand2 gate1364(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1365(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1366(.a(G1284), .O(gate511inter7));
  inv1  gate1367(.a(G1285), .O(gate511inter8));
  nand2 gate1368(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1369(.a(s_117), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1370(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1371(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1372(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate2311(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2312(.a(gate512inter0), .b(s_252), .O(gate512inter1));
  and2  gate2313(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2314(.a(s_252), .O(gate512inter3));
  inv1  gate2315(.a(s_253), .O(gate512inter4));
  nand2 gate2316(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2317(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2318(.a(G1286), .O(gate512inter7));
  inv1  gate2319(.a(G1287), .O(gate512inter8));
  nand2 gate2320(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2321(.a(s_253), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2322(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2323(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2324(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule