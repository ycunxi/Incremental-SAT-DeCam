module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1471(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1472(.a(gate12inter0), .b(s_132), .O(gate12inter1));
  and2  gate1473(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1474(.a(s_132), .O(gate12inter3));
  inv1  gate1475(.a(s_133), .O(gate12inter4));
  nand2 gate1476(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1477(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1478(.a(G7), .O(gate12inter7));
  inv1  gate1479(.a(G8), .O(gate12inter8));
  nand2 gate1480(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1481(.a(s_133), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1482(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1483(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1484(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1135(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1136(.a(gate14inter0), .b(s_84), .O(gate14inter1));
  and2  gate1137(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1138(.a(s_84), .O(gate14inter3));
  inv1  gate1139(.a(s_85), .O(gate14inter4));
  nand2 gate1140(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1141(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1142(.a(G11), .O(gate14inter7));
  inv1  gate1143(.a(G12), .O(gate14inter8));
  nand2 gate1144(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1145(.a(s_85), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1146(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1147(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1148(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2073(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2074(.a(gate17inter0), .b(s_218), .O(gate17inter1));
  and2  gate2075(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2076(.a(s_218), .O(gate17inter3));
  inv1  gate2077(.a(s_219), .O(gate17inter4));
  nand2 gate2078(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2079(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2080(.a(G17), .O(gate17inter7));
  inv1  gate2081(.a(G18), .O(gate17inter8));
  nand2 gate2082(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2083(.a(s_219), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2084(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2085(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2086(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1527(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1528(.a(gate22inter0), .b(s_140), .O(gate22inter1));
  and2  gate1529(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1530(.a(s_140), .O(gate22inter3));
  inv1  gate1531(.a(s_141), .O(gate22inter4));
  nand2 gate1532(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1533(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1534(.a(G27), .O(gate22inter7));
  inv1  gate1535(.a(G28), .O(gate22inter8));
  nand2 gate1536(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1537(.a(s_141), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1538(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1539(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1540(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1275(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1276(.a(gate24inter0), .b(s_104), .O(gate24inter1));
  and2  gate1277(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1278(.a(s_104), .O(gate24inter3));
  inv1  gate1279(.a(s_105), .O(gate24inter4));
  nand2 gate1280(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1281(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1282(.a(G31), .O(gate24inter7));
  inv1  gate1283(.a(G32), .O(gate24inter8));
  nand2 gate1284(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1285(.a(s_105), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1286(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1287(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1288(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1653(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1654(.a(gate26inter0), .b(s_158), .O(gate26inter1));
  and2  gate1655(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1656(.a(s_158), .O(gate26inter3));
  inv1  gate1657(.a(s_159), .O(gate26inter4));
  nand2 gate1658(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1659(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1660(.a(G9), .O(gate26inter7));
  inv1  gate1661(.a(G13), .O(gate26inter8));
  nand2 gate1662(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1663(.a(s_159), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1664(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1665(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1666(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate645(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate646(.a(gate27inter0), .b(s_14), .O(gate27inter1));
  and2  gate647(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate648(.a(s_14), .O(gate27inter3));
  inv1  gate649(.a(s_15), .O(gate27inter4));
  nand2 gate650(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate651(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate652(.a(G2), .O(gate27inter7));
  inv1  gate653(.a(G6), .O(gate27inter8));
  nand2 gate654(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate655(.a(s_15), .b(gate27inter3), .O(gate27inter10));
  nor2  gate656(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate657(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate658(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1163(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1164(.a(gate30inter0), .b(s_88), .O(gate30inter1));
  and2  gate1165(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1166(.a(s_88), .O(gate30inter3));
  inv1  gate1167(.a(s_89), .O(gate30inter4));
  nand2 gate1168(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1169(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1170(.a(G11), .O(gate30inter7));
  inv1  gate1171(.a(G15), .O(gate30inter8));
  nand2 gate1172(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1173(.a(s_89), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1174(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1175(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1176(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1373(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1374(.a(gate38inter0), .b(s_118), .O(gate38inter1));
  and2  gate1375(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1376(.a(s_118), .O(gate38inter3));
  inv1  gate1377(.a(s_119), .O(gate38inter4));
  nand2 gate1378(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1379(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1380(.a(G27), .O(gate38inter7));
  inv1  gate1381(.a(G31), .O(gate38inter8));
  nand2 gate1382(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1383(.a(s_119), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1384(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1385(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1386(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate617(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate618(.a(gate43inter0), .b(s_10), .O(gate43inter1));
  and2  gate619(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate620(.a(s_10), .O(gate43inter3));
  inv1  gate621(.a(s_11), .O(gate43inter4));
  nand2 gate622(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate623(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate624(.a(G3), .O(gate43inter7));
  inv1  gate625(.a(G269), .O(gate43inter8));
  nand2 gate626(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate627(.a(s_11), .b(gate43inter3), .O(gate43inter10));
  nor2  gate628(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate629(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate630(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1611(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1612(.a(gate51inter0), .b(s_152), .O(gate51inter1));
  and2  gate1613(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1614(.a(s_152), .O(gate51inter3));
  inv1  gate1615(.a(s_153), .O(gate51inter4));
  nand2 gate1616(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1617(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1618(.a(G11), .O(gate51inter7));
  inv1  gate1619(.a(G281), .O(gate51inter8));
  nand2 gate1620(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1621(.a(s_153), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1622(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1623(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1624(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate2129(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2130(.a(gate52inter0), .b(s_226), .O(gate52inter1));
  and2  gate2131(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2132(.a(s_226), .O(gate52inter3));
  inv1  gate2133(.a(s_227), .O(gate52inter4));
  nand2 gate2134(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2135(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2136(.a(G12), .O(gate52inter7));
  inv1  gate2137(.a(G281), .O(gate52inter8));
  nand2 gate2138(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2139(.a(s_227), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2140(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2141(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2142(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2115(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2116(.a(gate54inter0), .b(s_224), .O(gate54inter1));
  and2  gate2117(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2118(.a(s_224), .O(gate54inter3));
  inv1  gate2119(.a(s_225), .O(gate54inter4));
  nand2 gate2120(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2121(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2122(.a(G14), .O(gate54inter7));
  inv1  gate2123(.a(G284), .O(gate54inter8));
  nand2 gate2124(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2125(.a(s_225), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2126(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2127(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2128(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate953(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate954(.a(gate56inter0), .b(s_58), .O(gate56inter1));
  and2  gate955(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate956(.a(s_58), .O(gate56inter3));
  inv1  gate957(.a(s_59), .O(gate56inter4));
  nand2 gate958(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate959(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate960(.a(G16), .O(gate56inter7));
  inv1  gate961(.a(G287), .O(gate56inter8));
  nand2 gate962(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate963(.a(s_59), .b(gate56inter3), .O(gate56inter10));
  nor2  gate964(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate965(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate966(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1079(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1080(.a(gate62inter0), .b(s_76), .O(gate62inter1));
  and2  gate1081(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1082(.a(s_76), .O(gate62inter3));
  inv1  gate1083(.a(s_77), .O(gate62inter4));
  nand2 gate1084(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1085(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1086(.a(G22), .O(gate62inter7));
  inv1  gate1087(.a(G296), .O(gate62inter8));
  nand2 gate1088(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1089(.a(s_77), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1090(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1091(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1092(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate981(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate982(.a(gate65inter0), .b(s_62), .O(gate65inter1));
  and2  gate983(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate984(.a(s_62), .O(gate65inter3));
  inv1  gate985(.a(s_63), .O(gate65inter4));
  nand2 gate986(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate987(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate988(.a(G25), .O(gate65inter7));
  inv1  gate989(.a(G302), .O(gate65inter8));
  nand2 gate990(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate991(.a(s_63), .b(gate65inter3), .O(gate65inter10));
  nor2  gate992(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate993(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate994(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1429(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1430(.a(gate66inter0), .b(s_126), .O(gate66inter1));
  and2  gate1431(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1432(.a(s_126), .O(gate66inter3));
  inv1  gate1433(.a(s_127), .O(gate66inter4));
  nand2 gate1434(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1435(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1436(.a(G26), .O(gate66inter7));
  inv1  gate1437(.a(G302), .O(gate66inter8));
  nand2 gate1438(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1439(.a(s_127), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1440(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1441(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1442(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1177(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1178(.a(gate72inter0), .b(s_90), .O(gate72inter1));
  and2  gate1179(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1180(.a(s_90), .O(gate72inter3));
  inv1  gate1181(.a(s_91), .O(gate72inter4));
  nand2 gate1182(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1183(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1184(.a(G32), .O(gate72inter7));
  inv1  gate1185(.a(G311), .O(gate72inter8));
  nand2 gate1186(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1187(.a(s_91), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1188(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1189(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1190(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate827(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate828(.a(gate75inter0), .b(s_40), .O(gate75inter1));
  and2  gate829(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate830(.a(s_40), .O(gate75inter3));
  inv1  gate831(.a(s_41), .O(gate75inter4));
  nand2 gate832(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate833(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate834(.a(G9), .O(gate75inter7));
  inv1  gate835(.a(G317), .O(gate75inter8));
  nand2 gate836(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate837(.a(s_41), .b(gate75inter3), .O(gate75inter10));
  nor2  gate838(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate839(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate840(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1359(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1360(.a(gate76inter0), .b(s_116), .O(gate76inter1));
  and2  gate1361(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1362(.a(s_116), .O(gate76inter3));
  inv1  gate1363(.a(s_117), .O(gate76inter4));
  nand2 gate1364(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1365(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1366(.a(G13), .O(gate76inter7));
  inv1  gate1367(.a(G317), .O(gate76inter8));
  nand2 gate1368(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1369(.a(s_117), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1370(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1371(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1372(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate2213(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2214(.a(gate77inter0), .b(s_238), .O(gate77inter1));
  and2  gate2215(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2216(.a(s_238), .O(gate77inter3));
  inv1  gate2217(.a(s_239), .O(gate77inter4));
  nand2 gate2218(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2219(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2220(.a(G2), .O(gate77inter7));
  inv1  gate2221(.a(G320), .O(gate77inter8));
  nand2 gate2222(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2223(.a(s_239), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2224(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2225(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2226(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1639(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1640(.a(gate78inter0), .b(s_156), .O(gate78inter1));
  and2  gate1641(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1642(.a(s_156), .O(gate78inter3));
  inv1  gate1643(.a(s_157), .O(gate78inter4));
  nand2 gate1644(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1645(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1646(.a(G6), .O(gate78inter7));
  inv1  gate1647(.a(G320), .O(gate78inter8));
  nand2 gate1648(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1649(.a(s_157), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1650(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1651(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1652(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1569(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1570(.a(gate82inter0), .b(s_146), .O(gate82inter1));
  and2  gate1571(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1572(.a(s_146), .O(gate82inter3));
  inv1  gate1573(.a(s_147), .O(gate82inter4));
  nand2 gate1574(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1575(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1576(.a(G7), .O(gate82inter7));
  inv1  gate1577(.a(G326), .O(gate82inter8));
  nand2 gate1578(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1579(.a(s_147), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1580(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1581(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1582(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1387(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1388(.a(gate83inter0), .b(s_120), .O(gate83inter1));
  and2  gate1389(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1390(.a(s_120), .O(gate83inter3));
  inv1  gate1391(.a(s_121), .O(gate83inter4));
  nand2 gate1392(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1393(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1394(.a(G11), .O(gate83inter7));
  inv1  gate1395(.a(G329), .O(gate83inter8));
  nand2 gate1396(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1397(.a(s_121), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1398(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1399(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1400(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1009(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1010(.a(gate86inter0), .b(s_66), .O(gate86inter1));
  and2  gate1011(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1012(.a(s_66), .O(gate86inter3));
  inv1  gate1013(.a(s_67), .O(gate86inter4));
  nand2 gate1014(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1015(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1016(.a(G8), .O(gate86inter7));
  inv1  gate1017(.a(G332), .O(gate86inter8));
  nand2 gate1018(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1019(.a(s_67), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1020(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1021(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1022(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2185(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2186(.a(gate91inter0), .b(s_234), .O(gate91inter1));
  and2  gate2187(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2188(.a(s_234), .O(gate91inter3));
  inv1  gate2189(.a(s_235), .O(gate91inter4));
  nand2 gate2190(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2191(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2192(.a(G25), .O(gate91inter7));
  inv1  gate2193(.a(G341), .O(gate91inter8));
  nand2 gate2194(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2195(.a(s_235), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2196(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2197(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2198(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1121(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1122(.a(gate94inter0), .b(s_82), .O(gate94inter1));
  and2  gate1123(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1124(.a(s_82), .O(gate94inter3));
  inv1  gate1125(.a(s_83), .O(gate94inter4));
  nand2 gate1126(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1127(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1128(.a(G22), .O(gate94inter7));
  inv1  gate1129(.a(G344), .O(gate94inter8));
  nand2 gate1130(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1131(.a(s_83), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1132(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1133(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1134(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1205(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1206(.a(gate95inter0), .b(s_94), .O(gate95inter1));
  and2  gate1207(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1208(.a(s_94), .O(gate95inter3));
  inv1  gate1209(.a(s_95), .O(gate95inter4));
  nand2 gate1210(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1211(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1212(.a(G26), .O(gate95inter7));
  inv1  gate1213(.a(G347), .O(gate95inter8));
  nand2 gate1214(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1215(.a(s_95), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1216(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1217(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1218(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate701(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate702(.a(gate99inter0), .b(s_22), .O(gate99inter1));
  and2  gate703(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate704(.a(s_22), .O(gate99inter3));
  inv1  gate705(.a(s_23), .O(gate99inter4));
  nand2 gate706(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate707(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate708(.a(G27), .O(gate99inter7));
  inv1  gate709(.a(G353), .O(gate99inter8));
  nand2 gate710(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate711(.a(s_23), .b(gate99inter3), .O(gate99inter10));
  nor2  gate712(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate713(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate714(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2171(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2172(.a(gate102inter0), .b(s_232), .O(gate102inter1));
  and2  gate2173(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2174(.a(s_232), .O(gate102inter3));
  inv1  gate2175(.a(s_233), .O(gate102inter4));
  nand2 gate2176(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2177(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2178(.a(G24), .O(gate102inter7));
  inv1  gate2179(.a(G356), .O(gate102inter8));
  nand2 gate2180(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2181(.a(s_233), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2182(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2183(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2184(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1835(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1836(.a(gate107inter0), .b(s_184), .O(gate107inter1));
  and2  gate1837(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1838(.a(s_184), .O(gate107inter3));
  inv1  gate1839(.a(s_185), .O(gate107inter4));
  nand2 gate1840(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1841(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1842(.a(G366), .O(gate107inter7));
  inv1  gate1843(.a(G367), .O(gate107inter8));
  nand2 gate1844(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1845(.a(s_185), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1846(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1847(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1848(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1289(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1290(.a(gate109inter0), .b(s_106), .O(gate109inter1));
  and2  gate1291(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1292(.a(s_106), .O(gate109inter3));
  inv1  gate1293(.a(s_107), .O(gate109inter4));
  nand2 gate1294(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1295(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1296(.a(G370), .O(gate109inter7));
  inv1  gate1297(.a(G371), .O(gate109inter8));
  nand2 gate1298(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1299(.a(s_107), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1300(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1301(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1302(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1723(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1724(.a(gate110inter0), .b(s_168), .O(gate110inter1));
  and2  gate1725(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1726(.a(s_168), .O(gate110inter3));
  inv1  gate1727(.a(s_169), .O(gate110inter4));
  nand2 gate1728(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1729(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1730(.a(G372), .O(gate110inter7));
  inv1  gate1731(.a(G373), .O(gate110inter8));
  nand2 gate1732(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1733(.a(s_169), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1734(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1735(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1736(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1331(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1332(.a(gate115inter0), .b(s_112), .O(gate115inter1));
  and2  gate1333(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1334(.a(s_112), .O(gate115inter3));
  inv1  gate1335(.a(s_113), .O(gate115inter4));
  nand2 gate1336(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1337(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1338(.a(G382), .O(gate115inter7));
  inv1  gate1339(.a(G383), .O(gate115inter8));
  nand2 gate1340(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1341(.a(s_113), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1342(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1343(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1344(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1051(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1052(.a(gate121inter0), .b(s_72), .O(gate121inter1));
  and2  gate1053(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1054(.a(s_72), .O(gate121inter3));
  inv1  gate1055(.a(s_73), .O(gate121inter4));
  nand2 gate1056(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1057(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1058(.a(G394), .O(gate121inter7));
  inv1  gate1059(.a(G395), .O(gate121inter8));
  nand2 gate1060(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1061(.a(s_73), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1062(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1063(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1064(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1233(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1234(.a(gate122inter0), .b(s_98), .O(gate122inter1));
  and2  gate1235(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1236(.a(s_98), .O(gate122inter3));
  inv1  gate1237(.a(s_99), .O(gate122inter4));
  nand2 gate1238(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1239(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1240(.a(G396), .O(gate122inter7));
  inv1  gate1241(.a(G397), .O(gate122inter8));
  nand2 gate1242(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1243(.a(s_99), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1244(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1245(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1246(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1345(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1346(.a(gate123inter0), .b(s_114), .O(gate123inter1));
  and2  gate1347(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1348(.a(s_114), .O(gate123inter3));
  inv1  gate1349(.a(s_115), .O(gate123inter4));
  nand2 gate1350(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1351(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1352(.a(G398), .O(gate123inter7));
  inv1  gate1353(.a(G399), .O(gate123inter8));
  nand2 gate1354(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1355(.a(s_115), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1356(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1357(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1358(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate547(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate548(.a(gate126inter0), .b(s_0), .O(gate126inter1));
  and2  gate549(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate550(.a(s_0), .O(gate126inter3));
  inv1  gate551(.a(s_1), .O(gate126inter4));
  nand2 gate552(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate553(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate554(.a(G404), .O(gate126inter7));
  inv1  gate555(.a(G405), .O(gate126inter8));
  nand2 gate556(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate557(.a(s_1), .b(gate126inter3), .O(gate126inter10));
  nor2  gate558(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate559(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate560(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1597(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1598(.a(gate127inter0), .b(s_150), .O(gate127inter1));
  and2  gate1599(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1600(.a(s_150), .O(gate127inter3));
  inv1  gate1601(.a(s_151), .O(gate127inter4));
  nand2 gate1602(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1603(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1604(.a(G406), .O(gate127inter7));
  inv1  gate1605(.a(G407), .O(gate127inter8));
  nand2 gate1606(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1607(.a(s_151), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1608(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1609(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1610(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate813(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate814(.a(gate128inter0), .b(s_38), .O(gate128inter1));
  and2  gate815(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate816(.a(s_38), .O(gate128inter3));
  inv1  gate817(.a(s_39), .O(gate128inter4));
  nand2 gate818(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate819(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate820(.a(G408), .O(gate128inter7));
  inv1  gate821(.a(G409), .O(gate128inter8));
  nand2 gate822(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate823(.a(s_39), .b(gate128inter3), .O(gate128inter10));
  nor2  gate824(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate825(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate826(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate659(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate660(.a(gate130inter0), .b(s_16), .O(gate130inter1));
  and2  gate661(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate662(.a(s_16), .O(gate130inter3));
  inv1  gate663(.a(s_17), .O(gate130inter4));
  nand2 gate664(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate665(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate666(.a(G412), .O(gate130inter7));
  inv1  gate667(.a(G413), .O(gate130inter8));
  nand2 gate668(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate669(.a(s_17), .b(gate130inter3), .O(gate130inter10));
  nor2  gate670(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate671(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate672(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1709(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1710(.a(gate133inter0), .b(s_166), .O(gate133inter1));
  and2  gate1711(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1712(.a(s_166), .O(gate133inter3));
  inv1  gate1713(.a(s_167), .O(gate133inter4));
  nand2 gate1714(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1715(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1716(.a(G418), .O(gate133inter7));
  inv1  gate1717(.a(G419), .O(gate133inter8));
  nand2 gate1718(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1719(.a(s_167), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1720(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1721(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1722(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1513(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1514(.a(gate138inter0), .b(s_138), .O(gate138inter1));
  and2  gate1515(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1516(.a(s_138), .O(gate138inter3));
  inv1  gate1517(.a(s_139), .O(gate138inter4));
  nand2 gate1518(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1519(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1520(.a(G432), .O(gate138inter7));
  inv1  gate1521(.a(G435), .O(gate138inter8));
  nand2 gate1522(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1523(.a(s_139), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1524(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1525(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1526(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate855(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate856(.a(gate144inter0), .b(s_44), .O(gate144inter1));
  and2  gate857(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate858(.a(s_44), .O(gate144inter3));
  inv1  gate859(.a(s_45), .O(gate144inter4));
  nand2 gate860(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate861(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate862(.a(G468), .O(gate144inter7));
  inv1  gate863(.a(G471), .O(gate144inter8));
  nand2 gate864(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate865(.a(s_45), .b(gate144inter3), .O(gate144inter10));
  nor2  gate866(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate867(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate868(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1625(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1626(.a(gate146inter0), .b(s_154), .O(gate146inter1));
  and2  gate1627(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1628(.a(s_154), .O(gate146inter3));
  inv1  gate1629(.a(s_155), .O(gate146inter4));
  nand2 gate1630(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1631(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1632(.a(G480), .O(gate146inter7));
  inv1  gate1633(.a(G483), .O(gate146inter8));
  nand2 gate1634(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1635(.a(s_155), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1636(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1637(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1638(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2017(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2018(.a(gate147inter0), .b(s_210), .O(gate147inter1));
  and2  gate2019(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2020(.a(s_210), .O(gate147inter3));
  inv1  gate2021(.a(s_211), .O(gate147inter4));
  nand2 gate2022(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2023(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2024(.a(G486), .O(gate147inter7));
  inv1  gate2025(.a(G489), .O(gate147inter8));
  nand2 gate2026(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2027(.a(s_211), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2028(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2029(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2030(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2199(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2200(.a(gate149inter0), .b(s_236), .O(gate149inter1));
  and2  gate2201(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2202(.a(s_236), .O(gate149inter3));
  inv1  gate2203(.a(s_237), .O(gate149inter4));
  nand2 gate2204(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2205(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2206(.a(G498), .O(gate149inter7));
  inv1  gate2207(.a(G501), .O(gate149inter8));
  nand2 gate2208(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2209(.a(s_237), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2210(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2211(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2212(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1905(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1906(.a(gate154inter0), .b(s_194), .O(gate154inter1));
  and2  gate1907(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1908(.a(s_194), .O(gate154inter3));
  inv1  gate1909(.a(s_195), .O(gate154inter4));
  nand2 gate1910(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1911(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1912(.a(G429), .O(gate154inter7));
  inv1  gate1913(.a(G522), .O(gate154inter8));
  nand2 gate1914(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1915(.a(s_195), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1916(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1917(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1918(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1499(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1500(.a(gate155inter0), .b(s_136), .O(gate155inter1));
  and2  gate1501(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1502(.a(s_136), .O(gate155inter3));
  inv1  gate1503(.a(s_137), .O(gate155inter4));
  nand2 gate1504(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1505(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1506(.a(G432), .O(gate155inter7));
  inv1  gate1507(.a(G525), .O(gate155inter8));
  nand2 gate1508(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1509(.a(s_137), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1510(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1511(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1512(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2045(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2046(.a(gate157inter0), .b(s_214), .O(gate157inter1));
  and2  gate2047(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2048(.a(s_214), .O(gate157inter3));
  inv1  gate2049(.a(s_215), .O(gate157inter4));
  nand2 gate2050(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2051(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2052(.a(G438), .O(gate157inter7));
  inv1  gate2053(.a(G528), .O(gate157inter8));
  nand2 gate2054(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2055(.a(s_215), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2056(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2057(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2058(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate883(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate884(.a(gate161inter0), .b(s_48), .O(gate161inter1));
  and2  gate885(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate886(.a(s_48), .O(gate161inter3));
  inv1  gate887(.a(s_49), .O(gate161inter4));
  nand2 gate888(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate889(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate890(.a(G450), .O(gate161inter7));
  inv1  gate891(.a(G534), .O(gate161inter8));
  nand2 gate892(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate893(.a(s_49), .b(gate161inter3), .O(gate161inter10));
  nor2  gate894(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate895(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate896(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1779(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1780(.a(gate175inter0), .b(s_176), .O(gate175inter1));
  and2  gate1781(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1782(.a(s_176), .O(gate175inter3));
  inv1  gate1783(.a(s_177), .O(gate175inter4));
  nand2 gate1784(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1785(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1786(.a(G492), .O(gate175inter7));
  inv1  gate1787(.a(G555), .O(gate175inter8));
  nand2 gate1788(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1789(.a(s_177), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1790(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1791(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1792(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate939(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate940(.a(gate184inter0), .b(s_56), .O(gate184inter1));
  and2  gate941(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate942(.a(s_56), .O(gate184inter3));
  inv1  gate943(.a(s_57), .O(gate184inter4));
  nand2 gate944(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate945(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate946(.a(G519), .O(gate184inter7));
  inv1  gate947(.a(G567), .O(gate184inter8));
  nand2 gate948(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate949(.a(s_57), .b(gate184inter3), .O(gate184inter10));
  nor2  gate950(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate951(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate952(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1737(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1738(.a(gate185inter0), .b(s_170), .O(gate185inter1));
  and2  gate1739(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1740(.a(s_170), .O(gate185inter3));
  inv1  gate1741(.a(s_171), .O(gate185inter4));
  nand2 gate1742(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1743(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1744(.a(G570), .O(gate185inter7));
  inv1  gate1745(.a(G571), .O(gate185inter8));
  nand2 gate1746(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1747(.a(s_171), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1748(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1749(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1750(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate771(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate772(.a(gate188inter0), .b(s_32), .O(gate188inter1));
  and2  gate773(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate774(.a(s_32), .O(gate188inter3));
  inv1  gate775(.a(s_33), .O(gate188inter4));
  nand2 gate776(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate777(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate778(.a(G576), .O(gate188inter7));
  inv1  gate779(.a(G577), .O(gate188inter8));
  nand2 gate780(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate781(.a(s_33), .b(gate188inter3), .O(gate188inter10));
  nor2  gate782(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate783(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate784(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate673(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate674(.a(gate190inter0), .b(s_18), .O(gate190inter1));
  and2  gate675(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate676(.a(s_18), .O(gate190inter3));
  inv1  gate677(.a(s_19), .O(gate190inter4));
  nand2 gate678(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate679(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate680(.a(G580), .O(gate190inter7));
  inv1  gate681(.a(G581), .O(gate190inter8));
  nand2 gate682(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate683(.a(s_19), .b(gate190inter3), .O(gate190inter10));
  nor2  gate684(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate685(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate686(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1947(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1948(.a(gate193inter0), .b(s_200), .O(gate193inter1));
  and2  gate1949(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1950(.a(s_200), .O(gate193inter3));
  inv1  gate1951(.a(s_201), .O(gate193inter4));
  nand2 gate1952(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1953(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1954(.a(G586), .O(gate193inter7));
  inv1  gate1955(.a(G587), .O(gate193inter8));
  nand2 gate1956(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1957(.a(s_201), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1958(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1959(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1960(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2003(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2004(.a(gate201inter0), .b(s_208), .O(gate201inter1));
  and2  gate2005(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2006(.a(s_208), .O(gate201inter3));
  inv1  gate2007(.a(s_209), .O(gate201inter4));
  nand2 gate2008(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2009(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2010(.a(G602), .O(gate201inter7));
  inv1  gate2011(.a(G607), .O(gate201inter8));
  nand2 gate2012(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2013(.a(s_209), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2014(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2015(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2016(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate2059(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2060(.a(gate202inter0), .b(s_216), .O(gate202inter1));
  and2  gate2061(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2062(.a(s_216), .O(gate202inter3));
  inv1  gate2063(.a(s_217), .O(gate202inter4));
  nand2 gate2064(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2065(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2066(.a(G612), .O(gate202inter7));
  inv1  gate2067(.a(G617), .O(gate202inter8));
  nand2 gate2068(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2069(.a(s_217), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2070(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2071(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2072(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2227(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2228(.a(gate204inter0), .b(s_240), .O(gate204inter1));
  and2  gate2229(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2230(.a(s_240), .O(gate204inter3));
  inv1  gate2231(.a(s_241), .O(gate204inter4));
  nand2 gate2232(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2233(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2234(.a(G607), .O(gate204inter7));
  inv1  gate2235(.a(G617), .O(gate204inter8));
  nand2 gate2236(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2237(.a(s_241), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2238(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2239(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2240(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1765(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1766(.a(gate205inter0), .b(s_174), .O(gate205inter1));
  and2  gate1767(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1768(.a(s_174), .O(gate205inter3));
  inv1  gate1769(.a(s_175), .O(gate205inter4));
  nand2 gate1770(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1771(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1772(.a(G622), .O(gate205inter7));
  inv1  gate1773(.a(G627), .O(gate205inter8));
  nand2 gate1774(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1775(.a(s_175), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1776(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1777(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1778(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate799(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate800(.a(gate206inter0), .b(s_36), .O(gate206inter1));
  and2  gate801(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate802(.a(s_36), .O(gate206inter3));
  inv1  gate803(.a(s_37), .O(gate206inter4));
  nand2 gate804(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate805(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate806(.a(G632), .O(gate206inter7));
  inv1  gate807(.a(G637), .O(gate206inter8));
  nand2 gate808(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate809(.a(s_37), .b(gate206inter3), .O(gate206inter10));
  nor2  gate810(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate811(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate812(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1023(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1024(.a(gate217inter0), .b(s_68), .O(gate217inter1));
  and2  gate1025(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1026(.a(s_68), .O(gate217inter3));
  inv1  gate1027(.a(s_69), .O(gate217inter4));
  nand2 gate1028(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1029(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1030(.a(G622), .O(gate217inter7));
  inv1  gate1031(.a(G678), .O(gate217inter8));
  nand2 gate1032(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1033(.a(s_69), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1034(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1035(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1036(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate687(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate688(.a(gate219inter0), .b(s_20), .O(gate219inter1));
  and2  gate689(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate690(.a(s_20), .O(gate219inter3));
  inv1  gate691(.a(s_21), .O(gate219inter4));
  nand2 gate692(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate693(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate694(.a(G632), .O(gate219inter7));
  inv1  gate695(.a(G681), .O(gate219inter8));
  nand2 gate696(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate697(.a(s_21), .b(gate219inter3), .O(gate219inter10));
  nor2  gate698(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate699(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate700(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate715(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate716(.a(gate228inter0), .b(s_24), .O(gate228inter1));
  and2  gate717(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate718(.a(s_24), .O(gate228inter3));
  inv1  gate719(.a(s_25), .O(gate228inter4));
  nand2 gate720(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate721(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate722(.a(G696), .O(gate228inter7));
  inv1  gate723(.a(G697), .O(gate228inter8));
  nand2 gate724(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate725(.a(s_25), .b(gate228inter3), .O(gate228inter10));
  nor2  gate726(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate727(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate728(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1093(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1094(.a(gate232inter0), .b(s_78), .O(gate232inter1));
  and2  gate1095(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1096(.a(s_78), .O(gate232inter3));
  inv1  gate1097(.a(s_79), .O(gate232inter4));
  nand2 gate1098(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1099(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1100(.a(G704), .O(gate232inter7));
  inv1  gate1101(.a(G705), .O(gate232inter8));
  nand2 gate1102(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1103(.a(s_79), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1104(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1105(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1106(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1149(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1150(.a(gate236inter0), .b(s_86), .O(gate236inter1));
  and2  gate1151(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1152(.a(s_86), .O(gate236inter3));
  inv1  gate1153(.a(s_87), .O(gate236inter4));
  nand2 gate1154(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1155(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1156(.a(G251), .O(gate236inter7));
  inv1  gate1157(.a(G727), .O(gate236inter8));
  nand2 gate1158(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1159(.a(s_87), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1160(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1161(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1162(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate869(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate870(.a(gate237inter0), .b(s_46), .O(gate237inter1));
  and2  gate871(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate872(.a(s_46), .O(gate237inter3));
  inv1  gate873(.a(s_47), .O(gate237inter4));
  nand2 gate874(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate875(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate876(.a(G254), .O(gate237inter7));
  inv1  gate877(.a(G706), .O(gate237inter8));
  nand2 gate878(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate879(.a(s_47), .b(gate237inter3), .O(gate237inter10));
  nor2  gate880(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate881(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate882(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate603(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate604(.a(gate238inter0), .b(s_8), .O(gate238inter1));
  and2  gate605(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate606(.a(s_8), .O(gate238inter3));
  inv1  gate607(.a(s_9), .O(gate238inter4));
  nand2 gate608(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate609(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate610(.a(G257), .O(gate238inter7));
  inv1  gate611(.a(G709), .O(gate238inter8));
  nand2 gate612(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate613(.a(s_9), .b(gate238inter3), .O(gate238inter10));
  nor2  gate614(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate615(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate616(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1919(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1920(.a(gate241inter0), .b(s_196), .O(gate241inter1));
  and2  gate1921(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1922(.a(s_196), .O(gate241inter3));
  inv1  gate1923(.a(s_197), .O(gate241inter4));
  nand2 gate1924(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1925(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1926(.a(G242), .O(gate241inter7));
  inv1  gate1927(.a(G730), .O(gate241inter8));
  nand2 gate1928(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1929(.a(s_197), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1930(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1931(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1932(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate995(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate996(.a(gate244inter0), .b(s_64), .O(gate244inter1));
  and2  gate997(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate998(.a(s_64), .O(gate244inter3));
  inv1  gate999(.a(s_65), .O(gate244inter4));
  nand2 gate1000(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1001(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1002(.a(G721), .O(gate244inter7));
  inv1  gate1003(.a(G733), .O(gate244inter8));
  nand2 gate1004(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1005(.a(s_65), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1006(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1007(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1008(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1415(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1416(.a(gate250inter0), .b(s_124), .O(gate250inter1));
  and2  gate1417(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1418(.a(s_124), .O(gate250inter3));
  inv1  gate1419(.a(s_125), .O(gate250inter4));
  nand2 gate1420(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1421(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1422(.a(G706), .O(gate250inter7));
  inv1  gate1423(.a(G742), .O(gate250inter8));
  nand2 gate1424(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1425(.a(s_125), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1426(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1427(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1428(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1667(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1668(.a(gate258inter0), .b(s_160), .O(gate258inter1));
  and2  gate1669(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1670(.a(s_160), .O(gate258inter3));
  inv1  gate1671(.a(s_161), .O(gate258inter4));
  nand2 gate1672(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1673(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1674(.a(G756), .O(gate258inter7));
  inv1  gate1675(.a(G757), .O(gate258inter8));
  nand2 gate1676(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1677(.a(s_161), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1678(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1679(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1680(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate729(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate730(.a(gate263inter0), .b(s_26), .O(gate263inter1));
  and2  gate731(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate732(.a(s_26), .O(gate263inter3));
  inv1  gate733(.a(s_27), .O(gate263inter4));
  nand2 gate734(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate735(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate736(.a(G766), .O(gate263inter7));
  inv1  gate737(.a(G767), .O(gate263inter8));
  nand2 gate738(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate739(.a(s_27), .b(gate263inter3), .O(gate263inter10));
  nor2  gate740(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate741(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate742(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1261(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1262(.a(gate270inter0), .b(s_102), .O(gate270inter1));
  and2  gate1263(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1264(.a(s_102), .O(gate270inter3));
  inv1  gate1265(.a(s_103), .O(gate270inter4));
  nand2 gate1266(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1267(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1268(.a(G657), .O(gate270inter7));
  inv1  gate1269(.a(G785), .O(gate270inter8));
  nand2 gate1270(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1271(.a(s_103), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1272(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1273(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1274(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2031(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2032(.a(gate271inter0), .b(s_212), .O(gate271inter1));
  and2  gate2033(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2034(.a(s_212), .O(gate271inter3));
  inv1  gate2035(.a(s_213), .O(gate271inter4));
  nand2 gate2036(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2037(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2038(.a(G660), .O(gate271inter7));
  inv1  gate2039(.a(G788), .O(gate271inter8));
  nand2 gate2040(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2041(.a(s_213), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2042(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2043(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2044(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1975(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1976(.a(gate274inter0), .b(s_204), .O(gate274inter1));
  and2  gate1977(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1978(.a(s_204), .O(gate274inter3));
  inv1  gate1979(.a(s_205), .O(gate274inter4));
  nand2 gate1980(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1981(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1982(.a(G770), .O(gate274inter7));
  inv1  gate1983(.a(G794), .O(gate274inter8));
  nand2 gate1984(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1985(.a(s_205), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1986(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1987(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1988(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1863(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1864(.a(gate277inter0), .b(s_188), .O(gate277inter1));
  and2  gate1865(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1866(.a(s_188), .O(gate277inter3));
  inv1  gate1867(.a(s_189), .O(gate277inter4));
  nand2 gate1868(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1869(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1870(.a(G648), .O(gate277inter7));
  inv1  gate1871(.a(G800), .O(gate277inter8));
  nand2 gate1872(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1873(.a(s_189), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1874(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1875(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1876(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2087(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2088(.a(gate282inter0), .b(s_220), .O(gate282inter1));
  and2  gate2089(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2090(.a(s_220), .O(gate282inter3));
  inv1  gate2091(.a(s_221), .O(gate282inter4));
  nand2 gate2092(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2093(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2094(.a(G782), .O(gate282inter7));
  inv1  gate2095(.a(G806), .O(gate282inter8));
  nand2 gate2096(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2097(.a(s_221), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2098(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2099(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2100(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate561(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate562(.a(gate285inter0), .b(s_2), .O(gate285inter1));
  and2  gate563(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate564(.a(s_2), .O(gate285inter3));
  inv1  gate565(.a(s_3), .O(gate285inter4));
  nand2 gate566(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate567(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate568(.a(G660), .O(gate285inter7));
  inv1  gate569(.a(G812), .O(gate285inter8));
  nand2 gate570(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate571(.a(s_3), .b(gate285inter3), .O(gate285inter10));
  nor2  gate572(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate573(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate574(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1989(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1990(.a(gate286inter0), .b(s_206), .O(gate286inter1));
  and2  gate1991(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1992(.a(s_206), .O(gate286inter3));
  inv1  gate1993(.a(s_207), .O(gate286inter4));
  nand2 gate1994(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1995(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1996(.a(G788), .O(gate286inter7));
  inv1  gate1997(.a(G812), .O(gate286inter8));
  nand2 gate1998(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1999(.a(s_207), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2000(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2001(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2002(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1065(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1066(.a(gate288inter0), .b(s_74), .O(gate288inter1));
  and2  gate1067(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1068(.a(s_74), .O(gate288inter3));
  inv1  gate1069(.a(s_75), .O(gate288inter4));
  nand2 gate1070(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1071(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1072(.a(G791), .O(gate288inter7));
  inv1  gate1073(.a(G815), .O(gate288inter8));
  nand2 gate1074(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1075(.a(s_75), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1076(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1077(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1078(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1821(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1822(.a(gate289inter0), .b(s_182), .O(gate289inter1));
  and2  gate1823(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1824(.a(s_182), .O(gate289inter3));
  inv1  gate1825(.a(s_183), .O(gate289inter4));
  nand2 gate1826(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1827(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1828(.a(G818), .O(gate289inter7));
  inv1  gate1829(.a(G819), .O(gate289inter8));
  nand2 gate1830(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1831(.a(s_183), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1832(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1833(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1834(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1695(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1696(.a(gate388inter0), .b(s_164), .O(gate388inter1));
  and2  gate1697(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1698(.a(s_164), .O(gate388inter3));
  inv1  gate1699(.a(s_165), .O(gate388inter4));
  nand2 gate1700(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1701(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1702(.a(G2), .O(gate388inter7));
  inv1  gate1703(.a(G1039), .O(gate388inter8));
  nand2 gate1704(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1705(.a(s_165), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1706(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1707(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1708(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1219(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1220(.a(gate392inter0), .b(s_96), .O(gate392inter1));
  and2  gate1221(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1222(.a(s_96), .O(gate392inter3));
  inv1  gate1223(.a(s_97), .O(gate392inter4));
  nand2 gate1224(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1225(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1226(.a(G6), .O(gate392inter7));
  inv1  gate1227(.a(G1051), .O(gate392inter8));
  nand2 gate1228(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1229(.a(s_97), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1230(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1231(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1232(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1681(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1682(.a(gate393inter0), .b(s_162), .O(gate393inter1));
  and2  gate1683(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1684(.a(s_162), .O(gate393inter3));
  inv1  gate1685(.a(s_163), .O(gate393inter4));
  nand2 gate1686(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1687(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1688(.a(G7), .O(gate393inter7));
  inv1  gate1689(.a(G1054), .O(gate393inter8));
  nand2 gate1690(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1691(.a(s_163), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1692(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1693(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1694(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1555(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1556(.a(gate395inter0), .b(s_144), .O(gate395inter1));
  and2  gate1557(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1558(.a(s_144), .O(gate395inter3));
  inv1  gate1559(.a(s_145), .O(gate395inter4));
  nand2 gate1560(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1561(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1562(.a(G9), .O(gate395inter7));
  inv1  gate1563(.a(G1060), .O(gate395inter8));
  nand2 gate1564(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1565(.a(s_145), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1566(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1567(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1568(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1037(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1038(.a(gate399inter0), .b(s_70), .O(gate399inter1));
  and2  gate1039(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1040(.a(s_70), .O(gate399inter3));
  inv1  gate1041(.a(s_71), .O(gate399inter4));
  nand2 gate1042(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1043(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1044(.a(G13), .O(gate399inter7));
  inv1  gate1045(.a(G1072), .O(gate399inter8));
  nand2 gate1046(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1047(.a(s_71), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1048(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1049(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1050(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate631(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate632(.a(gate400inter0), .b(s_12), .O(gate400inter1));
  and2  gate633(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate634(.a(s_12), .O(gate400inter3));
  inv1  gate635(.a(s_13), .O(gate400inter4));
  nand2 gate636(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate637(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate638(.a(G14), .O(gate400inter7));
  inv1  gate639(.a(G1075), .O(gate400inter8));
  nand2 gate640(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate641(.a(s_13), .b(gate400inter3), .O(gate400inter10));
  nor2  gate642(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate643(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate644(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate589(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate590(.a(gate402inter0), .b(s_6), .O(gate402inter1));
  and2  gate591(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate592(.a(s_6), .O(gate402inter3));
  inv1  gate593(.a(s_7), .O(gate402inter4));
  nand2 gate594(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate595(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate596(.a(G16), .O(gate402inter7));
  inv1  gate597(.a(G1081), .O(gate402inter8));
  nand2 gate598(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate599(.a(s_7), .b(gate402inter3), .O(gate402inter10));
  nor2  gate600(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate601(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate602(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate575(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate576(.a(gate403inter0), .b(s_4), .O(gate403inter1));
  and2  gate577(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate578(.a(s_4), .O(gate403inter3));
  inv1  gate579(.a(s_5), .O(gate403inter4));
  nand2 gate580(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate581(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate582(.a(G17), .O(gate403inter7));
  inv1  gate583(.a(G1084), .O(gate403inter8));
  nand2 gate584(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate585(.a(s_5), .b(gate403inter3), .O(gate403inter10));
  nor2  gate586(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate587(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate588(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1247(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1248(.a(gate409inter0), .b(s_100), .O(gate409inter1));
  and2  gate1249(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1250(.a(s_100), .O(gate409inter3));
  inv1  gate1251(.a(s_101), .O(gate409inter4));
  nand2 gate1252(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1253(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1254(.a(G23), .O(gate409inter7));
  inv1  gate1255(.a(G1102), .O(gate409inter8));
  nand2 gate1256(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1257(.a(s_101), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1258(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1259(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1260(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2143(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2144(.a(gate410inter0), .b(s_228), .O(gate410inter1));
  and2  gate2145(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2146(.a(s_228), .O(gate410inter3));
  inv1  gate2147(.a(s_229), .O(gate410inter4));
  nand2 gate2148(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2149(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2150(.a(G24), .O(gate410inter7));
  inv1  gate2151(.a(G1105), .O(gate410inter8));
  nand2 gate2152(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2153(.a(s_229), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2154(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2155(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2156(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1443(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1444(.a(gate411inter0), .b(s_128), .O(gate411inter1));
  and2  gate1445(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1446(.a(s_128), .O(gate411inter3));
  inv1  gate1447(.a(s_129), .O(gate411inter4));
  nand2 gate1448(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1449(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1450(.a(G25), .O(gate411inter7));
  inv1  gate1451(.a(G1108), .O(gate411inter8));
  nand2 gate1452(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1453(.a(s_129), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1454(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1455(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1456(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1751(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1752(.a(gate412inter0), .b(s_172), .O(gate412inter1));
  and2  gate1753(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1754(.a(s_172), .O(gate412inter3));
  inv1  gate1755(.a(s_173), .O(gate412inter4));
  nand2 gate1756(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1757(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1758(.a(G26), .O(gate412inter7));
  inv1  gate1759(.a(G1111), .O(gate412inter8));
  nand2 gate1760(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1761(.a(s_173), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1762(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1763(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1764(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1849(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1850(.a(gate414inter0), .b(s_186), .O(gate414inter1));
  and2  gate1851(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1852(.a(s_186), .O(gate414inter3));
  inv1  gate1853(.a(s_187), .O(gate414inter4));
  nand2 gate1854(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1855(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1856(.a(G28), .O(gate414inter7));
  inv1  gate1857(.a(G1117), .O(gate414inter8));
  nand2 gate1858(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1859(.a(s_187), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1860(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1861(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1862(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1401(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1402(.a(gate419inter0), .b(s_122), .O(gate419inter1));
  and2  gate1403(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1404(.a(s_122), .O(gate419inter3));
  inv1  gate1405(.a(s_123), .O(gate419inter4));
  nand2 gate1406(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1407(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1408(.a(G1), .O(gate419inter7));
  inv1  gate1409(.a(G1132), .O(gate419inter8));
  nand2 gate1410(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1411(.a(s_123), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1412(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1413(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1414(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1933(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1934(.a(gate420inter0), .b(s_198), .O(gate420inter1));
  and2  gate1935(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1936(.a(s_198), .O(gate420inter3));
  inv1  gate1937(.a(s_199), .O(gate420inter4));
  nand2 gate1938(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1939(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1940(.a(G1036), .O(gate420inter7));
  inv1  gate1941(.a(G1132), .O(gate420inter8));
  nand2 gate1942(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1943(.a(s_199), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1944(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1945(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1946(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate757(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate758(.a(gate423inter0), .b(s_30), .O(gate423inter1));
  and2  gate759(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate760(.a(s_30), .O(gate423inter3));
  inv1  gate761(.a(s_31), .O(gate423inter4));
  nand2 gate762(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate763(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate764(.a(G3), .O(gate423inter7));
  inv1  gate765(.a(G1138), .O(gate423inter8));
  nand2 gate766(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate767(.a(s_31), .b(gate423inter3), .O(gate423inter10));
  nor2  gate768(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate769(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate770(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate785(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate786(.a(gate426inter0), .b(s_34), .O(gate426inter1));
  and2  gate787(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate788(.a(s_34), .O(gate426inter3));
  inv1  gate789(.a(s_35), .O(gate426inter4));
  nand2 gate790(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate791(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate792(.a(G1045), .O(gate426inter7));
  inv1  gate793(.a(G1141), .O(gate426inter8));
  nand2 gate794(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate795(.a(s_35), .b(gate426inter3), .O(gate426inter10));
  nor2  gate796(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate797(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate798(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1317(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1318(.a(gate430inter0), .b(s_110), .O(gate430inter1));
  and2  gate1319(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1320(.a(s_110), .O(gate430inter3));
  inv1  gate1321(.a(s_111), .O(gate430inter4));
  nand2 gate1322(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1323(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1324(.a(G1051), .O(gate430inter7));
  inv1  gate1325(.a(G1147), .O(gate430inter8));
  nand2 gate1326(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1327(.a(s_111), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1328(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1329(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1330(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1191(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1192(.a(gate436inter0), .b(s_92), .O(gate436inter1));
  and2  gate1193(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1194(.a(s_92), .O(gate436inter3));
  inv1  gate1195(.a(s_93), .O(gate436inter4));
  nand2 gate1196(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1197(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1198(.a(G1060), .O(gate436inter7));
  inv1  gate1199(.a(G1156), .O(gate436inter8));
  nand2 gate1200(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1201(.a(s_93), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1202(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1203(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1204(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate967(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate968(.a(gate437inter0), .b(s_60), .O(gate437inter1));
  and2  gate969(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate970(.a(s_60), .O(gate437inter3));
  inv1  gate971(.a(s_61), .O(gate437inter4));
  nand2 gate972(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate973(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate974(.a(G10), .O(gate437inter7));
  inv1  gate975(.a(G1159), .O(gate437inter8));
  nand2 gate976(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate977(.a(s_61), .b(gate437inter3), .O(gate437inter10));
  nor2  gate978(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate979(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate980(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1877(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1878(.a(gate442inter0), .b(s_190), .O(gate442inter1));
  and2  gate1879(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1880(.a(s_190), .O(gate442inter3));
  inv1  gate1881(.a(s_191), .O(gate442inter4));
  nand2 gate1882(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1883(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1884(.a(G1069), .O(gate442inter7));
  inv1  gate1885(.a(G1165), .O(gate442inter8));
  nand2 gate1886(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1887(.a(s_191), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1888(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1889(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1890(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate841(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate842(.a(gate444inter0), .b(s_42), .O(gate444inter1));
  and2  gate843(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate844(.a(s_42), .O(gate444inter3));
  inv1  gate845(.a(s_43), .O(gate444inter4));
  nand2 gate846(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate847(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate848(.a(G1072), .O(gate444inter7));
  inv1  gate849(.a(G1168), .O(gate444inter8));
  nand2 gate850(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate851(.a(s_43), .b(gate444inter3), .O(gate444inter10));
  nor2  gate852(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate853(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate854(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1457(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1458(.a(gate447inter0), .b(s_130), .O(gate447inter1));
  and2  gate1459(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1460(.a(s_130), .O(gate447inter3));
  inv1  gate1461(.a(s_131), .O(gate447inter4));
  nand2 gate1462(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1463(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1464(.a(G15), .O(gate447inter7));
  inv1  gate1465(.a(G1174), .O(gate447inter8));
  nand2 gate1466(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1467(.a(s_131), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1468(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1469(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1470(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2101(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2102(.a(gate448inter0), .b(s_222), .O(gate448inter1));
  and2  gate2103(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2104(.a(s_222), .O(gate448inter3));
  inv1  gate2105(.a(s_223), .O(gate448inter4));
  nand2 gate2106(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2107(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2108(.a(G1078), .O(gate448inter7));
  inv1  gate2109(.a(G1174), .O(gate448inter8));
  nand2 gate2110(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2111(.a(s_223), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2112(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2113(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2114(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate911(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate912(.a(gate450inter0), .b(s_52), .O(gate450inter1));
  and2  gate913(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate914(.a(s_52), .O(gate450inter3));
  inv1  gate915(.a(s_53), .O(gate450inter4));
  nand2 gate916(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate917(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate918(.a(G1081), .O(gate450inter7));
  inv1  gate919(.a(G1177), .O(gate450inter8));
  nand2 gate920(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate921(.a(s_53), .b(gate450inter3), .O(gate450inter10));
  nor2  gate922(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate923(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate924(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1583(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1584(.a(gate453inter0), .b(s_148), .O(gate453inter1));
  and2  gate1585(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1586(.a(s_148), .O(gate453inter3));
  inv1  gate1587(.a(s_149), .O(gate453inter4));
  nand2 gate1588(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1589(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1590(.a(G18), .O(gate453inter7));
  inv1  gate1591(.a(G1183), .O(gate453inter8));
  nand2 gate1592(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1593(.a(s_149), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1594(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1595(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1596(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate897(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate898(.a(gate456inter0), .b(s_50), .O(gate456inter1));
  and2  gate899(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate900(.a(s_50), .O(gate456inter3));
  inv1  gate901(.a(s_51), .O(gate456inter4));
  nand2 gate902(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate903(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate904(.a(G1090), .O(gate456inter7));
  inv1  gate905(.a(G1186), .O(gate456inter8));
  nand2 gate906(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate907(.a(s_51), .b(gate456inter3), .O(gate456inter10));
  nor2  gate908(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate909(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate910(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1541(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1542(.a(gate458inter0), .b(s_142), .O(gate458inter1));
  and2  gate1543(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1544(.a(s_142), .O(gate458inter3));
  inv1  gate1545(.a(s_143), .O(gate458inter4));
  nand2 gate1546(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1547(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1548(.a(G1093), .O(gate458inter7));
  inv1  gate1549(.a(G1189), .O(gate458inter8));
  nand2 gate1550(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1551(.a(s_143), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1552(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1553(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1554(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1807(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1808(.a(gate464inter0), .b(s_180), .O(gate464inter1));
  and2  gate1809(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1810(.a(s_180), .O(gate464inter3));
  inv1  gate1811(.a(s_181), .O(gate464inter4));
  nand2 gate1812(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1813(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1814(.a(G1102), .O(gate464inter7));
  inv1  gate1815(.a(G1198), .O(gate464inter8));
  nand2 gate1816(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1817(.a(s_181), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1818(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1819(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1820(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1961(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1962(.a(gate473inter0), .b(s_202), .O(gate473inter1));
  and2  gate1963(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1964(.a(s_202), .O(gate473inter3));
  inv1  gate1965(.a(s_203), .O(gate473inter4));
  nand2 gate1966(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1967(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1968(.a(G28), .O(gate473inter7));
  inv1  gate1969(.a(G1213), .O(gate473inter8));
  nand2 gate1970(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1971(.a(s_203), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1972(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1973(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1974(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate925(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate926(.a(gate475inter0), .b(s_54), .O(gate475inter1));
  and2  gate927(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate928(.a(s_54), .O(gate475inter3));
  inv1  gate929(.a(s_55), .O(gate475inter4));
  nand2 gate930(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate931(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate932(.a(G29), .O(gate475inter7));
  inv1  gate933(.a(G1216), .O(gate475inter8));
  nand2 gate934(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate935(.a(s_55), .b(gate475inter3), .O(gate475inter10));
  nor2  gate936(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate937(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate938(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1303(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1304(.a(gate476inter0), .b(s_108), .O(gate476inter1));
  and2  gate1305(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1306(.a(s_108), .O(gate476inter3));
  inv1  gate1307(.a(s_109), .O(gate476inter4));
  nand2 gate1308(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1309(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1310(.a(G1120), .O(gate476inter7));
  inv1  gate1311(.a(G1216), .O(gate476inter8));
  nand2 gate1312(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1313(.a(s_109), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1314(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1315(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1316(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1485(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1486(.a(gate477inter0), .b(s_134), .O(gate477inter1));
  and2  gate1487(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1488(.a(s_134), .O(gate477inter3));
  inv1  gate1489(.a(s_135), .O(gate477inter4));
  nand2 gate1490(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1491(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1492(.a(G30), .O(gate477inter7));
  inv1  gate1493(.a(G1219), .O(gate477inter8));
  nand2 gate1494(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1495(.a(s_135), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1496(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1497(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1498(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1793(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1794(.a(gate487inter0), .b(s_178), .O(gate487inter1));
  and2  gate1795(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1796(.a(s_178), .O(gate487inter3));
  inv1  gate1797(.a(s_179), .O(gate487inter4));
  nand2 gate1798(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1799(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1800(.a(G1236), .O(gate487inter7));
  inv1  gate1801(.a(G1237), .O(gate487inter8));
  nand2 gate1802(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1803(.a(s_179), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1804(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1805(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1806(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2157(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2158(.a(gate491inter0), .b(s_230), .O(gate491inter1));
  and2  gate2159(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2160(.a(s_230), .O(gate491inter3));
  inv1  gate2161(.a(s_231), .O(gate491inter4));
  nand2 gate2162(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2163(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2164(.a(G1244), .O(gate491inter7));
  inv1  gate2165(.a(G1245), .O(gate491inter8));
  nand2 gate2166(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2167(.a(s_231), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2168(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2169(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2170(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate743(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate744(.a(gate492inter0), .b(s_28), .O(gate492inter1));
  and2  gate745(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate746(.a(s_28), .O(gate492inter3));
  inv1  gate747(.a(s_29), .O(gate492inter4));
  nand2 gate748(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate749(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate750(.a(G1246), .O(gate492inter7));
  inv1  gate751(.a(G1247), .O(gate492inter8));
  nand2 gate752(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate753(.a(s_29), .b(gate492inter3), .O(gate492inter10));
  nor2  gate754(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate755(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate756(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1107(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1108(.a(gate508inter0), .b(s_80), .O(gate508inter1));
  and2  gate1109(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1110(.a(s_80), .O(gate508inter3));
  inv1  gate1111(.a(s_81), .O(gate508inter4));
  nand2 gate1112(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1113(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1114(.a(G1278), .O(gate508inter7));
  inv1  gate1115(.a(G1279), .O(gate508inter8));
  nand2 gate1116(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1117(.a(s_81), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1118(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1119(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1120(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1891(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1892(.a(gate509inter0), .b(s_192), .O(gate509inter1));
  and2  gate1893(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1894(.a(s_192), .O(gate509inter3));
  inv1  gate1895(.a(s_193), .O(gate509inter4));
  nand2 gate1896(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1897(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1898(.a(G1280), .O(gate509inter7));
  inv1  gate1899(.a(G1281), .O(gate509inter8));
  nand2 gate1900(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1901(.a(s_193), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1902(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1903(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1904(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule