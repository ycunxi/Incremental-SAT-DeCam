module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1667(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1668(.a(gate9inter0), .b(s_160), .O(gate9inter1));
  and2  gate1669(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1670(.a(s_160), .O(gate9inter3));
  inv1  gate1671(.a(s_161), .O(gate9inter4));
  nand2 gate1672(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1673(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1674(.a(G1), .O(gate9inter7));
  inv1  gate1675(.a(G2), .O(gate9inter8));
  nand2 gate1676(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1677(.a(s_161), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1678(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1679(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1680(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2227(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2228(.a(gate11inter0), .b(s_240), .O(gate11inter1));
  and2  gate2229(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2230(.a(s_240), .O(gate11inter3));
  inv1  gate2231(.a(s_241), .O(gate11inter4));
  nand2 gate2232(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2233(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2234(.a(G5), .O(gate11inter7));
  inv1  gate2235(.a(G6), .O(gate11inter8));
  nand2 gate2236(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2237(.a(s_241), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2238(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2239(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2240(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2339(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2340(.a(gate15inter0), .b(s_256), .O(gate15inter1));
  and2  gate2341(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2342(.a(s_256), .O(gate15inter3));
  inv1  gate2343(.a(s_257), .O(gate15inter4));
  nand2 gate2344(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2345(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2346(.a(G13), .O(gate15inter7));
  inv1  gate2347(.a(G14), .O(gate15inter8));
  nand2 gate2348(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2349(.a(s_257), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2350(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2351(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2352(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1275(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1276(.a(gate20inter0), .b(s_104), .O(gate20inter1));
  and2  gate1277(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1278(.a(s_104), .O(gate20inter3));
  inv1  gate1279(.a(s_105), .O(gate20inter4));
  nand2 gate1280(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1281(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1282(.a(G23), .O(gate20inter7));
  inv1  gate1283(.a(G24), .O(gate20inter8));
  nand2 gate1284(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1285(.a(s_105), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1286(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1287(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1288(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1975(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1976(.a(gate21inter0), .b(s_204), .O(gate21inter1));
  and2  gate1977(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1978(.a(s_204), .O(gate21inter3));
  inv1  gate1979(.a(s_205), .O(gate21inter4));
  nand2 gate1980(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1981(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1982(.a(G25), .O(gate21inter7));
  inv1  gate1983(.a(G26), .O(gate21inter8));
  nand2 gate1984(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1985(.a(s_205), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1986(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1987(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1988(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2297(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2298(.a(gate22inter0), .b(s_250), .O(gate22inter1));
  and2  gate2299(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2300(.a(s_250), .O(gate22inter3));
  inv1  gate2301(.a(s_251), .O(gate22inter4));
  nand2 gate2302(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2303(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2304(.a(G27), .O(gate22inter7));
  inv1  gate2305(.a(G28), .O(gate22inter8));
  nand2 gate2306(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2307(.a(s_251), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2308(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2309(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2310(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate659(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate660(.a(gate25inter0), .b(s_16), .O(gate25inter1));
  and2  gate661(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate662(.a(s_16), .O(gate25inter3));
  inv1  gate663(.a(s_17), .O(gate25inter4));
  nand2 gate664(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate665(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate666(.a(G1), .O(gate25inter7));
  inv1  gate667(.a(G5), .O(gate25inter8));
  nand2 gate668(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate669(.a(s_17), .b(gate25inter3), .O(gate25inter10));
  nor2  gate670(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate671(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate672(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1695(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1696(.a(gate27inter0), .b(s_164), .O(gate27inter1));
  and2  gate1697(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1698(.a(s_164), .O(gate27inter3));
  inv1  gate1699(.a(s_165), .O(gate27inter4));
  nand2 gate1700(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1701(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1702(.a(G2), .O(gate27inter7));
  inv1  gate1703(.a(G6), .O(gate27inter8));
  nand2 gate1704(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1705(.a(s_165), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1706(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1707(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1708(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1261(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1262(.a(gate37inter0), .b(s_102), .O(gate37inter1));
  and2  gate1263(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1264(.a(s_102), .O(gate37inter3));
  inv1  gate1265(.a(s_103), .O(gate37inter4));
  nand2 gate1266(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1267(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1268(.a(G19), .O(gate37inter7));
  inv1  gate1269(.a(G23), .O(gate37inter8));
  nand2 gate1270(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1271(.a(s_103), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1272(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1273(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1274(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate827(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate828(.a(gate39inter0), .b(s_40), .O(gate39inter1));
  and2  gate829(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate830(.a(s_40), .O(gate39inter3));
  inv1  gate831(.a(s_41), .O(gate39inter4));
  nand2 gate832(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate833(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate834(.a(G20), .O(gate39inter7));
  inv1  gate835(.a(G24), .O(gate39inter8));
  nand2 gate836(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate837(.a(s_41), .b(gate39inter3), .O(gate39inter10));
  nor2  gate838(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate839(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate840(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1779(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1780(.a(gate46inter0), .b(s_176), .O(gate46inter1));
  and2  gate1781(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1782(.a(s_176), .O(gate46inter3));
  inv1  gate1783(.a(s_177), .O(gate46inter4));
  nand2 gate1784(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1785(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1786(.a(G6), .O(gate46inter7));
  inv1  gate1787(.a(G272), .O(gate46inter8));
  nand2 gate1788(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1789(.a(s_177), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1790(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1791(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1792(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1653(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1654(.a(gate50inter0), .b(s_158), .O(gate50inter1));
  and2  gate1655(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1656(.a(s_158), .O(gate50inter3));
  inv1  gate1657(.a(s_159), .O(gate50inter4));
  nand2 gate1658(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1659(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1660(.a(G10), .O(gate50inter7));
  inv1  gate1661(.a(G278), .O(gate50inter8));
  nand2 gate1662(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1663(.a(s_159), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1664(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1665(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1666(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1121(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1122(.a(gate51inter0), .b(s_82), .O(gate51inter1));
  and2  gate1123(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1124(.a(s_82), .O(gate51inter3));
  inv1  gate1125(.a(s_83), .O(gate51inter4));
  nand2 gate1126(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1127(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1128(.a(G11), .O(gate51inter7));
  inv1  gate1129(.a(G281), .O(gate51inter8));
  nand2 gate1130(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1131(.a(s_83), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1132(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1133(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1134(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate771(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate772(.a(gate54inter0), .b(s_32), .O(gate54inter1));
  and2  gate773(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate774(.a(s_32), .O(gate54inter3));
  inv1  gate775(.a(s_33), .O(gate54inter4));
  nand2 gate776(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate777(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate778(.a(G14), .O(gate54inter7));
  inv1  gate779(.a(G284), .O(gate54inter8));
  nand2 gate780(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate781(.a(s_33), .b(gate54inter3), .O(gate54inter10));
  nor2  gate782(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate783(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate784(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1527(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1528(.a(gate59inter0), .b(s_140), .O(gate59inter1));
  and2  gate1529(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1530(.a(s_140), .O(gate59inter3));
  inv1  gate1531(.a(s_141), .O(gate59inter4));
  nand2 gate1532(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1533(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1534(.a(G19), .O(gate59inter7));
  inv1  gate1535(.a(G293), .O(gate59inter8));
  nand2 gate1536(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1537(.a(s_141), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1538(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1539(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1540(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2381(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2382(.a(gate64inter0), .b(s_262), .O(gate64inter1));
  and2  gate2383(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2384(.a(s_262), .O(gate64inter3));
  inv1  gate2385(.a(s_263), .O(gate64inter4));
  nand2 gate2386(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2387(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2388(.a(G24), .O(gate64inter7));
  inv1  gate2389(.a(G299), .O(gate64inter8));
  nand2 gate2390(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2391(.a(s_263), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2392(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2393(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2394(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate645(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate646(.a(gate66inter0), .b(s_14), .O(gate66inter1));
  and2  gate647(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate648(.a(s_14), .O(gate66inter3));
  inv1  gate649(.a(s_15), .O(gate66inter4));
  nand2 gate650(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate651(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate652(.a(G26), .O(gate66inter7));
  inv1  gate653(.a(G302), .O(gate66inter8));
  nand2 gate654(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate655(.a(s_15), .b(gate66inter3), .O(gate66inter10));
  nor2  gate656(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate657(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate658(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2073(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2074(.a(gate69inter0), .b(s_218), .O(gate69inter1));
  and2  gate2075(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2076(.a(s_218), .O(gate69inter3));
  inv1  gate2077(.a(s_219), .O(gate69inter4));
  nand2 gate2078(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2079(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2080(.a(G29), .O(gate69inter7));
  inv1  gate2081(.a(G308), .O(gate69inter8));
  nand2 gate2082(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2083(.a(s_219), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2084(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2085(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2086(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate589(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate590(.a(gate71inter0), .b(s_6), .O(gate71inter1));
  and2  gate591(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate592(.a(s_6), .O(gate71inter3));
  inv1  gate593(.a(s_7), .O(gate71inter4));
  nand2 gate594(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate595(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate596(.a(G31), .O(gate71inter7));
  inv1  gate597(.a(G311), .O(gate71inter8));
  nand2 gate598(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate599(.a(s_7), .b(gate71inter3), .O(gate71inter10));
  nor2  gate600(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate601(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate602(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate2353(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2354(.a(gate73inter0), .b(s_258), .O(gate73inter1));
  and2  gate2355(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2356(.a(s_258), .O(gate73inter3));
  inv1  gate2357(.a(s_259), .O(gate73inter4));
  nand2 gate2358(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2359(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2360(.a(G1), .O(gate73inter7));
  inv1  gate2361(.a(G314), .O(gate73inter8));
  nand2 gate2362(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2363(.a(s_259), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2364(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2365(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2366(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1135(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1136(.a(gate75inter0), .b(s_84), .O(gate75inter1));
  and2  gate1137(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1138(.a(s_84), .O(gate75inter3));
  inv1  gate1139(.a(s_85), .O(gate75inter4));
  nand2 gate1140(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1141(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1142(.a(G9), .O(gate75inter7));
  inv1  gate1143(.a(G317), .O(gate75inter8));
  nand2 gate1144(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1145(.a(s_85), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1146(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1147(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1148(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate925(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate926(.a(gate76inter0), .b(s_54), .O(gate76inter1));
  and2  gate927(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate928(.a(s_54), .O(gate76inter3));
  inv1  gate929(.a(s_55), .O(gate76inter4));
  nand2 gate930(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate931(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate932(.a(G13), .O(gate76inter7));
  inv1  gate933(.a(G317), .O(gate76inter8));
  nand2 gate934(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate935(.a(s_55), .b(gate76inter3), .O(gate76inter10));
  nor2  gate936(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate937(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate938(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1821(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1822(.a(gate81inter0), .b(s_182), .O(gate81inter1));
  and2  gate1823(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1824(.a(s_182), .O(gate81inter3));
  inv1  gate1825(.a(s_183), .O(gate81inter4));
  nand2 gate1826(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1827(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1828(.a(G3), .O(gate81inter7));
  inv1  gate1829(.a(G326), .O(gate81inter8));
  nand2 gate1830(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1831(.a(s_183), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1832(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1833(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1834(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate2255(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2256(.a(gate83inter0), .b(s_244), .O(gate83inter1));
  and2  gate2257(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2258(.a(s_244), .O(gate83inter3));
  inv1  gate2259(.a(s_245), .O(gate83inter4));
  nand2 gate2260(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2261(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2262(.a(G11), .O(gate83inter7));
  inv1  gate2263(.a(G329), .O(gate83inter8));
  nand2 gate2264(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2265(.a(s_245), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2266(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2267(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2268(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1933(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1934(.a(gate86inter0), .b(s_198), .O(gate86inter1));
  and2  gate1935(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1936(.a(s_198), .O(gate86inter3));
  inv1  gate1937(.a(s_199), .O(gate86inter4));
  nand2 gate1938(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1939(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1940(.a(G8), .O(gate86inter7));
  inv1  gate1941(.a(G332), .O(gate86inter8));
  nand2 gate1942(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1943(.a(s_199), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1944(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1945(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1946(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate855(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate856(.a(gate87inter0), .b(s_44), .O(gate87inter1));
  and2  gate857(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate858(.a(s_44), .O(gate87inter3));
  inv1  gate859(.a(s_45), .O(gate87inter4));
  nand2 gate860(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate861(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate862(.a(G12), .O(gate87inter7));
  inv1  gate863(.a(G335), .O(gate87inter8));
  nand2 gate864(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate865(.a(s_45), .b(gate87inter3), .O(gate87inter10));
  nor2  gate866(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate867(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate868(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2409(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2410(.a(gate91inter0), .b(s_266), .O(gate91inter1));
  and2  gate2411(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2412(.a(s_266), .O(gate91inter3));
  inv1  gate2413(.a(s_267), .O(gate91inter4));
  nand2 gate2414(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2415(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2416(.a(G25), .O(gate91inter7));
  inv1  gate2417(.a(G341), .O(gate91inter8));
  nand2 gate2418(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2419(.a(s_267), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2420(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2421(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2422(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate897(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate898(.a(gate94inter0), .b(s_50), .O(gate94inter1));
  and2  gate899(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate900(.a(s_50), .O(gate94inter3));
  inv1  gate901(.a(s_51), .O(gate94inter4));
  nand2 gate902(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate903(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate904(.a(G22), .O(gate94inter7));
  inv1  gate905(.a(G344), .O(gate94inter8));
  nand2 gate906(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate907(.a(s_51), .b(gate94inter3), .O(gate94inter10));
  nor2  gate908(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate909(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate910(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate869(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate870(.a(gate102inter0), .b(s_46), .O(gate102inter1));
  and2  gate871(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate872(.a(s_46), .O(gate102inter3));
  inv1  gate873(.a(s_47), .O(gate102inter4));
  nand2 gate874(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate875(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate876(.a(G24), .O(gate102inter7));
  inv1  gate877(.a(G356), .O(gate102inter8));
  nand2 gate878(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate879(.a(s_47), .b(gate102inter3), .O(gate102inter10));
  nor2  gate880(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate881(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate882(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2143(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2144(.a(gate108inter0), .b(s_228), .O(gate108inter1));
  and2  gate2145(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2146(.a(s_228), .O(gate108inter3));
  inv1  gate2147(.a(s_229), .O(gate108inter4));
  nand2 gate2148(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2149(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2150(.a(G368), .O(gate108inter7));
  inv1  gate2151(.a(G369), .O(gate108inter8));
  nand2 gate2152(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2153(.a(s_229), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2154(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2155(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2156(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1723(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1724(.a(gate109inter0), .b(s_168), .O(gate109inter1));
  and2  gate1725(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1726(.a(s_168), .O(gate109inter3));
  inv1  gate1727(.a(s_169), .O(gate109inter4));
  nand2 gate1728(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1729(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1730(.a(G370), .O(gate109inter7));
  inv1  gate1731(.a(G371), .O(gate109inter8));
  nand2 gate1732(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1733(.a(s_169), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1734(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1735(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1736(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate575(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate576(.a(gate111inter0), .b(s_4), .O(gate111inter1));
  and2  gate577(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate578(.a(s_4), .O(gate111inter3));
  inv1  gate579(.a(s_5), .O(gate111inter4));
  nand2 gate580(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate581(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate582(.a(G374), .O(gate111inter7));
  inv1  gate583(.a(G375), .O(gate111inter8));
  nand2 gate584(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate585(.a(s_5), .b(gate111inter3), .O(gate111inter10));
  nor2  gate586(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate587(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate588(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1233(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1234(.a(gate118inter0), .b(s_98), .O(gate118inter1));
  and2  gate1235(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1236(.a(s_98), .O(gate118inter3));
  inv1  gate1237(.a(s_99), .O(gate118inter4));
  nand2 gate1238(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1239(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1240(.a(G388), .O(gate118inter7));
  inv1  gate1241(.a(G389), .O(gate118inter8));
  nand2 gate1242(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1243(.a(s_99), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1244(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1245(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1246(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1499(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1500(.a(gate119inter0), .b(s_136), .O(gate119inter1));
  and2  gate1501(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1502(.a(s_136), .O(gate119inter3));
  inv1  gate1503(.a(s_137), .O(gate119inter4));
  nand2 gate1504(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1505(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1506(.a(G390), .O(gate119inter7));
  inv1  gate1507(.a(G391), .O(gate119inter8));
  nand2 gate1508(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1509(.a(s_137), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1510(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1511(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1512(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1345(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1346(.a(gate125inter0), .b(s_114), .O(gate125inter1));
  and2  gate1347(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1348(.a(s_114), .O(gate125inter3));
  inv1  gate1349(.a(s_115), .O(gate125inter4));
  nand2 gate1350(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1351(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1352(.a(G402), .O(gate125inter7));
  inv1  gate1353(.a(G403), .O(gate125inter8));
  nand2 gate1354(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1355(.a(s_115), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1356(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1357(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1358(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1387(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1388(.a(gate126inter0), .b(s_120), .O(gate126inter1));
  and2  gate1389(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1390(.a(s_120), .O(gate126inter3));
  inv1  gate1391(.a(s_121), .O(gate126inter4));
  nand2 gate1392(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1393(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1394(.a(G404), .O(gate126inter7));
  inv1  gate1395(.a(G405), .O(gate126inter8));
  nand2 gate1396(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1397(.a(s_121), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1398(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1399(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1400(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate799(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate800(.a(gate127inter0), .b(s_36), .O(gate127inter1));
  and2  gate801(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate802(.a(s_36), .O(gate127inter3));
  inv1  gate803(.a(s_37), .O(gate127inter4));
  nand2 gate804(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate805(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate806(.a(G406), .O(gate127inter7));
  inv1  gate807(.a(G407), .O(gate127inter8));
  nand2 gate808(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate809(.a(s_37), .b(gate127inter3), .O(gate127inter10));
  nor2  gate810(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate811(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate812(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1737(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1738(.a(gate132inter0), .b(s_170), .O(gate132inter1));
  and2  gate1739(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1740(.a(s_170), .O(gate132inter3));
  inv1  gate1741(.a(s_171), .O(gate132inter4));
  nand2 gate1742(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1743(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1744(.a(G416), .O(gate132inter7));
  inv1  gate1745(.a(G417), .O(gate132inter8));
  nand2 gate1746(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1747(.a(s_171), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1748(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1749(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1750(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1219(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1220(.a(gate133inter0), .b(s_96), .O(gate133inter1));
  and2  gate1221(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1222(.a(s_96), .O(gate133inter3));
  inv1  gate1223(.a(s_97), .O(gate133inter4));
  nand2 gate1224(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1225(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1226(.a(G418), .O(gate133inter7));
  inv1  gate1227(.a(G419), .O(gate133inter8));
  nand2 gate1228(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1229(.a(s_97), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1230(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1231(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1232(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1765(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1766(.a(gate136inter0), .b(s_174), .O(gate136inter1));
  and2  gate1767(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1768(.a(s_174), .O(gate136inter3));
  inv1  gate1769(.a(s_175), .O(gate136inter4));
  nand2 gate1770(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1771(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1772(.a(G424), .O(gate136inter7));
  inv1  gate1773(.a(G425), .O(gate136inter8));
  nand2 gate1774(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1775(.a(s_175), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1776(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1777(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1778(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1457(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1458(.a(gate137inter0), .b(s_130), .O(gate137inter1));
  and2  gate1459(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1460(.a(s_130), .O(gate137inter3));
  inv1  gate1461(.a(s_131), .O(gate137inter4));
  nand2 gate1462(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1463(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1464(.a(G426), .O(gate137inter7));
  inv1  gate1465(.a(G429), .O(gate137inter8));
  nand2 gate1466(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1467(.a(s_131), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1468(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1469(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1470(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1863(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1864(.a(gate140inter0), .b(s_188), .O(gate140inter1));
  and2  gate1865(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1866(.a(s_188), .O(gate140inter3));
  inv1  gate1867(.a(s_189), .O(gate140inter4));
  nand2 gate1868(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1869(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1870(.a(G444), .O(gate140inter7));
  inv1  gate1871(.a(G447), .O(gate140inter8));
  nand2 gate1872(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1873(.a(s_189), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1874(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1875(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1876(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1247(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1248(.a(gate141inter0), .b(s_100), .O(gate141inter1));
  and2  gate1249(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1250(.a(s_100), .O(gate141inter3));
  inv1  gate1251(.a(s_101), .O(gate141inter4));
  nand2 gate1252(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1253(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1254(.a(G450), .O(gate141inter7));
  inv1  gate1255(.a(G453), .O(gate141inter8));
  nand2 gate1256(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1257(.a(s_101), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1258(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1259(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1260(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate911(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate912(.a(gate143inter0), .b(s_52), .O(gate143inter1));
  and2  gate913(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate914(.a(s_52), .O(gate143inter3));
  inv1  gate915(.a(s_53), .O(gate143inter4));
  nand2 gate916(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate917(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate918(.a(G462), .O(gate143inter7));
  inv1  gate919(.a(G465), .O(gate143inter8));
  nand2 gate920(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate921(.a(s_53), .b(gate143inter3), .O(gate143inter10));
  nor2  gate922(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate923(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate924(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1079(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1080(.a(gate147inter0), .b(s_76), .O(gate147inter1));
  and2  gate1081(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1082(.a(s_76), .O(gate147inter3));
  inv1  gate1083(.a(s_77), .O(gate147inter4));
  nand2 gate1084(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1085(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1086(.a(G486), .O(gate147inter7));
  inv1  gate1087(.a(G489), .O(gate147inter8));
  nand2 gate1088(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1089(.a(s_77), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1090(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1091(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1092(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate785(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate786(.a(gate148inter0), .b(s_34), .O(gate148inter1));
  and2  gate787(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate788(.a(s_34), .O(gate148inter3));
  inv1  gate789(.a(s_35), .O(gate148inter4));
  nand2 gate790(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate791(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate792(.a(G492), .O(gate148inter7));
  inv1  gate793(.a(G495), .O(gate148inter8));
  nand2 gate794(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate795(.a(s_35), .b(gate148inter3), .O(gate148inter10));
  nor2  gate796(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate797(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate798(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate967(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate968(.a(gate150inter0), .b(s_60), .O(gate150inter1));
  and2  gate969(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate970(.a(s_60), .O(gate150inter3));
  inv1  gate971(.a(s_61), .O(gate150inter4));
  nand2 gate972(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate973(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate974(.a(G504), .O(gate150inter7));
  inv1  gate975(.a(G507), .O(gate150inter8));
  nand2 gate976(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate977(.a(s_61), .b(gate150inter3), .O(gate150inter10));
  nor2  gate978(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate979(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate980(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2115(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2116(.a(gate156inter0), .b(s_224), .O(gate156inter1));
  and2  gate2117(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2118(.a(s_224), .O(gate156inter3));
  inv1  gate2119(.a(s_225), .O(gate156inter4));
  nand2 gate2120(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2121(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2122(.a(G435), .O(gate156inter7));
  inv1  gate2123(.a(G525), .O(gate156inter8));
  nand2 gate2124(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2125(.a(s_225), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2126(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2127(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2128(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1359(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1360(.a(gate162inter0), .b(s_116), .O(gate162inter1));
  and2  gate1361(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1362(.a(s_116), .O(gate162inter3));
  inv1  gate1363(.a(s_117), .O(gate162inter4));
  nand2 gate1364(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1365(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1366(.a(G453), .O(gate162inter7));
  inv1  gate1367(.a(G534), .O(gate162inter8));
  nand2 gate1368(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1369(.a(s_117), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1370(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1371(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1372(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2045(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2046(.a(gate167inter0), .b(s_214), .O(gate167inter1));
  and2  gate2047(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2048(.a(s_214), .O(gate167inter3));
  inv1  gate2049(.a(s_215), .O(gate167inter4));
  nand2 gate2050(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2051(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2052(.a(G468), .O(gate167inter7));
  inv1  gate2053(.a(G543), .O(gate167inter8));
  nand2 gate2054(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2055(.a(s_215), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2056(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2057(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2058(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1891(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1892(.a(gate179inter0), .b(s_192), .O(gate179inter1));
  and2  gate1893(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1894(.a(s_192), .O(gate179inter3));
  inv1  gate1895(.a(s_193), .O(gate179inter4));
  nand2 gate1896(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1897(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1898(.a(G504), .O(gate179inter7));
  inv1  gate1899(.a(G561), .O(gate179inter8));
  nand2 gate1900(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1901(.a(s_193), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1902(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1903(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1904(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate701(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate702(.a(gate180inter0), .b(s_22), .O(gate180inter1));
  and2  gate703(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate704(.a(s_22), .O(gate180inter3));
  inv1  gate705(.a(s_23), .O(gate180inter4));
  nand2 gate706(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate707(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate708(.a(G507), .O(gate180inter7));
  inv1  gate709(.a(G561), .O(gate180inter8));
  nand2 gate710(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate711(.a(s_23), .b(gate180inter3), .O(gate180inter10));
  nor2  gate712(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate713(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate714(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate687(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate688(.a(gate181inter0), .b(s_20), .O(gate181inter1));
  and2  gate689(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate690(.a(s_20), .O(gate181inter3));
  inv1  gate691(.a(s_21), .O(gate181inter4));
  nand2 gate692(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate693(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate694(.a(G510), .O(gate181inter7));
  inv1  gate695(.a(G564), .O(gate181inter8));
  nand2 gate696(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate697(.a(s_21), .b(gate181inter3), .O(gate181inter10));
  nor2  gate698(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate699(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate700(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1569(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1570(.a(gate186inter0), .b(s_146), .O(gate186inter1));
  and2  gate1571(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1572(.a(s_146), .O(gate186inter3));
  inv1  gate1573(.a(s_147), .O(gate186inter4));
  nand2 gate1574(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1575(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1576(.a(G572), .O(gate186inter7));
  inv1  gate1577(.a(G573), .O(gate186inter8));
  nand2 gate1578(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1579(.a(s_147), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1580(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1581(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1582(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1331(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1332(.a(gate188inter0), .b(s_112), .O(gate188inter1));
  and2  gate1333(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1334(.a(s_112), .O(gate188inter3));
  inv1  gate1335(.a(s_113), .O(gate188inter4));
  nand2 gate1336(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1337(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1338(.a(G576), .O(gate188inter7));
  inv1  gate1339(.a(G577), .O(gate188inter8));
  nand2 gate1340(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1341(.a(s_113), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1342(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1343(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1344(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1037(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1038(.a(gate190inter0), .b(s_70), .O(gate190inter1));
  and2  gate1039(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1040(.a(s_70), .O(gate190inter3));
  inv1  gate1041(.a(s_71), .O(gate190inter4));
  nand2 gate1042(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1043(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1044(.a(G580), .O(gate190inter7));
  inv1  gate1045(.a(G581), .O(gate190inter8));
  nand2 gate1046(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1047(.a(s_71), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1048(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1049(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1050(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1443(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1444(.a(gate194inter0), .b(s_128), .O(gate194inter1));
  and2  gate1445(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1446(.a(s_128), .O(gate194inter3));
  inv1  gate1447(.a(s_129), .O(gate194inter4));
  nand2 gate1448(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1449(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1450(.a(G588), .O(gate194inter7));
  inv1  gate1451(.a(G589), .O(gate194inter8));
  nand2 gate1452(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1453(.a(s_129), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1454(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1455(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1456(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2171(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2172(.a(gate195inter0), .b(s_232), .O(gate195inter1));
  and2  gate2173(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2174(.a(s_232), .O(gate195inter3));
  inv1  gate2175(.a(s_233), .O(gate195inter4));
  nand2 gate2176(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2177(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2178(.a(G590), .O(gate195inter7));
  inv1  gate2179(.a(G591), .O(gate195inter8));
  nand2 gate2180(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2181(.a(s_233), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2182(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2183(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2184(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate743(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate744(.a(gate196inter0), .b(s_28), .O(gate196inter1));
  and2  gate745(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate746(.a(s_28), .O(gate196inter3));
  inv1  gate747(.a(s_29), .O(gate196inter4));
  nand2 gate748(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate749(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate750(.a(G592), .O(gate196inter7));
  inv1  gate751(.a(G593), .O(gate196inter8));
  nand2 gate752(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate753(.a(s_29), .b(gate196inter3), .O(gate196inter10));
  nor2  gate754(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate755(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate756(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1625(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1626(.a(gate197inter0), .b(s_154), .O(gate197inter1));
  and2  gate1627(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1628(.a(s_154), .O(gate197inter3));
  inv1  gate1629(.a(s_155), .O(gate197inter4));
  nand2 gate1630(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1631(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1632(.a(G594), .O(gate197inter7));
  inv1  gate1633(.a(G595), .O(gate197inter8));
  nand2 gate1634(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1635(.a(s_155), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1636(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1637(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1638(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1191(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1192(.a(gate199inter0), .b(s_92), .O(gate199inter1));
  and2  gate1193(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1194(.a(s_92), .O(gate199inter3));
  inv1  gate1195(.a(s_93), .O(gate199inter4));
  nand2 gate1196(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1197(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1198(.a(G598), .O(gate199inter7));
  inv1  gate1199(.a(G599), .O(gate199inter8));
  nand2 gate1200(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1201(.a(s_93), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1202(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1203(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1204(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1583(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1584(.a(gate201inter0), .b(s_148), .O(gate201inter1));
  and2  gate1585(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1586(.a(s_148), .O(gate201inter3));
  inv1  gate1587(.a(s_149), .O(gate201inter4));
  nand2 gate1588(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1589(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1590(.a(G602), .O(gate201inter7));
  inv1  gate1591(.a(G607), .O(gate201inter8));
  nand2 gate1592(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1593(.a(s_149), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1594(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1595(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1596(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1905(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1906(.a(gate202inter0), .b(s_194), .O(gate202inter1));
  and2  gate1907(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1908(.a(s_194), .O(gate202inter3));
  inv1  gate1909(.a(s_195), .O(gate202inter4));
  nand2 gate1910(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1911(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1912(.a(G612), .O(gate202inter7));
  inv1  gate1913(.a(G617), .O(gate202inter8));
  nand2 gate1914(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1915(.a(s_195), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1916(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1917(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1918(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate939(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate940(.a(gate204inter0), .b(s_56), .O(gate204inter1));
  and2  gate941(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate942(.a(s_56), .O(gate204inter3));
  inv1  gate943(.a(s_57), .O(gate204inter4));
  nand2 gate944(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate945(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate946(.a(G607), .O(gate204inter7));
  inv1  gate947(.a(G617), .O(gate204inter8));
  nand2 gate948(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate949(.a(s_57), .b(gate204inter3), .O(gate204inter10));
  nor2  gate950(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate951(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate952(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate2059(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2060(.a(gate205inter0), .b(s_216), .O(gate205inter1));
  and2  gate2061(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2062(.a(s_216), .O(gate205inter3));
  inv1  gate2063(.a(s_217), .O(gate205inter4));
  nand2 gate2064(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2065(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2066(.a(G622), .O(gate205inter7));
  inv1  gate2067(.a(G627), .O(gate205inter8));
  nand2 gate2068(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2069(.a(s_217), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2070(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2071(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2072(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2311(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2312(.a(gate207inter0), .b(s_252), .O(gate207inter1));
  and2  gate2313(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2314(.a(s_252), .O(gate207inter3));
  inv1  gate2315(.a(s_253), .O(gate207inter4));
  nand2 gate2316(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2317(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2318(.a(G622), .O(gate207inter7));
  inv1  gate2319(.a(G632), .O(gate207inter8));
  nand2 gate2320(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2321(.a(s_253), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2322(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2323(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2324(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1751(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1752(.a(gate211inter0), .b(s_172), .O(gate211inter1));
  and2  gate1753(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1754(.a(s_172), .O(gate211inter3));
  inv1  gate1755(.a(s_173), .O(gate211inter4));
  nand2 gate1756(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1757(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1758(.a(G612), .O(gate211inter7));
  inv1  gate1759(.a(G669), .O(gate211inter8));
  nand2 gate1760(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1761(.a(s_173), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1762(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1763(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1764(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2031(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2032(.a(gate212inter0), .b(s_212), .O(gate212inter1));
  and2  gate2033(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2034(.a(s_212), .O(gate212inter3));
  inv1  gate2035(.a(s_213), .O(gate212inter4));
  nand2 gate2036(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2037(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2038(.a(G617), .O(gate212inter7));
  inv1  gate2039(.a(G669), .O(gate212inter8));
  nand2 gate2040(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2041(.a(s_213), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2042(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2043(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2044(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1835(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1836(.a(gate215inter0), .b(s_184), .O(gate215inter1));
  and2  gate1837(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1838(.a(s_184), .O(gate215inter3));
  inv1  gate1839(.a(s_185), .O(gate215inter4));
  nand2 gate1840(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1841(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1842(.a(G607), .O(gate215inter7));
  inv1  gate1843(.a(G675), .O(gate215inter8));
  nand2 gate1844(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1845(.a(s_185), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1846(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1847(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1848(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate673(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate674(.a(gate218inter0), .b(s_18), .O(gate218inter1));
  and2  gate675(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate676(.a(s_18), .O(gate218inter3));
  inv1  gate677(.a(s_19), .O(gate218inter4));
  nand2 gate678(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate679(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate680(.a(G627), .O(gate218inter7));
  inv1  gate681(.a(G678), .O(gate218inter8));
  nand2 gate682(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate683(.a(s_19), .b(gate218inter3), .O(gate218inter10));
  nor2  gate684(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate685(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate686(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1793(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1794(.a(gate219inter0), .b(s_178), .O(gate219inter1));
  and2  gate1795(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1796(.a(s_178), .O(gate219inter3));
  inv1  gate1797(.a(s_179), .O(gate219inter4));
  nand2 gate1798(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1799(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1800(.a(G632), .O(gate219inter7));
  inv1  gate1801(.a(G681), .O(gate219inter8));
  nand2 gate1802(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1803(.a(s_179), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1804(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1805(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1806(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate841(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate842(.a(gate222inter0), .b(s_42), .O(gate222inter1));
  and2  gate843(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate844(.a(s_42), .O(gate222inter3));
  inv1  gate845(.a(s_43), .O(gate222inter4));
  nand2 gate846(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate847(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate848(.a(G632), .O(gate222inter7));
  inv1  gate849(.a(G684), .O(gate222inter8));
  nand2 gate850(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate851(.a(s_43), .b(gate222inter3), .O(gate222inter10));
  nor2  gate852(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate853(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate854(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2185(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2186(.a(gate223inter0), .b(s_234), .O(gate223inter1));
  and2  gate2187(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2188(.a(s_234), .O(gate223inter3));
  inv1  gate2189(.a(s_235), .O(gate223inter4));
  nand2 gate2190(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2191(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2192(.a(G627), .O(gate223inter7));
  inv1  gate2193(.a(G687), .O(gate223inter8));
  nand2 gate2194(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2195(.a(s_235), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2196(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2197(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2198(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1947(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1948(.a(gate224inter0), .b(s_200), .O(gate224inter1));
  and2  gate1949(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1950(.a(s_200), .O(gate224inter3));
  inv1  gate1951(.a(s_201), .O(gate224inter4));
  nand2 gate1952(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1953(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1954(.a(G637), .O(gate224inter7));
  inv1  gate1955(.a(G687), .O(gate224inter8));
  nand2 gate1956(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1957(.a(s_201), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1958(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1959(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1960(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1541(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1542(.a(gate230inter0), .b(s_142), .O(gate230inter1));
  and2  gate1543(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1544(.a(s_142), .O(gate230inter3));
  inv1  gate1545(.a(s_143), .O(gate230inter4));
  nand2 gate1546(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1547(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1548(.a(G700), .O(gate230inter7));
  inv1  gate1549(.a(G701), .O(gate230inter8));
  nand2 gate1550(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1551(.a(s_143), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1552(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1553(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1554(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2283(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2284(.a(gate231inter0), .b(s_248), .O(gate231inter1));
  and2  gate2285(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2286(.a(s_248), .O(gate231inter3));
  inv1  gate2287(.a(s_249), .O(gate231inter4));
  nand2 gate2288(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2289(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2290(.a(G702), .O(gate231inter7));
  inv1  gate2291(.a(G703), .O(gate231inter8));
  nand2 gate2292(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2293(.a(s_249), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2294(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2295(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2296(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2395(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2396(.a(gate233inter0), .b(s_264), .O(gate233inter1));
  and2  gate2397(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2398(.a(s_264), .O(gate233inter3));
  inv1  gate2399(.a(s_265), .O(gate233inter4));
  nand2 gate2400(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2401(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2402(.a(G242), .O(gate233inter7));
  inv1  gate2403(.a(G718), .O(gate233inter8));
  nand2 gate2404(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2405(.a(s_265), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2406(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2407(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2408(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1177(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1178(.a(gate245inter0), .b(s_90), .O(gate245inter1));
  and2  gate1179(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1180(.a(s_90), .O(gate245inter3));
  inv1  gate1181(.a(s_91), .O(gate245inter4));
  nand2 gate1182(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1183(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1184(.a(G248), .O(gate245inter7));
  inv1  gate1185(.a(G736), .O(gate245inter8));
  nand2 gate1186(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1187(.a(s_91), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1188(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1189(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1190(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2101(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2102(.a(gate252inter0), .b(s_222), .O(gate252inter1));
  and2  gate2103(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2104(.a(s_222), .O(gate252inter3));
  inv1  gate2105(.a(s_223), .O(gate252inter4));
  nand2 gate2106(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2107(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2108(.a(G709), .O(gate252inter7));
  inv1  gate2109(.a(G745), .O(gate252inter8));
  nand2 gate2110(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2111(.a(s_223), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2112(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2113(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2114(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1877(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1878(.a(gate257inter0), .b(s_190), .O(gate257inter1));
  and2  gate1879(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1880(.a(s_190), .O(gate257inter3));
  inv1  gate1881(.a(s_191), .O(gate257inter4));
  nand2 gate1882(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1883(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1884(.a(G754), .O(gate257inter7));
  inv1  gate1885(.a(G755), .O(gate257inter8));
  nand2 gate1886(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1887(.a(s_191), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1888(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1889(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1890(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1961(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1962(.a(gate261inter0), .b(s_202), .O(gate261inter1));
  and2  gate1963(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1964(.a(s_202), .O(gate261inter3));
  inv1  gate1965(.a(s_203), .O(gate261inter4));
  nand2 gate1966(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1967(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1968(.a(G762), .O(gate261inter7));
  inv1  gate1969(.a(G763), .O(gate261inter8));
  nand2 gate1970(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1971(.a(s_203), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1972(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1973(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1974(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2213(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2214(.a(gate262inter0), .b(s_238), .O(gate262inter1));
  and2  gate2215(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2216(.a(s_238), .O(gate262inter3));
  inv1  gate2217(.a(s_239), .O(gate262inter4));
  nand2 gate2218(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2219(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2220(.a(G764), .O(gate262inter7));
  inv1  gate2221(.a(G765), .O(gate262inter8));
  nand2 gate2222(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2223(.a(s_239), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2224(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2225(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2226(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1023(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1024(.a(gate267inter0), .b(s_68), .O(gate267inter1));
  and2  gate1025(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1026(.a(s_68), .O(gate267inter3));
  inv1  gate1027(.a(s_69), .O(gate267inter4));
  nand2 gate1028(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1029(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1030(.a(G648), .O(gate267inter7));
  inv1  gate1031(.a(G776), .O(gate267inter8));
  nand2 gate1032(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1033(.a(s_69), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1034(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1035(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1036(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate953(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate954(.a(gate274inter0), .b(s_58), .O(gate274inter1));
  and2  gate955(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate956(.a(s_58), .O(gate274inter3));
  inv1  gate957(.a(s_59), .O(gate274inter4));
  nand2 gate958(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate959(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate960(.a(G770), .O(gate274inter7));
  inv1  gate961(.a(G794), .O(gate274inter8));
  nand2 gate962(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate963(.a(s_59), .b(gate274inter3), .O(gate274inter10));
  nor2  gate964(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate965(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate966(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1009(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1010(.a(gate279inter0), .b(s_66), .O(gate279inter1));
  and2  gate1011(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1012(.a(s_66), .O(gate279inter3));
  inv1  gate1013(.a(s_67), .O(gate279inter4));
  nand2 gate1014(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1015(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1016(.a(G651), .O(gate279inter7));
  inv1  gate1017(.a(G803), .O(gate279inter8));
  nand2 gate1018(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1019(.a(s_67), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1020(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1021(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1022(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2129(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2130(.a(gate283inter0), .b(s_226), .O(gate283inter1));
  and2  gate2131(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2132(.a(s_226), .O(gate283inter3));
  inv1  gate2133(.a(s_227), .O(gate283inter4));
  nand2 gate2134(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2135(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2136(.a(G657), .O(gate283inter7));
  inv1  gate2137(.a(G809), .O(gate283inter8));
  nand2 gate2138(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2139(.a(s_227), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2140(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2141(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2142(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2423(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2424(.a(gate289inter0), .b(s_268), .O(gate289inter1));
  and2  gate2425(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2426(.a(s_268), .O(gate289inter3));
  inv1  gate2427(.a(s_269), .O(gate289inter4));
  nand2 gate2428(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2429(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2430(.a(G818), .O(gate289inter7));
  inv1  gate2431(.a(G819), .O(gate289inter8));
  nand2 gate2432(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2433(.a(s_269), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2434(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2435(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2436(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate757(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate758(.a(gate292inter0), .b(s_30), .O(gate292inter1));
  and2  gate759(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate760(.a(s_30), .O(gate292inter3));
  inv1  gate761(.a(s_31), .O(gate292inter4));
  nand2 gate762(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate763(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate764(.a(G824), .O(gate292inter7));
  inv1  gate765(.a(G825), .O(gate292inter8));
  nand2 gate766(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate767(.a(s_31), .b(gate292inter3), .O(gate292inter10));
  nor2  gate768(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate769(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate770(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate883(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate884(.a(gate294inter0), .b(s_48), .O(gate294inter1));
  and2  gate885(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate886(.a(s_48), .O(gate294inter3));
  inv1  gate887(.a(s_49), .O(gate294inter4));
  nand2 gate888(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate889(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate890(.a(G832), .O(gate294inter7));
  inv1  gate891(.a(G833), .O(gate294inter8));
  nand2 gate892(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate893(.a(s_49), .b(gate294inter3), .O(gate294inter10));
  nor2  gate894(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate895(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate896(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2157(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2158(.a(gate296inter0), .b(s_230), .O(gate296inter1));
  and2  gate2159(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2160(.a(s_230), .O(gate296inter3));
  inv1  gate2161(.a(s_231), .O(gate296inter4));
  nand2 gate2162(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2163(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2164(.a(G826), .O(gate296inter7));
  inv1  gate2165(.a(G827), .O(gate296inter8));
  nand2 gate2166(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2167(.a(s_231), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2168(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2169(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2170(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1989(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1990(.a(gate389inter0), .b(s_206), .O(gate389inter1));
  and2  gate1991(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1992(.a(s_206), .O(gate389inter3));
  inv1  gate1993(.a(s_207), .O(gate389inter4));
  nand2 gate1994(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1995(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1996(.a(G3), .O(gate389inter7));
  inv1  gate1997(.a(G1042), .O(gate389inter8));
  nand2 gate1998(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1999(.a(s_207), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2000(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2001(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2002(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1513(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1514(.a(gate392inter0), .b(s_138), .O(gate392inter1));
  and2  gate1515(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1516(.a(s_138), .O(gate392inter3));
  inv1  gate1517(.a(s_139), .O(gate392inter4));
  nand2 gate1518(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1519(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1520(.a(G6), .O(gate392inter7));
  inv1  gate1521(.a(G1051), .O(gate392inter8));
  nand2 gate1522(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1523(.a(s_139), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1524(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1525(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1526(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1051(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1052(.a(gate393inter0), .b(s_72), .O(gate393inter1));
  and2  gate1053(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1054(.a(s_72), .O(gate393inter3));
  inv1  gate1055(.a(s_73), .O(gate393inter4));
  nand2 gate1056(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1057(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1058(.a(G7), .O(gate393inter7));
  inv1  gate1059(.a(G1054), .O(gate393inter8));
  nand2 gate1060(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1061(.a(s_73), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1062(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1063(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1064(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate547(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate548(.a(gate399inter0), .b(s_0), .O(gate399inter1));
  and2  gate549(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate550(.a(s_0), .O(gate399inter3));
  inv1  gate551(.a(s_1), .O(gate399inter4));
  nand2 gate552(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate553(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate554(.a(G13), .O(gate399inter7));
  inv1  gate555(.a(G1072), .O(gate399inter8));
  nand2 gate556(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate557(.a(s_1), .b(gate399inter3), .O(gate399inter10));
  nor2  gate558(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate559(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate560(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2003(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2004(.a(gate402inter0), .b(s_208), .O(gate402inter1));
  and2  gate2005(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2006(.a(s_208), .O(gate402inter3));
  inv1  gate2007(.a(s_209), .O(gate402inter4));
  nand2 gate2008(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2009(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2010(.a(G16), .O(gate402inter7));
  inv1  gate2011(.a(G1081), .O(gate402inter8));
  nand2 gate2012(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2013(.a(s_209), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2014(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2015(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2016(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate617(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate618(.a(gate403inter0), .b(s_10), .O(gate403inter1));
  and2  gate619(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate620(.a(s_10), .O(gate403inter3));
  inv1  gate621(.a(s_11), .O(gate403inter4));
  nand2 gate622(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate623(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate624(.a(G17), .O(gate403inter7));
  inv1  gate625(.a(G1084), .O(gate403inter8));
  nand2 gate626(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate627(.a(s_11), .b(gate403inter3), .O(gate403inter10));
  nor2  gate628(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate629(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate630(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1163(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1164(.a(gate404inter0), .b(s_88), .O(gate404inter1));
  and2  gate1165(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1166(.a(s_88), .O(gate404inter3));
  inv1  gate1167(.a(s_89), .O(gate404inter4));
  nand2 gate1168(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1169(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1170(.a(G18), .O(gate404inter7));
  inv1  gate1171(.a(G1087), .O(gate404inter8));
  nand2 gate1172(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1173(.a(s_89), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1174(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1175(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1176(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1709(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1710(.a(gate405inter0), .b(s_166), .O(gate405inter1));
  and2  gate1711(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1712(.a(s_166), .O(gate405inter3));
  inv1  gate1713(.a(s_167), .O(gate405inter4));
  nand2 gate1714(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1715(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1716(.a(G19), .O(gate405inter7));
  inv1  gate1717(.a(G1090), .O(gate405inter8));
  nand2 gate1718(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1719(.a(s_167), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1720(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1721(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1722(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1401(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1402(.a(gate409inter0), .b(s_122), .O(gate409inter1));
  and2  gate1403(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1404(.a(s_122), .O(gate409inter3));
  inv1  gate1405(.a(s_123), .O(gate409inter4));
  nand2 gate1406(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1407(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1408(.a(G23), .O(gate409inter7));
  inv1  gate1409(.a(G1102), .O(gate409inter8));
  nand2 gate1410(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1411(.a(s_123), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1412(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1413(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1414(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1149(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1150(.a(gate411inter0), .b(s_86), .O(gate411inter1));
  and2  gate1151(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1152(.a(s_86), .O(gate411inter3));
  inv1  gate1153(.a(s_87), .O(gate411inter4));
  nand2 gate1154(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1155(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1156(.a(G25), .O(gate411inter7));
  inv1  gate1157(.a(G1108), .O(gate411inter8));
  nand2 gate1158(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1159(.a(s_87), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1160(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1161(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1162(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1555(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1556(.a(gate417inter0), .b(s_144), .O(gate417inter1));
  and2  gate1557(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1558(.a(s_144), .O(gate417inter3));
  inv1  gate1559(.a(s_145), .O(gate417inter4));
  nand2 gate1560(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1561(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1562(.a(G31), .O(gate417inter7));
  inv1  gate1563(.a(G1126), .O(gate417inter8));
  nand2 gate1564(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1565(.a(s_145), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1566(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1567(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1568(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate813(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate814(.a(gate418inter0), .b(s_38), .O(gate418inter1));
  and2  gate815(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate816(.a(s_38), .O(gate418inter3));
  inv1  gate817(.a(s_39), .O(gate418inter4));
  nand2 gate818(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate819(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate820(.a(G32), .O(gate418inter7));
  inv1  gate821(.a(G1129), .O(gate418inter8));
  nand2 gate822(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate823(.a(s_39), .b(gate418inter3), .O(gate418inter10));
  nor2  gate824(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate825(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate826(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1471(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1472(.a(gate422inter0), .b(s_132), .O(gate422inter1));
  and2  gate1473(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1474(.a(s_132), .O(gate422inter3));
  inv1  gate1475(.a(s_133), .O(gate422inter4));
  nand2 gate1476(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1477(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1478(.a(G1039), .O(gate422inter7));
  inv1  gate1479(.a(G1135), .O(gate422inter8));
  nand2 gate1480(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1481(.a(s_133), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1482(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1483(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1484(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2325(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2326(.a(gate429inter0), .b(s_254), .O(gate429inter1));
  and2  gate2327(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2328(.a(s_254), .O(gate429inter3));
  inv1  gate2329(.a(s_255), .O(gate429inter4));
  nand2 gate2330(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2331(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2332(.a(G6), .O(gate429inter7));
  inv1  gate2333(.a(G1147), .O(gate429inter8));
  nand2 gate2334(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2335(.a(s_255), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2336(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2337(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2338(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1485(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1486(.a(gate437inter0), .b(s_134), .O(gate437inter1));
  and2  gate1487(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1488(.a(s_134), .O(gate437inter3));
  inv1  gate1489(.a(s_135), .O(gate437inter4));
  nand2 gate1490(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1491(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1492(.a(G10), .O(gate437inter7));
  inv1  gate1493(.a(G1159), .O(gate437inter8));
  nand2 gate1494(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1495(.a(s_135), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1496(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1497(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1498(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate715(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate716(.a(gate440inter0), .b(s_24), .O(gate440inter1));
  and2  gate717(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate718(.a(s_24), .O(gate440inter3));
  inv1  gate719(.a(s_25), .O(gate440inter4));
  nand2 gate720(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate721(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate722(.a(G1066), .O(gate440inter7));
  inv1  gate723(.a(G1162), .O(gate440inter8));
  nand2 gate724(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate725(.a(s_25), .b(gate440inter3), .O(gate440inter10));
  nor2  gate726(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate727(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate728(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate561(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate562(.a(gate441inter0), .b(s_2), .O(gate441inter1));
  and2  gate563(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate564(.a(s_2), .O(gate441inter3));
  inv1  gate565(.a(s_3), .O(gate441inter4));
  nand2 gate566(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate567(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate568(.a(G12), .O(gate441inter7));
  inv1  gate569(.a(G1165), .O(gate441inter8));
  nand2 gate570(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate571(.a(s_3), .b(gate441inter3), .O(gate441inter10));
  nor2  gate572(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate573(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate574(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate729(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate730(.a(gate442inter0), .b(s_26), .O(gate442inter1));
  and2  gate731(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate732(.a(s_26), .O(gate442inter3));
  inv1  gate733(.a(s_27), .O(gate442inter4));
  nand2 gate734(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate735(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate736(.a(G1069), .O(gate442inter7));
  inv1  gate737(.a(G1165), .O(gate442inter8));
  nand2 gate738(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate739(.a(s_27), .b(gate442inter3), .O(gate442inter10));
  nor2  gate740(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate741(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate742(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1205(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1206(.a(gate448inter0), .b(s_94), .O(gate448inter1));
  and2  gate1207(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1208(.a(s_94), .O(gate448inter3));
  inv1  gate1209(.a(s_95), .O(gate448inter4));
  nand2 gate1210(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1211(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1212(.a(G1078), .O(gate448inter7));
  inv1  gate1213(.a(G1174), .O(gate448inter8));
  nand2 gate1214(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1215(.a(s_95), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1216(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1217(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1218(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1681(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1682(.a(gate453inter0), .b(s_162), .O(gate453inter1));
  and2  gate1683(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1684(.a(s_162), .O(gate453inter3));
  inv1  gate1685(.a(s_163), .O(gate453inter4));
  nand2 gate1686(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1687(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1688(.a(G18), .O(gate453inter7));
  inv1  gate1689(.a(G1183), .O(gate453inter8));
  nand2 gate1690(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1691(.a(s_163), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1692(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1693(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1694(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate995(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate996(.a(gate454inter0), .b(s_64), .O(gate454inter1));
  and2  gate997(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate998(.a(s_64), .O(gate454inter3));
  inv1  gate999(.a(s_65), .O(gate454inter4));
  nand2 gate1000(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1001(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1002(.a(G1087), .O(gate454inter7));
  inv1  gate1003(.a(G1183), .O(gate454inter8));
  nand2 gate1004(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1005(.a(s_65), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1006(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1007(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1008(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1639(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1640(.a(gate455inter0), .b(s_156), .O(gate455inter1));
  and2  gate1641(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1642(.a(s_156), .O(gate455inter3));
  inv1  gate1643(.a(s_157), .O(gate455inter4));
  nand2 gate1644(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1645(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1646(.a(G19), .O(gate455inter7));
  inv1  gate1647(.a(G1186), .O(gate455inter8));
  nand2 gate1648(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1649(.a(s_157), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1650(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1651(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1652(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2199(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2200(.a(gate458inter0), .b(s_236), .O(gate458inter1));
  and2  gate2201(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2202(.a(s_236), .O(gate458inter3));
  inv1  gate2203(.a(s_237), .O(gate458inter4));
  nand2 gate2204(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2205(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2206(.a(G1093), .O(gate458inter7));
  inv1  gate2207(.a(G1189), .O(gate458inter8));
  nand2 gate2208(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2209(.a(s_237), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2210(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2211(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2212(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2241(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2242(.a(gate460inter0), .b(s_242), .O(gate460inter1));
  and2  gate2243(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2244(.a(s_242), .O(gate460inter3));
  inv1  gate2245(.a(s_243), .O(gate460inter4));
  nand2 gate2246(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2247(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2248(.a(G1096), .O(gate460inter7));
  inv1  gate2249(.a(G1192), .O(gate460inter8));
  nand2 gate2250(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2251(.a(s_243), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2252(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2253(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2254(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1597(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1598(.a(gate463inter0), .b(s_150), .O(gate463inter1));
  and2  gate1599(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1600(.a(s_150), .O(gate463inter3));
  inv1  gate1601(.a(s_151), .O(gate463inter4));
  nand2 gate1602(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1603(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1604(.a(G23), .O(gate463inter7));
  inv1  gate1605(.a(G1198), .O(gate463inter8));
  nand2 gate1606(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1607(.a(s_151), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1608(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1609(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1610(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate981(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate982(.a(gate469inter0), .b(s_62), .O(gate469inter1));
  and2  gate983(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate984(.a(s_62), .O(gate469inter3));
  inv1  gate985(.a(s_63), .O(gate469inter4));
  nand2 gate986(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate987(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate988(.a(G26), .O(gate469inter7));
  inv1  gate989(.a(G1207), .O(gate469inter8));
  nand2 gate990(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate991(.a(s_63), .b(gate469inter3), .O(gate469inter10));
  nor2  gate992(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate993(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate994(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2367(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2368(.a(gate471inter0), .b(s_260), .O(gate471inter1));
  and2  gate2369(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2370(.a(s_260), .O(gate471inter3));
  inv1  gate2371(.a(s_261), .O(gate471inter4));
  nand2 gate2372(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2373(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2374(.a(G27), .O(gate471inter7));
  inv1  gate2375(.a(G1210), .O(gate471inter8));
  nand2 gate2376(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2377(.a(s_261), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2378(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2379(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2380(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate631(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate632(.a(gate472inter0), .b(s_12), .O(gate472inter1));
  and2  gate633(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate634(.a(s_12), .O(gate472inter3));
  inv1  gate635(.a(s_13), .O(gate472inter4));
  nand2 gate636(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate637(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate638(.a(G1114), .O(gate472inter7));
  inv1  gate639(.a(G1210), .O(gate472inter8));
  nand2 gate640(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate641(.a(s_13), .b(gate472inter3), .O(gate472inter10));
  nor2  gate642(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate643(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate644(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1373(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1374(.a(gate474inter0), .b(s_118), .O(gate474inter1));
  and2  gate1375(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1376(.a(s_118), .O(gate474inter3));
  inv1  gate1377(.a(s_119), .O(gate474inter4));
  nand2 gate1378(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1379(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1380(.a(G1117), .O(gate474inter7));
  inv1  gate1381(.a(G1213), .O(gate474inter8));
  nand2 gate1382(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1383(.a(s_119), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1384(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1385(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1386(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1093(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1094(.a(gate475inter0), .b(s_78), .O(gate475inter1));
  and2  gate1095(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1096(.a(s_78), .O(gate475inter3));
  inv1  gate1097(.a(s_79), .O(gate475inter4));
  nand2 gate1098(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1099(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1100(.a(G29), .O(gate475inter7));
  inv1  gate1101(.a(G1216), .O(gate475inter8));
  nand2 gate1102(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1103(.a(s_79), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1104(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1105(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1106(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1919(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1920(.a(gate479inter0), .b(s_196), .O(gate479inter1));
  and2  gate1921(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1922(.a(s_196), .O(gate479inter3));
  inv1  gate1923(.a(s_197), .O(gate479inter4));
  nand2 gate1924(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1925(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1926(.a(G31), .O(gate479inter7));
  inv1  gate1927(.a(G1222), .O(gate479inter8));
  nand2 gate1928(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1929(.a(s_197), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1930(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1931(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1932(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1303(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1304(.a(gate480inter0), .b(s_108), .O(gate480inter1));
  and2  gate1305(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1306(.a(s_108), .O(gate480inter3));
  inv1  gate1307(.a(s_109), .O(gate480inter4));
  nand2 gate1308(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1309(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1310(.a(G1126), .O(gate480inter7));
  inv1  gate1311(.a(G1222), .O(gate480inter8));
  nand2 gate1312(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1313(.a(s_109), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1314(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1315(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1316(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1415(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1416(.a(gate481inter0), .b(s_124), .O(gate481inter1));
  and2  gate1417(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1418(.a(s_124), .O(gate481inter3));
  inv1  gate1419(.a(s_125), .O(gate481inter4));
  nand2 gate1420(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1421(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1422(.a(G32), .O(gate481inter7));
  inv1  gate1423(.a(G1225), .O(gate481inter8));
  nand2 gate1424(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1425(.a(s_125), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1426(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1427(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1428(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate603(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate604(.a(gate483inter0), .b(s_8), .O(gate483inter1));
  and2  gate605(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate606(.a(s_8), .O(gate483inter3));
  inv1  gate607(.a(s_9), .O(gate483inter4));
  nand2 gate608(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate609(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate610(.a(G1228), .O(gate483inter7));
  inv1  gate611(.a(G1229), .O(gate483inter8));
  nand2 gate612(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate613(.a(s_9), .b(gate483inter3), .O(gate483inter10));
  nor2  gate614(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate615(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate616(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1317(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1318(.a(gate484inter0), .b(s_110), .O(gate484inter1));
  and2  gate1319(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1320(.a(s_110), .O(gate484inter3));
  inv1  gate1321(.a(s_111), .O(gate484inter4));
  nand2 gate1322(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1323(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1324(.a(G1230), .O(gate484inter7));
  inv1  gate1325(.a(G1231), .O(gate484inter8));
  nand2 gate1326(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1327(.a(s_111), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1328(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1329(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1330(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2437(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2438(.a(gate485inter0), .b(s_270), .O(gate485inter1));
  and2  gate2439(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2440(.a(s_270), .O(gate485inter3));
  inv1  gate2441(.a(s_271), .O(gate485inter4));
  nand2 gate2442(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2443(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2444(.a(G1232), .O(gate485inter7));
  inv1  gate2445(.a(G1233), .O(gate485inter8));
  nand2 gate2446(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2447(.a(s_271), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2448(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2449(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2450(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1289(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1290(.a(gate487inter0), .b(s_106), .O(gate487inter1));
  and2  gate1291(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1292(.a(s_106), .O(gate487inter3));
  inv1  gate1293(.a(s_107), .O(gate487inter4));
  nand2 gate1294(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1295(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1296(.a(G1236), .O(gate487inter7));
  inv1  gate1297(.a(G1237), .O(gate487inter8));
  nand2 gate1298(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1299(.a(s_107), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1300(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1301(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1302(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2017(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2018(.a(gate488inter0), .b(s_210), .O(gate488inter1));
  and2  gate2019(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2020(.a(s_210), .O(gate488inter3));
  inv1  gate2021(.a(s_211), .O(gate488inter4));
  nand2 gate2022(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2023(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2024(.a(G1238), .O(gate488inter7));
  inv1  gate2025(.a(G1239), .O(gate488inter8));
  nand2 gate2026(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2027(.a(s_211), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2028(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2029(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2030(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2087(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2088(.a(gate490inter0), .b(s_220), .O(gate490inter1));
  and2  gate2089(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2090(.a(s_220), .O(gate490inter3));
  inv1  gate2091(.a(s_221), .O(gate490inter4));
  nand2 gate2092(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2093(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2094(.a(G1242), .O(gate490inter7));
  inv1  gate2095(.a(G1243), .O(gate490inter8));
  nand2 gate2096(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2097(.a(s_221), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2098(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2099(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2100(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1107(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1108(.a(gate491inter0), .b(s_80), .O(gate491inter1));
  and2  gate1109(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1110(.a(s_80), .O(gate491inter3));
  inv1  gate1111(.a(s_81), .O(gate491inter4));
  nand2 gate1112(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1113(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1114(.a(G1244), .O(gate491inter7));
  inv1  gate1115(.a(G1245), .O(gate491inter8));
  nand2 gate1116(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1117(.a(s_81), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1118(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1119(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1120(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1065(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1066(.a(gate495inter0), .b(s_74), .O(gate495inter1));
  and2  gate1067(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1068(.a(s_74), .O(gate495inter3));
  inv1  gate1069(.a(s_75), .O(gate495inter4));
  nand2 gate1070(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1071(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1072(.a(G1252), .O(gate495inter7));
  inv1  gate1073(.a(G1253), .O(gate495inter8));
  nand2 gate1074(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1075(.a(s_75), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1076(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1077(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1078(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate1849(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1850(.a(gate496inter0), .b(s_186), .O(gate496inter1));
  and2  gate1851(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1852(.a(s_186), .O(gate496inter3));
  inv1  gate1853(.a(s_187), .O(gate496inter4));
  nand2 gate1854(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1855(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1856(.a(G1254), .O(gate496inter7));
  inv1  gate1857(.a(G1255), .O(gate496inter8));
  nand2 gate1858(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1859(.a(s_187), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1860(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1861(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1862(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1429(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1430(.a(gate497inter0), .b(s_126), .O(gate497inter1));
  and2  gate1431(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1432(.a(s_126), .O(gate497inter3));
  inv1  gate1433(.a(s_127), .O(gate497inter4));
  nand2 gate1434(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1435(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1436(.a(G1256), .O(gate497inter7));
  inv1  gate1437(.a(G1257), .O(gate497inter8));
  nand2 gate1438(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1439(.a(s_127), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1440(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1441(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1442(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1611(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1612(.a(gate500inter0), .b(s_152), .O(gate500inter1));
  and2  gate1613(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1614(.a(s_152), .O(gate500inter3));
  inv1  gate1615(.a(s_153), .O(gate500inter4));
  nand2 gate1616(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1617(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1618(.a(G1262), .O(gate500inter7));
  inv1  gate1619(.a(G1263), .O(gate500inter8));
  nand2 gate1620(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1621(.a(s_153), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1622(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1623(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1624(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1807(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1808(.a(gate502inter0), .b(s_180), .O(gate502inter1));
  and2  gate1809(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1810(.a(s_180), .O(gate502inter3));
  inv1  gate1811(.a(s_181), .O(gate502inter4));
  nand2 gate1812(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1813(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1814(.a(G1266), .O(gate502inter7));
  inv1  gate1815(.a(G1267), .O(gate502inter8));
  nand2 gate1816(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1817(.a(s_181), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1818(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1819(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1820(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2269(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2270(.a(gate510inter0), .b(s_246), .O(gate510inter1));
  and2  gate2271(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2272(.a(s_246), .O(gate510inter3));
  inv1  gate2273(.a(s_247), .O(gate510inter4));
  nand2 gate2274(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2275(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2276(.a(G1282), .O(gate510inter7));
  inv1  gate2277(.a(G1283), .O(gate510inter8));
  nand2 gate2278(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2279(.a(s_247), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2280(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2281(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2282(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule