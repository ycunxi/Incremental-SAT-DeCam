module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1401(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1402(.a(gate10inter0), .b(s_122), .O(gate10inter1));
  and2  gate1403(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1404(.a(s_122), .O(gate10inter3));
  inv1  gate1405(.a(s_123), .O(gate10inter4));
  nand2 gate1406(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1407(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1408(.a(G3), .O(gate10inter7));
  inv1  gate1409(.a(G4), .O(gate10inter8));
  nand2 gate1410(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1411(.a(s_123), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1412(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1413(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1414(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate575(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate576(.a(gate12inter0), .b(s_4), .O(gate12inter1));
  and2  gate577(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate578(.a(s_4), .O(gate12inter3));
  inv1  gate579(.a(s_5), .O(gate12inter4));
  nand2 gate580(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate581(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate582(.a(G7), .O(gate12inter7));
  inv1  gate583(.a(G8), .O(gate12inter8));
  nand2 gate584(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate585(.a(s_5), .b(gate12inter3), .O(gate12inter10));
  nor2  gate586(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate587(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate588(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate799(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate800(.a(gate20inter0), .b(s_36), .O(gate20inter1));
  and2  gate801(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate802(.a(s_36), .O(gate20inter3));
  inv1  gate803(.a(s_37), .O(gate20inter4));
  nand2 gate804(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate805(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate806(.a(G23), .O(gate20inter7));
  inv1  gate807(.a(G24), .O(gate20inter8));
  nand2 gate808(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate809(.a(s_37), .b(gate20inter3), .O(gate20inter10));
  nor2  gate810(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate811(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate812(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1177(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1178(.a(gate28inter0), .b(s_90), .O(gate28inter1));
  and2  gate1179(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1180(.a(s_90), .O(gate28inter3));
  inv1  gate1181(.a(s_91), .O(gate28inter4));
  nand2 gate1182(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1183(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1184(.a(G10), .O(gate28inter7));
  inv1  gate1185(.a(G14), .O(gate28inter8));
  nand2 gate1186(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1187(.a(s_91), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1188(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1189(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1190(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate701(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate702(.a(gate31inter0), .b(s_22), .O(gate31inter1));
  and2  gate703(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate704(.a(s_22), .O(gate31inter3));
  inv1  gate705(.a(s_23), .O(gate31inter4));
  nand2 gate706(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate707(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate708(.a(G4), .O(gate31inter7));
  inv1  gate709(.a(G8), .O(gate31inter8));
  nand2 gate710(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate711(.a(s_23), .b(gate31inter3), .O(gate31inter10));
  nor2  gate712(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate713(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate714(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate883(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate884(.a(gate44inter0), .b(s_48), .O(gate44inter1));
  and2  gate885(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate886(.a(s_48), .O(gate44inter3));
  inv1  gate887(.a(s_49), .O(gate44inter4));
  nand2 gate888(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate889(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate890(.a(G4), .O(gate44inter7));
  inv1  gate891(.a(G269), .O(gate44inter8));
  nand2 gate892(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate893(.a(s_49), .b(gate44inter3), .O(gate44inter10));
  nor2  gate894(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate895(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate896(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1121(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1122(.a(gate56inter0), .b(s_82), .O(gate56inter1));
  and2  gate1123(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1124(.a(s_82), .O(gate56inter3));
  inv1  gate1125(.a(s_83), .O(gate56inter4));
  nand2 gate1126(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1127(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1128(.a(G16), .O(gate56inter7));
  inv1  gate1129(.a(G287), .O(gate56inter8));
  nand2 gate1130(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1131(.a(s_83), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1132(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1133(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1134(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1191(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1192(.a(gate57inter0), .b(s_92), .O(gate57inter1));
  and2  gate1193(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1194(.a(s_92), .O(gate57inter3));
  inv1  gate1195(.a(s_93), .O(gate57inter4));
  nand2 gate1196(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1197(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1198(.a(G17), .O(gate57inter7));
  inv1  gate1199(.a(G290), .O(gate57inter8));
  nand2 gate1200(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1201(.a(s_93), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1202(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1203(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1204(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate673(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate674(.a(gate69inter0), .b(s_18), .O(gate69inter1));
  and2  gate675(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate676(.a(s_18), .O(gate69inter3));
  inv1  gate677(.a(s_19), .O(gate69inter4));
  nand2 gate678(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate679(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate680(.a(G29), .O(gate69inter7));
  inv1  gate681(.a(G308), .O(gate69inter8));
  nand2 gate682(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate683(.a(s_19), .b(gate69inter3), .O(gate69inter10));
  nor2  gate684(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate685(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate686(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1387(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1388(.a(gate75inter0), .b(s_120), .O(gate75inter1));
  and2  gate1389(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1390(.a(s_120), .O(gate75inter3));
  inv1  gate1391(.a(s_121), .O(gate75inter4));
  nand2 gate1392(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1393(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1394(.a(G9), .O(gate75inter7));
  inv1  gate1395(.a(G317), .O(gate75inter8));
  nand2 gate1396(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1397(.a(s_121), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1398(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1399(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1400(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1023(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1024(.a(gate79inter0), .b(s_68), .O(gate79inter1));
  and2  gate1025(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1026(.a(s_68), .O(gate79inter3));
  inv1  gate1027(.a(s_69), .O(gate79inter4));
  nand2 gate1028(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1029(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1030(.a(G10), .O(gate79inter7));
  inv1  gate1031(.a(G323), .O(gate79inter8));
  nand2 gate1032(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1033(.a(s_69), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1034(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1035(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1036(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate659(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate660(.a(gate80inter0), .b(s_16), .O(gate80inter1));
  and2  gate661(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate662(.a(s_16), .O(gate80inter3));
  inv1  gate663(.a(s_17), .O(gate80inter4));
  nand2 gate664(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate665(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate666(.a(G14), .O(gate80inter7));
  inv1  gate667(.a(G323), .O(gate80inter8));
  nand2 gate668(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate669(.a(s_17), .b(gate80inter3), .O(gate80inter10));
  nor2  gate670(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate671(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate672(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate757(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate758(.a(gate86inter0), .b(s_30), .O(gate86inter1));
  and2  gate759(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate760(.a(s_30), .O(gate86inter3));
  inv1  gate761(.a(s_31), .O(gate86inter4));
  nand2 gate762(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate763(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate764(.a(G8), .O(gate86inter7));
  inv1  gate765(.a(G332), .O(gate86inter8));
  nand2 gate766(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate767(.a(s_31), .b(gate86inter3), .O(gate86inter10));
  nor2  gate768(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate769(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate770(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate743(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate744(.a(gate103inter0), .b(s_28), .O(gate103inter1));
  and2  gate745(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate746(.a(s_28), .O(gate103inter3));
  inv1  gate747(.a(s_29), .O(gate103inter4));
  nand2 gate748(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate749(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate750(.a(G28), .O(gate103inter7));
  inv1  gate751(.a(G359), .O(gate103inter8));
  nand2 gate752(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate753(.a(s_29), .b(gate103inter3), .O(gate103inter10));
  nor2  gate754(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate755(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate756(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate561(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate562(.a(gate115inter0), .b(s_2), .O(gate115inter1));
  and2  gate563(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate564(.a(s_2), .O(gate115inter3));
  inv1  gate565(.a(s_3), .O(gate115inter4));
  nand2 gate566(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate567(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate568(.a(G382), .O(gate115inter7));
  inv1  gate569(.a(G383), .O(gate115inter8));
  nand2 gate570(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate571(.a(s_3), .b(gate115inter3), .O(gate115inter10));
  nor2  gate572(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate573(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate574(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate855(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate856(.a(gate135inter0), .b(s_44), .O(gate135inter1));
  and2  gate857(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate858(.a(s_44), .O(gate135inter3));
  inv1  gate859(.a(s_45), .O(gate135inter4));
  nand2 gate860(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate861(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate862(.a(G422), .O(gate135inter7));
  inv1  gate863(.a(G423), .O(gate135inter8));
  nand2 gate864(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate865(.a(s_45), .b(gate135inter3), .O(gate135inter10));
  nor2  gate866(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate867(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate868(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1037(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1038(.a(gate137inter0), .b(s_70), .O(gate137inter1));
  and2  gate1039(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1040(.a(s_70), .O(gate137inter3));
  inv1  gate1041(.a(s_71), .O(gate137inter4));
  nand2 gate1042(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1043(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1044(.a(G426), .O(gate137inter7));
  inv1  gate1045(.a(G429), .O(gate137inter8));
  nand2 gate1046(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1047(.a(s_71), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1048(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1049(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1050(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate911(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate912(.a(gate164inter0), .b(s_52), .O(gate164inter1));
  and2  gate913(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate914(.a(s_52), .O(gate164inter3));
  inv1  gate915(.a(s_53), .O(gate164inter4));
  nand2 gate916(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate917(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate918(.a(G459), .O(gate164inter7));
  inv1  gate919(.a(G537), .O(gate164inter8));
  nand2 gate920(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate921(.a(s_53), .b(gate164inter3), .O(gate164inter10));
  nor2  gate922(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate923(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate924(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1331(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1332(.a(gate167inter0), .b(s_112), .O(gate167inter1));
  and2  gate1333(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1334(.a(s_112), .O(gate167inter3));
  inv1  gate1335(.a(s_113), .O(gate167inter4));
  nand2 gate1336(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1337(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1338(.a(G468), .O(gate167inter7));
  inv1  gate1339(.a(G543), .O(gate167inter8));
  nand2 gate1340(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1341(.a(s_113), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1342(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1343(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1344(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate771(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate772(.a(gate169inter0), .b(s_32), .O(gate169inter1));
  and2  gate773(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate774(.a(s_32), .O(gate169inter3));
  inv1  gate775(.a(s_33), .O(gate169inter4));
  nand2 gate776(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate777(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate778(.a(G474), .O(gate169inter7));
  inv1  gate779(.a(G546), .O(gate169inter8));
  nand2 gate780(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate781(.a(s_33), .b(gate169inter3), .O(gate169inter10));
  nor2  gate782(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate783(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate784(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate785(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate786(.a(gate170inter0), .b(s_34), .O(gate170inter1));
  and2  gate787(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate788(.a(s_34), .O(gate170inter3));
  inv1  gate789(.a(s_35), .O(gate170inter4));
  nand2 gate790(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate791(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate792(.a(G477), .O(gate170inter7));
  inv1  gate793(.a(G546), .O(gate170inter8));
  nand2 gate794(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate795(.a(s_35), .b(gate170inter3), .O(gate170inter10));
  nor2  gate796(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate797(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate798(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1359(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1360(.a(gate177inter0), .b(s_116), .O(gate177inter1));
  and2  gate1361(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1362(.a(s_116), .O(gate177inter3));
  inv1  gate1363(.a(s_117), .O(gate177inter4));
  nand2 gate1364(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1365(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1366(.a(G498), .O(gate177inter7));
  inv1  gate1367(.a(G558), .O(gate177inter8));
  nand2 gate1368(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1369(.a(s_117), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1370(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1371(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1372(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1093(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1094(.a(gate179inter0), .b(s_78), .O(gate179inter1));
  and2  gate1095(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1096(.a(s_78), .O(gate179inter3));
  inv1  gate1097(.a(s_79), .O(gate179inter4));
  nand2 gate1098(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1099(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1100(.a(G504), .O(gate179inter7));
  inv1  gate1101(.a(G561), .O(gate179inter8));
  nand2 gate1102(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1103(.a(s_79), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1104(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1105(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1106(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate589(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate590(.a(gate181inter0), .b(s_6), .O(gate181inter1));
  and2  gate591(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate592(.a(s_6), .O(gate181inter3));
  inv1  gate593(.a(s_7), .O(gate181inter4));
  nand2 gate594(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate595(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate596(.a(G510), .O(gate181inter7));
  inv1  gate597(.a(G564), .O(gate181inter8));
  nand2 gate598(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate599(.a(s_7), .b(gate181inter3), .O(gate181inter10));
  nor2  gate600(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate601(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate602(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1233(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1234(.a(gate183inter0), .b(s_98), .O(gate183inter1));
  and2  gate1235(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1236(.a(s_98), .O(gate183inter3));
  inv1  gate1237(.a(s_99), .O(gate183inter4));
  nand2 gate1238(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1239(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1240(.a(G516), .O(gate183inter7));
  inv1  gate1241(.a(G567), .O(gate183inter8));
  nand2 gate1242(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1243(.a(s_99), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1244(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1245(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1246(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1149(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1150(.a(gate184inter0), .b(s_86), .O(gate184inter1));
  and2  gate1151(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1152(.a(s_86), .O(gate184inter3));
  inv1  gate1153(.a(s_87), .O(gate184inter4));
  nand2 gate1154(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1155(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1156(.a(G519), .O(gate184inter7));
  inv1  gate1157(.a(G567), .O(gate184inter8));
  nand2 gate1158(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1159(.a(s_87), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1160(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1161(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1162(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1079(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1080(.a(gate185inter0), .b(s_76), .O(gate185inter1));
  and2  gate1081(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1082(.a(s_76), .O(gate185inter3));
  inv1  gate1083(.a(s_77), .O(gate185inter4));
  nand2 gate1084(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1085(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1086(.a(G570), .O(gate185inter7));
  inv1  gate1087(.a(G571), .O(gate185inter8));
  nand2 gate1088(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1089(.a(s_77), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1090(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1091(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1092(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate995(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate996(.a(gate188inter0), .b(s_64), .O(gate188inter1));
  and2  gate997(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate998(.a(s_64), .O(gate188inter3));
  inv1  gate999(.a(s_65), .O(gate188inter4));
  nand2 gate1000(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1001(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1002(.a(G576), .O(gate188inter7));
  inv1  gate1003(.a(G577), .O(gate188inter8));
  nand2 gate1004(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1005(.a(s_65), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1006(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1007(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1008(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1289(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1290(.a(gate195inter0), .b(s_106), .O(gate195inter1));
  and2  gate1291(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1292(.a(s_106), .O(gate195inter3));
  inv1  gate1293(.a(s_107), .O(gate195inter4));
  nand2 gate1294(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1295(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1296(.a(G590), .O(gate195inter7));
  inv1  gate1297(.a(G591), .O(gate195inter8));
  nand2 gate1298(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1299(.a(s_107), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1300(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1301(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1302(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate897(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate898(.a(gate208inter0), .b(s_50), .O(gate208inter1));
  and2  gate899(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate900(.a(s_50), .O(gate208inter3));
  inv1  gate901(.a(s_51), .O(gate208inter4));
  nand2 gate902(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate903(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate904(.a(G627), .O(gate208inter7));
  inv1  gate905(.a(G637), .O(gate208inter8));
  nand2 gate906(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate907(.a(s_51), .b(gate208inter3), .O(gate208inter10));
  nor2  gate908(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate909(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate910(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate729(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate730(.a(gate212inter0), .b(s_26), .O(gate212inter1));
  and2  gate731(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate732(.a(s_26), .O(gate212inter3));
  inv1  gate733(.a(s_27), .O(gate212inter4));
  nand2 gate734(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate735(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate736(.a(G617), .O(gate212inter7));
  inv1  gate737(.a(G669), .O(gate212inter8));
  nand2 gate738(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate739(.a(s_27), .b(gate212inter3), .O(gate212inter10));
  nor2  gate740(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate741(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate742(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate645(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate646(.a(gate221inter0), .b(s_14), .O(gate221inter1));
  and2  gate647(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate648(.a(s_14), .O(gate221inter3));
  inv1  gate649(.a(s_15), .O(gate221inter4));
  nand2 gate650(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate651(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate652(.a(G622), .O(gate221inter7));
  inv1  gate653(.a(G684), .O(gate221inter8));
  nand2 gate654(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate655(.a(s_15), .b(gate221inter3), .O(gate221inter10));
  nor2  gate656(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate657(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate658(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate869(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate870(.a(gate226inter0), .b(s_46), .O(gate226inter1));
  and2  gate871(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate872(.a(s_46), .O(gate226inter3));
  inv1  gate873(.a(s_47), .O(gate226inter4));
  nand2 gate874(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate875(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate876(.a(G692), .O(gate226inter7));
  inv1  gate877(.a(G693), .O(gate226inter8));
  nand2 gate878(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate879(.a(s_47), .b(gate226inter3), .O(gate226inter10));
  nor2  gate880(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate881(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate882(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate939(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate940(.a(gate227inter0), .b(s_56), .O(gate227inter1));
  and2  gate941(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate942(.a(s_56), .O(gate227inter3));
  inv1  gate943(.a(s_57), .O(gate227inter4));
  nand2 gate944(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate945(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate946(.a(G694), .O(gate227inter7));
  inv1  gate947(.a(G695), .O(gate227inter8));
  nand2 gate948(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate949(.a(s_57), .b(gate227inter3), .O(gate227inter10));
  nor2  gate950(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate951(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate952(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1303(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1304(.a(gate228inter0), .b(s_108), .O(gate228inter1));
  and2  gate1305(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1306(.a(s_108), .O(gate228inter3));
  inv1  gate1307(.a(s_109), .O(gate228inter4));
  nand2 gate1308(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1309(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1310(.a(G696), .O(gate228inter7));
  inv1  gate1311(.a(G697), .O(gate228inter8));
  nand2 gate1312(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1313(.a(s_109), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1314(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1315(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1316(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate967(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate968(.a(gate230inter0), .b(s_60), .O(gate230inter1));
  and2  gate969(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate970(.a(s_60), .O(gate230inter3));
  inv1  gate971(.a(s_61), .O(gate230inter4));
  nand2 gate972(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate973(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate974(.a(G700), .O(gate230inter7));
  inv1  gate975(.a(G701), .O(gate230inter8));
  nand2 gate976(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate977(.a(s_61), .b(gate230inter3), .O(gate230inter10));
  nor2  gate978(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate979(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate980(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate687(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate688(.a(gate231inter0), .b(s_20), .O(gate231inter1));
  and2  gate689(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate690(.a(s_20), .O(gate231inter3));
  inv1  gate691(.a(s_21), .O(gate231inter4));
  nand2 gate692(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate693(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate694(.a(G702), .O(gate231inter7));
  inv1  gate695(.a(G703), .O(gate231inter8));
  nand2 gate696(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate697(.a(s_21), .b(gate231inter3), .O(gate231inter10));
  nor2  gate698(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate699(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate700(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1373(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1374(.a(gate236inter0), .b(s_118), .O(gate236inter1));
  and2  gate1375(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1376(.a(s_118), .O(gate236inter3));
  inv1  gate1377(.a(s_119), .O(gate236inter4));
  nand2 gate1378(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1379(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1380(.a(G251), .O(gate236inter7));
  inv1  gate1381(.a(G727), .O(gate236inter8));
  nand2 gate1382(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1383(.a(s_119), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1384(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1385(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1386(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate827(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate828(.a(gate242inter0), .b(s_40), .O(gate242inter1));
  and2  gate829(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate830(.a(s_40), .O(gate242inter3));
  inv1  gate831(.a(s_41), .O(gate242inter4));
  nand2 gate832(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate833(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate834(.a(G718), .O(gate242inter7));
  inv1  gate835(.a(G730), .O(gate242inter8));
  nand2 gate836(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate837(.a(s_41), .b(gate242inter3), .O(gate242inter10));
  nor2  gate838(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate839(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate840(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate981(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate982(.a(gate248inter0), .b(s_62), .O(gate248inter1));
  and2  gate983(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate984(.a(s_62), .O(gate248inter3));
  inv1  gate985(.a(s_63), .O(gate248inter4));
  nand2 gate986(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate987(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate988(.a(G727), .O(gate248inter7));
  inv1  gate989(.a(G739), .O(gate248inter8));
  nand2 gate990(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate991(.a(s_63), .b(gate248inter3), .O(gate248inter10));
  nor2  gate992(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate993(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate994(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1135(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1136(.a(gate276inter0), .b(s_84), .O(gate276inter1));
  and2  gate1137(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1138(.a(s_84), .O(gate276inter3));
  inv1  gate1139(.a(s_85), .O(gate276inter4));
  nand2 gate1140(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1141(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1142(.a(G773), .O(gate276inter7));
  inv1  gate1143(.a(G797), .O(gate276inter8));
  nand2 gate1144(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1145(.a(s_85), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1146(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1147(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1148(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1107(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1108(.a(gate286inter0), .b(s_80), .O(gate286inter1));
  and2  gate1109(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1110(.a(s_80), .O(gate286inter3));
  inv1  gate1111(.a(s_81), .O(gate286inter4));
  nand2 gate1112(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1113(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1114(.a(G788), .O(gate286inter7));
  inv1  gate1115(.a(G812), .O(gate286inter8));
  nand2 gate1116(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1117(.a(s_81), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1118(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1119(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1120(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1247(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1248(.a(gate290inter0), .b(s_100), .O(gate290inter1));
  and2  gate1249(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1250(.a(s_100), .O(gate290inter3));
  inv1  gate1251(.a(s_101), .O(gate290inter4));
  nand2 gate1252(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1253(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1254(.a(G820), .O(gate290inter7));
  inv1  gate1255(.a(G821), .O(gate290inter8));
  nand2 gate1256(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1257(.a(s_101), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1258(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1259(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1260(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1219(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1220(.a(gate292inter0), .b(s_96), .O(gate292inter1));
  and2  gate1221(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1222(.a(s_96), .O(gate292inter3));
  inv1  gate1223(.a(s_97), .O(gate292inter4));
  nand2 gate1224(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1225(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1226(.a(G824), .O(gate292inter7));
  inv1  gate1227(.a(G825), .O(gate292inter8));
  nand2 gate1228(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1229(.a(s_97), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1230(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1231(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1232(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1317(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1318(.a(gate296inter0), .b(s_110), .O(gate296inter1));
  and2  gate1319(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1320(.a(s_110), .O(gate296inter3));
  inv1  gate1321(.a(s_111), .O(gate296inter4));
  nand2 gate1322(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1323(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1324(.a(G826), .O(gate296inter7));
  inv1  gate1325(.a(G827), .O(gate296inter8));
  nand2 gate1326(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1327(.a(s_111), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1328(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1329(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1330(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1261(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1262(.a(gate389inter0), .b(s_102), .O(gate389inter1));
  and2  gate1263(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1264(.a(s_102), .O(gate389inter3));
  inv1  gate1265(.a(s_103), .O(gate389inter4));
  nand2 gate1266(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1267(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1268(.a(G3), .O(gate389inter7));
  inv1  gate1269(.a(G1042), .O(gate389inter8));
  nand2 gate1270(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1271(.a(s_103), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1272(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1273(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1274(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate547(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate548(.a(gate392inter0), .b(s_0), .O(gate392inter1));
  and2  gate549(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate550(.a(s_0), .O(gate392inter3));
  inv1  gate551(.a(s_1), .O(gate392inter4));
  nand2 gate552(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate553(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate554(.a(G6), .O(gate392inter7));
  inv1  gate555(.a(G1051), .O(gate392inter8));
  nand2 gate556(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate557(.a(s_1), .b(gate392inter3), .O(gate392inter10));
  nor2  gate558(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate559(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate560(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1163(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1164(.a(gate394inter0), .b(s_88), .O(gate394inter1));
  and2  gate1165(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1166(.a(s_88), .O(gate394inter3));
  inv1  gate1167(.a(s_89), .O(gate394inter4));
  nand2 gate1168(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1169(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1170(.a(G8), .O(gate394inter7));
  inv1  gate1171(.a(G1057), .O(gate394inter8));
  nand2 gate1172(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1173(.a(s_89), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1174(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1175(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1176(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1345(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1346(.a(gate396inter0), .b(s_114), .O(gate396inter1));
  and2  gate1347(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1348(.a(s_114), .O(gate396inter3));
  inv1  gate1349(.a(s_115), .O(gate396inter4));
  nand2 gate1350(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1351(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1352(.a(G10), .O(gate396inter7));
  inv1  gate1353(.a(G1063), .O(gate396inter8));
  nand2 gate1354(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1355(.a(s_115), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1356(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1357(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1358(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1205(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1206(.a(gate398inter0), .b(s_94), .O(gate398inter1));
  and2  gate1207(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1208(.a(s_94), .O(gate398inter3));
  inv1  gate1209(.a(s_95), .O(gate398inter4));
  nand2 gate1210(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1211(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1212(.a(G12), .O(gate398inter7));
  inv1  gate1213(.a(G1069), .O(gate398inter8));
  nand2 gate1214(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1215(.a(s_95), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1216(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1217(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1218(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1457(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1458(.a(gate403inter0), .b(s_130), .O(gate403inter1));
  and2  gate1459(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1460(.a(s_130), .O(gate403inter3));
  inv1  gate1461(.a(s_131), .O(gate403inter4));
  nand2 gate1462(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1463(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1464(.a(G17), .O(gate403inter7));
  inv1  gate1465(.a(G1084), .O(gate403inter8));
  nand2 gate1466(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1467(.a(s_131), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1468(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1469(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1470(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1009(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1010(.a(gate414inter0), .b(s_66), .O(gate414inter1));
  and2  gate1011(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1012(.a(s_66), .O(gate414inter3));
  inv1  gate1013(.a(s_67), .O(gate414inter4));
  nand2 gate1014(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1015(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1016(.a(G28), .O(gate414inter7));
  inv1  gate1017(.a(G1117), .O(gate414inter8));
  nand2 gate1018(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1019(.a(s_67), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1020(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1021(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1022(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate603(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate604(.a(gate418inter0), .b(s_8), .O(gate418inter1));
  and2  gate605(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate606(.a(s_8), .O(gate418inter3));
  inv1  gate607(.a(s_9), .O(gate418inter4));
  nand2 gate608(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate609(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate610(.a(G32), .O(gate418inter7));
  inv1  gate611(.a(G1129), .O(gate418inter8));
  nand2 gate612(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate613(.a(s_9), .b(gate418inter3), .O(gate418inter10));
  nor2  gate614(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate615(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate616(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1065(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1066(.a(gate423inter0), .b(s_74), .O(gate423inter1));
  and2  gate1067(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1068(.a(s_74), .O(gate423inter3));
  inv1  gate1069(.a(s_75), .O(gate423inter4));
  nand2 gate1070(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1071(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1072(.a(G3), .O(gate423inter7));
  inv1  gate1073(.a(G1138), .O(gate423inter8));
  nand2 gate1074(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1075(.a(s_75), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1076(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1077(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1078(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate631(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate632(.a(gate425inter0), .b(s_12), .O(gate425inter1));
  and2  gate633(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate634(.a(s_12), .O(gate425inter3));
  inv1  gate635(.a(s_13), .O(gate425inter4));
  nand2 gate636(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate637(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate638(.a(G4), .O(gate425inter7));
  inv1  gate639(.a(G1141), .O(gate425inter8));
  nand2 gate640(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate641(.a(s_13), .b(gate425inter3), .O(gate425inter10));
  nor2  gate642(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate643(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate644(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate715(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate716(.a(gate432inter0), .b(s_24), .O(gate432inter1));
  and2  gate717(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate718(.a(s_24), .O(gate432inter3));
  inv1  gate719(.a(s_25), .O(gate432inter4));
  nand2 gate720(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate721(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate722(.a(G1054), .O(gate432inter7));
  inv1  gate723(.a(G1150), .O(gate432inter8));
  nand2 gate724(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate725(.a(s_25), .b(gate432inter3), .O(gate432inter10));
  nor2  gate726(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate727(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate728(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1443(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1444(.a(gate445inter0), .b(s_128), .O(gate445inter1));
  and2  gate1445(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1446(.a(s_128), .O(gate445inter3));
  inv1  gate1447(.a(s_129), .O(gate445inter4));
  nand2 gate1448(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1449(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1450(.a(G14), .O(gate445inter7));
  inv1  gate1451(.a(G1171), .O(gate445inter8));
  nand2 gate1452(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1453(.a(s_129), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1454(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1455(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1456(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate953(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate954(.a(gate449inter0), .b(s_58), .O(gate449inter1));
  and2  gate955(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate956(.a(s_58), .O(gate449inter3));
  inv1  gate957(.a(s_59), .O(gate449inter4));
  nand2 gate958(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate959(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate960(.a(G16), .O(gate449inter7));
  inv1  gate961(.a(G1177), .O(gate449inter8));
  nand2 gate962(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate963(.a(s_59), .b(gate449inter3), .O(gate449inter10));
  nor2  gate964(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate965(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate966(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate841(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate842(.a(gate452inter0), .b(s_42), .O(gate452inter1));
  and2  gate843(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate844(.a(s_42), .O(gate452inter3));
  inv1  gate845(.a(s_43), .O(gate452inter4));
  nand2 gate846(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate847(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate848(.a(G1084), .O(gate452inter7));
  inv1  gate849(.a(G1180), .O(gate452inter8));
  nand2 gate850(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate851(.a(s_43), .b(gate452inter3), .O(gate452inter10));
  nor2  gate852(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate853(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate854(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1415(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1416(.a(gate467inter0), .b(s_124), .O(gate467inter1));
  and2  gate1417(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1418(.a(s_124), .O(gate467inter3));
  inv1  gate1419(.a(s_125), .O(gate467inter4));
  nand2 gate1420(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1421(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1422(.a(G25), .O(gate467inter7));
  inv1  gate1423(.a(G1204), .O(gate467inter8));
  nand2 gate1424(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1425(.a(s_125), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1426(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1427(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1428(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate925(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate926(.a(gate471inter0), .b(s_54), .O(gate471inter1));
  and2  gate927(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate928(.a(s_54), .O(gate471inter3));
  inv1  gate929(.a(s_55), .O(gate471inter4));
  nand2 gate930(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate931(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate932(.a(G27), .O(gate471inter7));
  inv1  gate933(.a(G1210), .O(gate471inter8));
  nand2 gate934(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate935(.a(s_55), .b(gate471inter3), .O(gate471inter10));
  nor2  gate936(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate937(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate938(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate813(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate814(.a(gate480inter0), .b(s_38), .O(gate480inter1));
  and2  gate815(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate816(.a(s_38), .O(gate480inter3));
  inv1  gate817(.a(s_39), .O(gate480inter4));
  nand2 gate818(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate819(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate820(.a(G1126), .O(gate480inter7));
  inv1  gate821(.a(G1222), .O(gate480inter8));
  nand2 gate822(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate823(.a(s_39), .b(gate480inter3), .O(gate480inter10));
  nor2  gate824(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate825(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate826(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate617(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate618(.a(gate488inter0), .b(s_10), .O(gate488inter1));
  and2  gate619(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate620(.a(s_10), .O(gate488inter3));
  inv1  gate621(.a(s_11), .O(gate488inter4));
  nand2 gate622(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate623(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate624(.a(G1238), .O(gate488inter7));
  inv1  gate625(.a(G1239), .O(gate488inter8));
  nand2 gate626(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate627(.a(s_11), .b(gate488inter3), .O(gate488inter10));
  nor2  gate628(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate629(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate630(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1051(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1052(.a(gate492inter0), .b(s_72), .O(gate492inter1));
  and2  gate1053(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1054(.a(s_72), .O(gate492inter3));
  inv1  gate1055(.a(s_73), .O(gate492inter4));
  nand2 gate1056(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1057(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1058(.a(G1246), .O(gate492inter7));
  inv1  gate1059(.a(G1247), .O(gate492inter8));
  nand2 gate1060(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1061(.a(s_73), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1062(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1063(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1064(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1275(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1276(.a(gate507inter0), .b(s_104), .O(gate507inter1));
  and2  gate1277(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1278(.a(s_104), .O(gate507inter3));
  inv1  gate1279(.a(s_105), .O(gate507inter4));
  nand2 gate1280(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1281(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1282(.a(G1276), .O(gate507inter7));
  inv1  gate1283(.a(G1277), .O(gate507inter8));
  nand2 gate1284(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1285(.a(s_105), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1286(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1287(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1288(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1429(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1430(.a(gate509inter0), .b(s_126), .O(gate509inter1));
  and2  gate1431(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1432(.a(s_126), .O(gate509inter3));
  inv1  gate1433(.a(s_127), .O(gate509inter4));
  nand2 gate1434(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1435(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1436(.a(G1280), .O(gate509inter7));
  inv1  gate1437(.a(G1281), .O(gate509inter8));
  nand2 gate1438(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1439(.a(s_127), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1440(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1441(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1442(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule