module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1779(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1780(.a(gate10inter0), .b(s_176), .O(gate10inter1));
  and2  gate1781(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1782(.a(s_176), .O(gate10inter3));
  inv1  gate1783(.a(s_177), .O(gate10inter4));
  nand2 gate1784(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1785(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1786(.a(G3), .O(gate10inter7));
  inv1  gate1787(.a(G4), .O(gate10inter8));
  nand2 gate1788(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1789(.a(s_177), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1790(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1791(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1792(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate1849(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1850(.a(gate11inter0), .b(s_186), .O(gate11inter1));
  and2  gate1851(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1852(.a(s_186), .O(gate11inter3));
  inv1  gate1853(.a(s_187), .O(gate11inter4));
  nand2 gate1854(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1855(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1856(.a(G5), .O(gate11inter7));
  inv1  gate1857(.a(G6), .O(gate11inter8));
  nand2 gate1858(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1859(.a(s_187), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1860(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1861(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1862(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate631(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate632(.a(gate12inter0), .b(s_12), .O(gate12inter1));
  and2  gate633(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate634(.a(s_12), .O(gate12inter3));
  inv1  gate635(.a(s_13), .O(gate12inter4));
  nand2 gate636(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate637(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate638(.a(G7), .O(gate12inter7));
  inv1  gate639(.a(G8), .O(gate12inter8));
  nand2 gate640(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate641(.a(s_13), .b(gate12inter3), .O(gate12inter10));
  nor2  gate642(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate643(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate644(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate715(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate716(.a(gate15inter0), .b(s_24), .O(gate15inter1));
  and2  gate717(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate718(.a(s_24), .O(gate15inter3));
  inv1  gate719(.a(s_25), .O(gate15inter4));
  nand2 gate720(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate721(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate722(.a(G13), .O(gate15inter7));
  inv1  gate723(.a(G14), .O(gate15inter8));
  nand2 gate724(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate725(.a(s_25), .b(gate15inter3), .O(gate15inter10));
  nor2  gate726(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate727(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate728(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate645(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate646(.a(gate17inter0), .b(s_14), .O(gate17inter1));
  and2  gate647(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate648(.a(s_14), .O(gate17inter3));
  inv1  gate649(.a(s_15), .O(gate17inter4));
  nand2 gate650(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate651(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate652(.a(G17), .O(gate17inter7));
  inv1  gate653(.a(G18), .O(gate17inter8));
  nand2 gate654(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate655(.a(s_15), .b(gate17inter3), .O(gate17inter10));
  nor2  gate656(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate657(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate658(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1765(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1766(.a(gate24inter0), .b(s_174), .O(gate24inter1));
  and2  gate1767(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1768(.a(s_174), .O(gate24inter3));
  inv1  gate1769(.a(s_175), .O(gate24inter4));
  nand2 gate1770(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1771(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1772(.a(G31), .O(gate24inter7));
  inv1  gate1773(.a(G32), .O(gate24inter8));
  nand2 gate1774(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1775(.a(s_175), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1776(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1777(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1778(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate701(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate702(.a(gate32inter0), .b(s_22), .O(gate32inter1));
  and2  gate703(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate704(.a(s_22), .O(gate32inter3));
  inv1  gate705(.a(s_23), .O(gate32inter4));
  nand2 gate706(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate707(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate708(.a(G12), .O(gate32inter7));
  inv1  gate709(.a(G16), .O(gate32inter8));
  nand2 gate710(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate711(.a(s_23), .b(gate32inter3), .O(gate32inter10));
  nor2  gate712(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate713(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate714(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1429(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1430(.a(gate40inter0), .b(s_126), .O(gate40inter1));
  and2  gate1431(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1432(.a(s_126), .O(gate40inter3));
  inv1  gate1433(.a(s_127), .O(gate40inter4));
  nand2 gate1434(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1435(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1436(.a(G28), .O(gate40inter7));
  inv1  gate1437(.a(G32), .O(gate40inter8));
  nand2 gate1438(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1439(.a(s_127), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1440(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1441(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1442(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate995(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate996(.a(gate49inter0), .b(s_64), .O(gate49inter1));
  and2  gate997(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate998(.a(s_64), .O(gate49inter3));
  inv1  gate999(.a(s_65), .O(gate49inter4));
  nand2 gate1000(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1001(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1002(.a(G9), .O(gate49inter7));
  inv1  gate1003(.a(G278), .O(gate49inter8));
  nand2 gate1004(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1005(.a(s_65), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1006(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1007(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1008(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1471(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1472(.a(gate50inter0), .b(s_132), .O(gate50inter1));
  and2  gate1473(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1474(.a(s_132), .O(gate50inter3));
  inv1  gate1475(.a(s_133), .O(gate50inter4));
  nand2 gate1476(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1477(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1478(.a(G10), .O(gate50inter7));
  inv1  gate1479(.a(G278), .O(gate50inter8));
  nand2 gate1480(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1481(.a(s_133), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1482(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1483(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1484(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1933(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1934(.a(gate57inter0), .b(s_198), .O(gate57inter1));
  and2  gate1935(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1936(.a(s_198), .O(gate57inter3));
  inv1  gate1937(.a(s_199), .O(gate57inter4));
  nand2 gate1938(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1939(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1940(.a(G17), .O(gate57inter7));
  inv1  gate1941(.a(G290), .O(gate57inter8));
  nand2 gate1942(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1943(.a(s_199), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1944(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1945(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1946(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1947(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1948(.a(gate67inter0), .b(s_200), .O(gate67inter1));
  and2  gate1949(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1950(.a(s_200), .O(gate67inter3));
  inv1  gate1951(.a(s_201), .O(gate67inter4));
  nand2 gate1952(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1953(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1954(.a(G27), .O(gate67inter7));
  inv1  gate1955(.a(G305), .O(gate67inter8));
  nand2 gate1956(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1957(.a(s_201), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1958(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1959(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1960(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1205(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1206(.a(gate69inter0), .b(s_94), .O(gate69inter1));
  and2  gate1207(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1208(.a(s_94), .O(gate69inter3));
  inv1  gate1209(.a(s_95), .O(gate69inter4));
  nand2 gate1210(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1211(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1212(.a(G29), .O(gate69inter7));
  inv1  gate1213(.a(G308), .O(gate69inter8));
  nand2 gate1214(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1215(.a(s_95), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1216(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1217(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1218(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1751(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1752(.a(gate70inter0), .b(s_172), .O(gate70inter1));
  and2  gate1753(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1754(.a(s_172), .O(gate70inter3));
  inv1  gate1755(.a(s_173), .O(gate70inter4));
  nand2 gate1756(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1757(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1758(.a(G30), .O(gate70inter7));
  inv1  gate1759(.a(G308), .O(gate70inter8));
  nand2 gate1760(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1761(.a(s_173), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1762(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1763(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1764(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate743(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate744(.a(gate73inter0), .b(s_28), .O(gate73inter1));
  and2  gate745(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate746(.a(s_28), .O(gate73inter3));
  inv1  gate747(.a(s_29), .O(gate73inter4));
  nand2 gate748(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate749(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate750(.a(G1), .O(gate73inter7));
  inv1  gate751(.a(G314), .O(gate73inter8));
  nand2 gate752(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate753(.a(s_29), .b(gate73inter3), .O(gate73inter10));
  nor2  gate754(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate755(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate756(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1331(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1332(.a(gate76inter0), .b(s_112), .O(gate76inter1));
  and2  gate1333(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1334(.a(s_112), .O(gate76inter3));
  inv1  gate1335(.a(s_113), .O(gate76inter4));
  nand2 gate1336(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1337(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1338(.a(G13), .O(gate76inter7));
  inv1  gate1339(.a(G317), .O(gate76inter8));
  nand2 gate1340(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1341(.a(s_113), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1342(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1343(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1344(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate967(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate968(.a(gate78inter0), .b(s_60), .O(gate78inter1));
  and2  gate969(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate970(.a(s_60), .O(gate78inter3));
  inv1  gate971(.a(s_61), .O(gate78inter4));
  nand2 gate972(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate973(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate974(.a(G6), .O(gate78inter7));
  inv1  gate975(.a(G320), .O(gate78inter8));
  nand2 gate976(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate977(.a(s_61), .b(gate78inter3), .O(gate78inter10));
  nor2  gate978(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate979(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate980(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1345(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1346(.a(gate85inter0), .b(s_114), .O(gate85inter1));
  and2  gate1347(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1348(.a(s_114), .O(gate85inter3));
  inv1  gate1349(.a(s_115), .O(gate85inter4));
  nand2 gate1350(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1351(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1352(.a(G4), .O(gate85inter7));
  inv1  gate1353(.a(G332), .O(gate85inter8));
  nand2 gate1354(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1355(.a(s_115), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1356(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1357(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1358(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate603(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate604(.a(gate86inter0), .b(s_8), .O(gate86inter1));
  and2  gate605(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate606(.a(s_8), .O(gate86inter3));
  inv1  gate607(.a(s_9), .O(gate86inter4));
  nand2 gate608(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate609(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate610(.a(G8), .O(gate86inter7));
  inv1  gate611(.a(G332), .O(gate86inter8));
  nand2 gate612(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate613(.a(s_9), .b(gate86inter3), .O(gate86inter10));
  nor2  gate614(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate615(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate616(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate659(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate660(.a(gate87inter0), .b(s_16), .O(gate87inter1));
  and2  gate661(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate662(.a(s_16), .O(gate87inter3));
  inv1  gate663(.a(s_17), .O(gate87inter4));
  nand2 gate664(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate665(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate666(.a(G12), .O(gate87inter7));
  inv1  gate667(.a(G335), .O(gate87inter8));
  nand2 gate668(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate669(.a(s_17), .b(gate87inter3), .O(gate87inter10));
  nor2  gate670(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate671(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate672(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate953(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate954(.a(gate89inter0), .b(s_58), .O(gate89inter1));
  and2  gate955(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate956(.a(s_58), .O(gate89inter3));
  inv1  gate957(.a(s_59), .O(gate89inter4));
  nand2 gate958(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate959(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate960(.a(G17), .O(gate89inter7));
  inv1  gate961(.a(G338), .O(gate89inter8));
  nand2 gate962(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate963(.a(s_59), .b(gate89inter3), .O(gate89inter10));
  nor2  gate964(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate965(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate966(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1583(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1584(.a(gate94inter0), .b(s_148), .O(gate94inter1));
  and2  gate1585(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1586(.a(s_148), .O(gate94inter3));
  inv1  gate1587(.a(s_149), .O(gate94inter4));
  nand2 gate1588(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1589(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1590(.a(G22), .O(gate94inter7));
  inv1  gate1591(.a(G344), .O(gate94inter8));
  nand2 gate1592(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1593(.a(s_149), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1594(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1595(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1596(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate981(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate982(.a(gate98inter0), .b(s_62), .O(gate98inter1));
  and2  gate983(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate984(.a(s_62), .O(gate98inter3));
  inv1  gate985(.a(s_63), .O(gate98inter4));
  nand2 gate986(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate987(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate988(.a(G23), .O(gate98inter7));
  inv1  gate989(.a(G350), .O(gate98inter8));
  nand2 gate990(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate991(.a(s_63), .b(gate98inter3), .O(gate98inter10));
  nor2  gate992(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate993(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate994(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1877(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1878(.a(gate102inter0), .b(s_190), .O(gate102inter1));
  and2  gate1879(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1880(.a(s_190), .O(gate102inter3));
  inv1  gate1881(.a(s_191), .O(gate102inter4));
  nand2 gate1882(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1883(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1884(.a(G24), .O(gate102inter7));
  inv1  gate1885(.a(G356), .O(gate102inter8));
  nand2 gate1886(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1887(.a(s_191), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1888(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1889(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1890(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate897(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate898(.a(gate108inter0), .b(s_50), .O(gate108inter1));
  and2  gate899(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate900(.a(s_50), .O(gate108inter3));
  inv1  gate901(.a(s_51), .O(gate108inter4));
  nand2 gate902(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate903(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate904(.a(G368), .O(gate108inter7));
  inv1  gate905(.a(G369), .O(gate108inter8));
  nand2 gate906(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate907(.a(s_51), .b(gate108inter3), .O(gate108inter10));
  nor2  gate908(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate909(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate910(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1065(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1066(.a(gate109inter0), .b(s_74), .O(gate109inter1));
  and2  gate1067(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1068(.a(s_74), .O(gate109inter3));
  inv1  gate1069(.a(s_75), .O(gate109inter4));
  nand2 gate1070(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1071(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1072(.a(G370), .O(gate109inter7));
  inv1  gate1073(.a(G371), .O(gate109inter8));
  nand2 gate1074(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1075(.a(s_75), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1076(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1077(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1078(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1555(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1556(.a(gate110inter0), .b(s_144), .O(gate110inter1));
  and2  gate1557(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1558(.a(s_144), .O(gate110inter3));
  inv1  gate1559(.a(s_145), .O(gate110inter4));
  nand2 gate1560(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1561(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1562(.a(G372), .O(gate110inter7));
  inv1  gate1563(.a(G373), .O(gate110inter8));
  nand2 gate1564(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1565(.a(s_145), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1566(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1567(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1568(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate561(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate562(.a(gate114inter0), .b(s_2), .O(gate114inter1));
  and2  gate563(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate564(.a(s_2), .O(gate114inter3));
  inv1  gate565(.a(s_3), .O(gate114inter4));
  nand2 gate566(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate567(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate568(.a(G380), .O(gate114inter7));
  inv1  gate569(.a(G381), .O(gate114inter8));
  nand2 gate570(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate571(.a(s_3), .b(gate114inter3), .O(gate114inter10));
  nor2  gate572(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate573(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate574(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1639(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1640(.a(gate118inter0), .b(s_156), .O(gate118inter1));
  and2  gate1641(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1642(.a(s_156), .O(gate118inter3));
  inv1  gate1643(.a(s_157), .O(gate118inter4));
  nand2 gate1644(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1645(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1646(.a(G388), .O(gate118inter7));
  inv1  gate1647(.a(G389), .O(gate118inter8));
  nand2 gate1648(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1649(.a(s_157), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1650(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1651(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1652(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1793(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1794(.a(gate119inter0), .b(s_178), .O(gate119inter1));
  and2  gate1795(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1796(.a(s_178), .O(gate119inter3));
  inv1  gate1797(.a(s_179), .O(gate119inter4));
  nand2 gate1798(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1799(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1800(.a(G390), .O(gate119inter7));
  inv1  gate1801(.a(G391), .O(gate119inter8));
  nand2 gate1802(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1803(.a(s_179), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1804(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1805(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1806(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate589(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate590(.a(gate120inter0), .b(s_6), .O(gate120inter1));
  and2  gate591(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate592(.a(s_6), .O(gate120inter3));
  inv1  gate593(.a(s_7), .O(gate120inter4));
  nand2 gate594(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate595(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate596(.a(G392), .O(gate120inter7));
  inv1  gate597(.a(G393), .O(gate120inter8));
  nand2 gate598(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate599(.a(s_7), .b(gate120inter3), .O(gate120inter10));
  nor2  gate600(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate601(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate602(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate939(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate940(.a(gate121inter0), .b(s_56), .O(gate121inter1));
  and2  gate941(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate942(.a(s_56), .O(gate121inter3));
  inv1  gate943(.a(s_57), .O(gate121inter4));
  nand2 gate944(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate945(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate946(.a(G394), .O(gate121inter7));
  inv1  gate947(.a(G395), .O(gate121inter8));
  nand2 gate948(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate949(.a(s_57), .b(gate121inter3), .O(gate121inter10));
  nor2  gate950(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate951(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate952(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1219(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1220(.a(gate128inter0), .b(s_96), .O(gate128inter1));
  and2  gate1221(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1222(.a(s_96), .O(gate128inter3));
  inv1  gate1223(.a(s_97), .O(gate128inter4));
  nand2 gate1224(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1225(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1226(.a(G408), .O(gate128inter7));
  inv1  gate1227(.a(G409), .O(gate128inter8));
  nand2 gate1228(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1229(.a(s_97), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1230(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1231(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1232(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1569(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1570(.a(gate130inter0), .b(s_146), .O(gate130inter1));
  and2  gate1571(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1572(.a(s_146), .O(gate130inter3));
  inv1  gate1573(.a(s_147), .O(gate130inter4));
  nand2 gate1574(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1575(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1576(.a(G412), .O(gate130inter7));
  inv1  gate1577(.a(G413), .O(gate130inter8));
  nand2 gate1578(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1579(.a(s_147), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1580(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1581(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1582(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1737(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1738(.a(gate131inter0), .b(s_170), .O(gate131inter1));
  and2  gate1739(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1740(.a(s_170), .O(gate131inter3));
  inv1  gate1741(.a(s_171), .O(gate131inter4));
  nand2 gate1742(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1743(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1744(.a(G414), .O(gate131inter7));
  inv1  gate1745(.a(G415), .O(gate131inter8));
  nand2 gate1746(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1747(.a(s_171), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1748(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1749(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1750(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate855(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate856(.a(gate135inter0), .b(s_44), .O(gate135inter1));
  and2  gate857(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate858(.a(s_44), .O(gate135inter3));
  inv1  gate859(.a(s_45), .O(gate135inter4));
  nand2 gate860(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate861(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate862(.a(G422), .O(gate135inter7));
  inv1  gate863(.a(G423), .O(gate135inter8));
  nand2 gate864(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate865(.a(s_45), .b(gate135inter3), .O(gate135inter10));
  nor2  gate866(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate867(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate868(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1163(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1164(.a(gate137inter0), .b(s_88), .O(gate137inter1));
  and2  gate1165(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1166(.a(s_88), .O(gate137inter3));
  inv1  gate1167(.a(s_89), .O(gate137inter4));
  nand2 gate1168(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1169(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1170(.a(G426), .O(gate137inter7));
  inv1  gate1171(.a(G429), .O(gate137inter8));
  nand2 gate1172(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1173(.a(s_89), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1174(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1175(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1176(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1919(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1920(.a(gate145inter0), .b(s_196), .O(gate145inter1));
  and2  gate1921(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1922(.a(s_196), .O(gate145inter3));
  inv1  gate1923(.a(s_197), .O(gate145inter4));
  nand2 gate1924(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1925(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1926(.a(G474), .O(gate145inter7));
  inv1  gate1927(.a(G477), .O(gate145inter8));
  nand2 gate1928(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1929(.a(s_197), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1930(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1931(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1932(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1135(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1136(.a(gate150inter0), .b(s_84), .O(gate150inter1));
  and2  gate1137(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1138(.a(s_84), .O(gate150inter3));
  inv1  gate1139(.a(s_85), .O(gate150inter4));
  nand2 gate1140(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1141(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1142(.a(G504), .O(gate150inter7));
  inv1  gate1143(.a(G507), .O(gate150inter8));
  nand2 gate1144(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1145(.a(s_85), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1146(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1147(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1148(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate729(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate730(.a(gate159inter0), .b(s_26), .O(gate159inter1));
  and2  gate731(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate732(.a(s_26), .O(gate159inter3));
  inv1  gate733(.a(s_27), .O(gate159inter4));
  nand2 gate734(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate735(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate736(.a(G444), .O(gate159inter7));
  inv1  gate737(.a(G531), .O(gate159inter8));
  nand2 gate738(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate739(.a(s_27), .b(gate159inter3), .O(gate159inter10));
  nor2  gate740(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate741(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate742(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1233(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1234(.a(gate162inter0), .b(s_98), .O(gate162inter1));
  and2  gate1235(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1236(.a(s_98), .O(gate162inter3));
  inv1  gate1237(.a(s_99), .O(gate162inter4));
  nand2 gate1238(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1239(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1240(.a(G453), .O(gate162inter7));
  inv1  gate1241(.a(G534), .O(gate162inter8));
  nand2 gate1242(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1243(.a(s_99), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1244(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1245(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1246(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1415(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1416(.a(gate171inter0), .b(s_124), .O(gate171inter1));
  and2  gate1417(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1418(.a(s_124), .O(gate171inter3));
  inv1  gate1419(.a(s_125), .O(gate171inter4));
  nand2 gate1420(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1421(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1422(.a(G480), .O(gate171inter7));
  inv1  gate1423(.a(G549), .O(gate171inter8));
  nand2 gate1424(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1425(.a(s_125), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1426(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1427(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1428(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate575(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate576(.a(gate172inter0), .b(s_4), .O(gate172inter1));
  and2  gate577(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate578(.a(s_4), .O(gate172inter3));
  inv1  gate579(.a(s_5), .O(gate172inter4));
  nand2 gate580(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate581(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate582(.a(G483), .O(gate172inter7));
  inv1  gate583(.a(G549), .O(gate172inter8));
  nand2 gate584(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate585(.a(s_5), .b(gate172inter3), .O(gate172inter10));
  nor2  gate586(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate587(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate588(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1667(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1668(.a(gate192inter0), .b(s_160), .O(gate192inter1));
  and2  gate1669(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1670(.a(s_160), .O(gate192inter3));
  inv1  gate1671(.a(s_161), .O(gate192inter4));
  nand2 gate1672(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1673(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1674(.a(G584), .O(gate192inter7));
  inv1  gate1675(.a(G585), .O(gate192inter8));
  nand2 gate1676(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1677(.a(s_161), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1678(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1679(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1680(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1527(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1528(.a(gate201inter0), .b(s_140), .O(gate201inter1));
  and2  gate1529(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1530(.a(s_140), .O(gate201inter3));
  inv1  gate1531(.a(s_141), .O(gate201inter4));
  nand2 gate1532(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1533(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1534(.a(G602), .O(gate201inter7));
  inv1  gate1535(.a(G607), .O(gate201inter8));
  nand2 gate1536(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1537(.a(s_141), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1538(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1539(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1540(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1807(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1808(.a(gate203inter0), .b(s_180), .O(gate203inter1));
  and2  gate1809(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1810(.a(s_180), .O(gate203inter3));
  inv1  gate1811(.a(s_181), .O(gate203inter4));
  nand2 gate1812(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1813(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1814(.a(G602), .O(gate203inter7));
  inv1  gate1815(.a(G612), .O(gate203inter8));
  nand2 gate1816(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1817(.a(s_181), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1818(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1819(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1820(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1191(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1192(.a(gate205inter0), .b(s_92), .O(gate205inter1));
  and2  gate1193(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1194(.a(s_92), .O(gate205inter3));
  inv1  gate1195(.a(s_93), .O(gate205inter4));
  nand2 gate1196(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1197(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1198(.a(G622), .O(gate205inter7));
  inv1  gate1199(.a(G627), .O(gate205inter8));
  nand2 gate1200(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1201(.a(s_93), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1202(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1203(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1204(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1093(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1094(.a(gate214inter0), .b(s_78), .O(gate214inter1));
  and2  gate1095(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1096(.a(s_78), .O(gate214inter3));
  inv1  gate1097(.a(s_79), .O(gate214inter4));
  nand2 gate1098(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1099(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1100(.a(G612), .O(gate214inter7));
  inv1  gate1101(.a(G672), .O(gate214inter8));
  nand2 gate1102(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1103(.a(s_79), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1104(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1105(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1106(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate687(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate688(.a(gate217inter0), .b(s_20), .O(gate217inter1));
  and2  gate689(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate690(.a(s_20), .O(gate217inter3));
  inv1  gate691(.a(s_21), .O(gate217inter4));
  nand2 gate692(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate693(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate694(.a(G622), .O(gate217inter7));
  inv1  gate695(.a(G678), .O(gate217inter8));
  nand2 gate696(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate697(.a(s_21), .b(gate217inter3), .O(gate217inter10));
  nor2  gate698(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate699(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate700(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate911(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate912(.a(gate219inter0), .b(s_52), .O(gate219inter1));
  and2  gate913(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate914(.a(s_52), .O(gate219inter3));
  inv1  gate915(.a(s_53), .O(gate219inter4));
  nand2 gate916(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate917(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate918(.a(G632), .O(gate219inter7));
  inv1  gate919(.a(G681), .O(gate219inter8));
  nand2 gate920(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate921(.a(s_53), .b(gate219inter3), .O(gate219inter10));
  nor2  gate922(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate923(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate924(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1401(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1402(.a(gate221inter0), .b(s_122), .O(gate221inter1));
  and2  gate1403(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1404(.a(s_122), .O(gate221inter3));
  inv1  gate1405(.a(s_123), .O(gate221inter4));
  nand2 gate1406(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1407(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1408(.a(G622), .O(gate221inter7));
  inv1  gate1409(.a(G684), .O(gate221inter8));
  nand2 gate1410(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1411(.a(s_123), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1412(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1413(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1414(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1359(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1360(.a(gate222inter0), .b(s_116), .O(gate222inter1));
  and2  gate1361(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1362(.a(s_116), .O(gate222inter3));
  inv1  gate1363(.a(s_117), .O(gate222inter4));
  nand2 gate1364(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1365(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1366(.a(G632), .O(gate222inter7));
  inv1  gate1367(.a(G684), .O(gate222inter8));
  nand2 gate1368(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1369(.a(s_117), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1370(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1371(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1372(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1625(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1626(.a(gate230inter0), .b(s_154), .O(gate230inter1));
  and2  gate1627(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1628(.a(s_154), .O(gate230inter3));
  inv1  gate1629(.a(s_155), .O(gate230inter4));
  nand2 gate1630(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1631(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1632(.a(G700), .O(gate230inter7));
  inv1  gate1633(.a(G701), .O(gate230inter8));
  nand2 gate1634(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1635(.a(s_155), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1636(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1637(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1638(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1891(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1892(.a(gate234inter0), .b(s_192), .O(gate234inter1));
  and2  gate1893(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1894(.a(s_192), .O(gate234inter3));
  inv1  gate1895(.a(s_193), .O(gate234inter4));
  nand2 gate1896(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1897(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1898(.a(G245), .O(gate234inter7));
  inv1  gate1899(.a(G721), .O(gate234inter8));
  nand2 gate1900(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1901(.a(s_193), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1902(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1903(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1904(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate673(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate674(.a(gate244inter0), .b(s_18), .O(gate244inter1));
  and2  gate675(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate676(.a(s_18), .O(gate244inter3));
  inv1  gate677(.a(s_19), .O(gate244inter4));
  nand2 gate678(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate679(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate680(.a(G721), .O(gate244inter7));
  inv1  gate681(.a(G733), .O(gate244inter8));
  nand2 gate682(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate683(.a(s_19), .b(gate244inter3), .O(gate244inter10));
  nor2  gate684(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate685(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate686(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1317(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1318(.a(gate255inter0), .b(s_110), .O(gate255inter1));
  and2  gate1319(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1320(.a(s_110), .O(gate255inter3));
  inv1  gate1321(.a(s_111), .O(gate255inter4));
  nand2 gate1322(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1323(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1324(.a(G263), .O(gate255inter7));
  inv1  gate1325(.a(G751), .O(gate255inter8));
  nand2 gate1326(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1327(.a(s_111), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1328(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1329(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1330(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate925(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate926(.a(gate256inter0), .b(s_54), .O(gate256inter1));
  and2  gate927(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate928(.a(s_54), .O(gate256inter3));
  inv1  gate929(.a(s_55), .O(gate256inter4));
  nand2 gate930(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate931(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate932(.a(G715), .O(gate256inter7));
  inv1  gate933(.a(G751), .O(gate256inter8));
  nand2 gate934(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate935(.a(s_55), .b(gate256inter3), .O(gate256inter10));
  nor2  gate936(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate937(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate938(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1709(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1710(.a(gate258inter0), .b(s_166), .O(gate258inter1));
  and2  gate1711(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1712(.a(s_166), .O(gate258inter3));
  inv1  gate1713(.a(s_167), .O(gate258inter4));
  nand2 gate1714(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1715(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1716(.a(G756), .O(gate258inter7));
  inv1  gate1717(.a(G757), .O(gate258inter8));
  nand2 gate1718(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1719(.a(s_167), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1720(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1721(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1722(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1247(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1248(.a(gate264inter0), .b(s_100), .O(gate264inter1));
  and2  gate1249(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1250(.a(s_100), .O(gate264inter3));
  inv1  gate1251(.a(s_101), .O(gate264inter4));
  nand2 gate1252(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1253(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1254(.a(G768), .O(gate264inter7));
  inv1  gate1255(.a(G769), .O(gate264inter8));
  nand2 gate1256(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1257(.a(s_101), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1258(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1259(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1260(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1009(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1010(.a(gate265inter0), .b(s_66), .O(gate265inter1));
  and2  gate1011(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1012(.a(s_66), .O(gate265inter3));
  inv1  gate1013(.a(s_67), .O(gate265inter4));
  nand2 gate1014(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1015(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1016(.a(G642), .O(gate265inter7));
  inv1  gate1017(.a(G770), .O(gate265inter8));
  nand2 gate1018(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1019(.a(s_67), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1020(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1021(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1022(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1695(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1696(.a(gate267inter0), .b(s_164), .O(gate267inter1));
  and2  gate1697(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1698(.a(s_164), .O(gate267inter3));
  inv1  gate1699(.a(s_165), .O(gate267inter4));
  nand2 gate1700(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1701(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1702(.a(G648), .O(gate267inter7));
  inv1  gate1703(.a(G776), .O(gate267inter8));
  nand2 gate1704(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1705(.a(s_165), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1706(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1707(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1708(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1485(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1486(.a(gate269inter0), .b(s_134), .O(gate269inter1));
  and2  gate1487(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1488(.a(s_134), .O(gate269inter3));
  inv1  gate1489(.a(s_135), .O(gate269inter4));
  nand2 gate1490(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1491(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1492(.a(G654), .O(gate269inter7));
  inv1  gate1493(.a(G782), .O(gate269inter8));
  nand2 gate1494(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1495(.a(s_135), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1496(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1497(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1498(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1541(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1542(.a(gate273inter0), .b(s_142), .O(gate273inter1));
  and2  gate1543(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1544(.a(s_142), .O(gate273inter3));
  inv1  gate1545(.a(s_143), .O(gate273inter4));
  nand2 gate1546(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1547(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1548(.a(G642), .O(gate273inter7));
  inv1  gate1549(.a(G794), .O(gate273inter8));
  nand2 gate1550(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1551(.a(s_143), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1552(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1553(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1554(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1289(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1290(.a(gate277inter0), .b(s_106), .O(gate277inter1));
  and2  gate1291(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1292(.a(s_106), .O(gate277inter3));
  inv1  gate1293(.a(s_107), .O(gate277inter4));
  nand2 gate1294(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1295(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1296(.a(G648), .O(gate277inter7));
  inv1  gate1297(.a(G800), .O(gate277inter8));
  nand2 gate1298(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1299(.a(s_107), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1300(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1301(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1302(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1037(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1038(.a(gate282inter0), .b(s_70), .O(gate282inter1));
  and2  gate1039(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1040(.a(s_70), .O(gate282inter3));
  inv1  gate1041(.a(s_71), .O(gate282inter4));
  nand2 gate1042(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1043(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1044(.a(G782), .O(gate282inter7));
  inv1  gate1045(.a(G806), .O(gate282inter8));
  nand2 gate1046(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1047(.a(s_71), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1048(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1049(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1050(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1387(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1388(.a(gate286inter0), .b(s_120), .O(gate286inter1));
  and2  gate1389(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1390(.a(s_120), .O(gate286inter3));
  inv1  gate1391(.a(s_121), .O(gate286inter4));
  nand2 gate1392(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1393(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1394(.a(G788), .O(gate286inter7));
  inv1  gate1395(.a(G812), .O(gate286inter8));
  nand2 gate1396(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1397(.a(s_121), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1398(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1399(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1400(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1653(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1654(.a(gate290inter0), .b(s_158), .O(gate290inter1));
  and2  gate1655(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1656(.a(s_158), .O(gate290inter3));
  inv1  gate1657(.a(s_159), .O(gate290inter4));
  nand2 gate1658(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1659(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1660(.a(G820), .O(gate290inter7));
  inv1  gate1661(.a(G821), .O(gate290inter8));
  nand2 gate1662(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1663(.a(s_159), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1664(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1665(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1666(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1611(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1612(.a(gate291inter0), .b(s_152), .O(gate291inter1));
  and2  gate1613(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1614(.a(s_152), .O(gate291inter3));
  inv1  gate1615(.a(s_153), .O(gate291inter4));
  nand2 gate1616(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1617(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1618(.a(G822), .O(gate291inter7));
  inv1  gate1619(.a(G823), .O(gate291inter8));
  nand2 gate1620(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1621(.a(s_153), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1622(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1623(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1624(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1863(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1864(.a(gate293inter0), .b(s_188), .O(gate293inter1));
  and2  gate1865(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1866(.a(s_188), .O(gate293inter3));
  inv1  gate1867(.a(s_189), .O(gate293inter4));
  nand2 gate1868(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1869(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1870(.a(G828), .O(gate293inter7));
  inv1  gate1871(.a(G829), .O(gate293inter8));
  nand2 gate1872(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1873(.a(s_189), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1874(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1875(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1876(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1275(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1276(.a(gate387inter0), .b(s_104), .O(gate387inter1));
  and2  gate1277(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1278(.a(s_104), .O(gate387inter3));
  inv1  gate1279(.a(s_105), .O(gate387inter4));
  nand2 gate1280(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1281(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1282(.a(G1), .O(gate387inter7));
  inv1  gate1283(.a(G1036), .O(gate387inter8));
  nand2 gate1284(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1285(.a(s_105), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1286(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1287(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1288(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1905(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1906(.a(gate389inter0), .b(s_194), .O(gate389inter1));
  and2  gate1907(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1908(.a(s_194), .O(gate389inter3));
  inv1  gate1909(.a(s_195), .O(gate389inter4));
  nand2 gate1910(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1911(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1912(.a(G3), .O(gate389inter7));
  inv1  gate1913(.a(G1042), .O(gate389inter8));
  nand2 gate1914(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1915(.a(s_195), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1916(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1917(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1918(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate617(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate618(.a(gate391inter0), .b(s_10), .O(gate391inter1));
  and2  gate619(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate620(.a(s_10), .O(gate391inter3));
  inv1  gate621(.a(s_11), .O(gate391inter4));
  nand2 gate622(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate623(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate624(.a(G5), .O(gate391inter7));
  inv1  gate625(.a(G1048), .O(gate391inter8));
  nand2 gate626(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate627(.a(s_11), .b(gate391inter3), .O(gate391inter10));
  nor2  gate628(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate629(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate630(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1107(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1108(.a(gate396inter0), .b(s_80), .O(gate396inter1));
  and2  gate1109(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1110(.a(s_80), .O(gate396inter3));
  inv1  gate1111(.a(s_81), .O(gate396inter4));
  nand2 gate1112(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1113(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1114(.a(G10), .O(gate396inter7));
  inv1  gate1115(.a(G1063), .O(gate396inter8));
  nand2 gate1116(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1117(.a(s_81), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1118(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1119(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1120(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1443(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1444(.a(gate399inter0), .b(s_128), .O(gate399inter1));
  and2  gate1445(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1446(.a(s_128), .O(gate399inter3));
  inv1  gate1447(.a(s_129), .O(gate399inter4));
  nand2 gate1448(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1449(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1450(.a(G13), .O(gate399inter7));
  inv1  gate1451(.a(G1072), .O(gate399inter8));
  nand2 gate1452(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1453(.a(s_129), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1454(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1455(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1456(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1835(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1836(.a(gate400inter0), .b(s_184), .O(gate400inter1));
  and2  gate1837(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1838(.a(s_184), .O(gate400inter3));
  inv1  gate1839(.a(s_185), .O(gate400inter4));
  nand2 gate1840(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1841(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1842(.a(G14), .O(gate400inter7));
  inv1  gate1843(.a(G1075), .O(gate400inter8));
  nand2 gate1844(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1845(.a(s_185), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1846(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1847(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1848(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate827(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate828(.a(gate411inter0), .b(s_40), .O(gate411inter1));
  and2  gate829(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate830(.a(s_40), .O(gate411inter3));
  inv1  gate831(.a(s_41), .O(gate411inter4));
  nand2 gate832(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate833(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate834(.a(G25), .O(gate411inter7));
  inv1  gate835(.a(G1108), .O(gate411inter8));
  nand2 gate836(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate837(.a(s_41), .b(gate411inter3), .O(gate411inter10));
  nor2  gate838(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate839(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate840(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1499(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1500(.a(gate420inter0), .b(s_136), .O(gate420inter1));
  and2  gate1501(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1502(.a(s_136), .O(gate420inter3));
  inv1  gate1503(.a(s_137), .O(gate420inter4));
  nand2 gate1504(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1505(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1506(.a(G1036), .O(gate420inter7));
  inv1  gate1507(.a(G1132), .O(gate420inter8));
  nand2 gate1508(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1509(.a(s_137), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1510(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1511(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1512(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate813(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate814(.a(gate421inter0), .b(s_38), .O(gate421inter1));
  and2  gate815(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate816(.a(s_38), .O(gate421inter3));
  inv1  gate817(.a(s_39), .O(gate421inter4));
  nand2 gate818(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate819(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate820(.a(G2), .O(gate421inter7));
  inv1  gate821(.a(G1135), .O(gate421inter8));
  nand2 gate822(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate823(.a(s_39), .b(gate421inter3), .O(gate421inter10));
  nor2  gate824(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate825(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate826(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1261(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1262(.a(gate425inter0), .b(s_102), .O(gate425inter1));
  and2  gate1263(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1264(.a(s_102), .O(gate425inter3));
  inv1  gate1265(.a(s_103), .O(gate425inter4));
  nand2 gate1266(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1267(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1268(.a(G4), .O(gate425inter7));
  inv1  gate1269(.a(G1141), .O(gate425inter8));
  nand2 gate1270(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1271(.a(s_103), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1272(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1273(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1274(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate771(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate772(.a(gate433inter0), .b(s_32), .O(gate433inter1));
  and2  gate773(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate774(.a(s_32), .O(gate433inter3));
  inv1  gate775(.a(s_33), .O(gate433inter4));
  nand2 gate776(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate777(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate778(.a(G8), .O(gate433inter7));
  inv1  gate779(.a(G1153), .O(gate433inter8));
  nand2 gate780(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate781(.a(s_33), .b(gate433inter3), .O(gate433inter10));
  nor2  gate782(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate783(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate784(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1051(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1052(.a(gate435inter0), .b(s_72), .O(gate435inter1));
  and2  gate1053(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1054(.a(s_72), .O(gate435inter3));
  inv1  gate1055(.a(s_73), .O(gate435inter4));
  nand2 gate1056(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1057(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1058(.a(G9), .O(gate435inter7));
  inv1  gate1059(.a(G1156), .O(gate435inter8));
  nand2 gate1060(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1061(.a(s_73), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1062(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1063(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1064(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate841(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate842(.a(gate448inter0), .b(s_42), .O(gate448inter1));
  and2  gate843(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate844(.a(s_42), .O(gate448inter3));
  inv1  gate845(.a(s_43), .O(gate448inter4));
  nand2 gate846(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate847(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate848(.a(G1078), .O(gate448inter7));
  inv1  gate849(.a(G1174), .O(gate448inter8));
  nand2 gate850(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate851(.a(s_43), .b(gate448inter3), .O(gate448inter10));
  nor2  gate852(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate853(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate854(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1121(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1122(.a(gate450inter0), .b(s_82), .O(gate450inter1));
  and2  gate1123(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1124(.a(s_82), .O(gate450inter3));
  inv1  gate1125(.a(s_83), .O(gate450inter4));
  nand2 gate1126(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1127(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1128(.a(G1081), .O(gate450inter7));
  inv1  gate1129(.a(G1177), .O(gate450inter8));
  nand2 gate1130(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1131(.a(s_83), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1132(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1133(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1134(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1023(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1024(.a(gate451inter0), .b(s_68), .O(gate451inter1));
  and2  gate1025(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1026(.a(s_68), .O(gate451inter3));
  inv1  gate1027(.a(s_69), .O(gate451inter4));
  nand2 gate1028(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1029(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1030(.a(G17), .O(gate451inter7));
  inv1  gate1031(.a(G1180), .O(gate451inter8));
  nand2 gate1032(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1033(.a(s_69), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1034(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1035(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1036(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1723(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1724(.a(gate453inter0), .b(s_168), .O(gate453inter1));
  and2  gate1725(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1726(.a(s_168), .O(gate453inter3));
  inv1  gate1727(.a(s_169), .O(gate453inter4));
  nand2 gate1728(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1729(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1730(.a(G18), .O(gate453inter7));
  inv1  gate1731(.a(G1183), .O(gate453inter8));
  nand2 gate1732(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1733(.a(s_169), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1734(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1735(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1736(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate883(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate884(.a(gate461inter0), .b(s_48), .O(gate461inter1));
  and2  gate885(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate886(.a(s_48), .O(gate461inter3));
  inv1  gate887(.a(s_49), .O(gate461inter4));
  nand2 gate888(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate889(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate890(.a(G22), .O(gate461inter7));
  inv1  gate891(.a(G1195), .O(gate461inter8));
  nand2 gate892(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate893(.a(s_49), .b(gate461inter3), .O(gate461inter10));
  nor2  gate894(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate895(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate896(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate547(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate548(.a(gate468inter0), .b(s_0), .O(gate468inter1));
  and2  gate549(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate550(.a(s_0), .O(gate468inter3));
  inv1  gate551(.a(s_1), .O(gate468inter4));
  nand2 gate552(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate553(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate554(.a(G1108), .O(gate468inter7));
  inv1  gate555(.a(G1204), .O(gate468inter8));
  nand2 gate556(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate557(.a(s_1), .b(gate468inter3), .O(gate468inter10));
  nor2  gate558(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate559(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate560(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1597(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1598(.a(gate477inter0), .b(s_150), .O(gate477inter1));
  and2  gate1599(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1600(.a(s_150), .O(gate477inter3));
  inv1  gate1601(.a(s_151), .O(gate477inter4));
  nand2 gate1602(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1603(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1604(.a(G30), .O(gate477inter7));
  inv1  gate1605(.a(G1219), .O(gate477inter8));
  nand2 gate1606(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1607(.a(s_151), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1608(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1609(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1610(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate785(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate786(.a(gate478inter0), .b(s_34), .O(gate478inter1));
  and2  gate787(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate788(.a(s_34), .O(gate478inter3));
  inv1  gate789(.a(s_35), .O(gate478inter4));
  nand2 gate790(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate791(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate792(.a(G1123), .O(gate478inter7));
  inv1  gate793(.a(G1219), .O(gate478inter8));
  nand2 gate794(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate795(.a(s_35), .b(gate478inter3), .O(gate478inter10));
  nor2  gate796(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate797(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate798(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1681(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1682(.a(gate486inter0), .b(s_162), .O(gate486inter1));
  and2  gate1683(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1684(.a(s_162), .O(gate486inter3));
  inv1  gate1685(.a(s_163), .O(gate486inter4));
  nand2 gate1686(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1687(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1688(.a(G1234), .O(gate486inter7));
  inv1  gate1689(.a(G1235), .O(gate486inter8));
  nand2 gate1690(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1691(.a(s_163), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1692(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1693(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1694(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1149(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1150(.a(gate489inter0), .b(s_86), .O(gate489inter1));
  and2  gate1151(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1152(.a(s_86), .O(gate489inter3));
  inv1  gate1153(.a(s_87), .O(gate489inter4));
  nand2 gate1154(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1155(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1156(.a(G1240), .O(gate489inter7));
  inv1  gate1157(.a(G1241), .O(gate489inter8));
  nand2 gate1158(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1159(.a(s_87), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1160(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1161(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1162(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1303(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1304(.a(gate493inter0), .b(s_108), .O(gate493inter1));
  and2  gate1305(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1306(.a(s_108), .O(gate493inter3));
  inv1  gate1307(.a(s_109), .O(gate493inter4));
  nand2 gate1308(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1309(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1310(.a(G1248), .O(gate493inter7));
  inv1  gate1311(.a(G1249), .O(gate493inter8));
  nand2 gate1312(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1313(.a(s_109), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1314(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1315(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1316(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1177(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1178(.a(gate494inter0), .b(s_90), .O(gate494inter1));
  and2  gate1179(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1180(.a(s_90), .O(gate494inter3));
  inv1  gate1181(.a(s_91), .O(gate494inter4));
  nand2 gate1182(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1183(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1184(.a(G1250), .O(gate494inter7));
  inv1  gate1185(.a(G1251), .O(gate494inter8));
  nand2 gate1186(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1187(.a(s_91), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1188(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1189(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1190(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate869(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate870(.a(gate497inter0), .b(s_46), .O(gate497inter1));
  and2  gate871(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate872(.a(s_46), .O(gate497inter3));
  inv1  gate873(.a(s_47), .O(gate497inter4));
  nand2 gate874(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate875(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate876(.a(G1256), .O(gate497inter7));
  inv1  gate877(.a(G1257), .O(gate497inter8));
  nand2 gate878(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate879(.a(s_47), .b(gate497inter3), .O(gate497inter10));
  nor2  gate880(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate881(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate882(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1821(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1822(.a(gate498inter0), .b(s_182), .O(gate498inter1));
  and2  gate1823(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1824(.a(s_182), .O(gate498inter3));
  inv1  gate1825(.a(s_183), .O(gate498inter4));
  nand2 gate1826(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1827(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1828(.a(G1258), .O(gate498inter7));
  inv1  gate1829(.a(G1259), .O(gate498inter8));
  nand2 gate1830(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1831(.a(s_183), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1832(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1833(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1834(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate799(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate800(.a(gate500inter0), .b(s_36), .O(gate500inter1));
  and2  gate801(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate802(.a(s_36), .O(gate500inter3));
  inv1  gate803(.a(s_37), .O(gate500inter4));
  nand2 gate804(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate805(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate806(.a(G1262), .O(gate500inter7));
  inv1  gate807(.a(G1263), .O(gate500inter8));
  nand2 gate808(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate809(.a(s_37), .b(gate500inter3), .O(gate500inter10));
  nor2  gate810(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate811(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate812(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate757(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate758(.a(gate504inter0), .b(s_30), .O(gate504inter1));
  and2  gate759(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate760(.a(s_30), .O(gate504inter3));
  inv1  gate761(.a(s_31), .O(gate504inter4));
  nand2 gate762(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate763(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate764(.a(G1270), .O(gate504inter7));
  inv1  gate765(.a(G1271), .O(gate504inter8));
  nand2 gate766(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate767(.a(s_31), .b(gate504inter3), .O(gate504inter10));
  nor2  gate768(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate769(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate770(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1373(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1374(.a(gate505inter0), .b(s_118), .O(gate505inter1));
  and2  gate1375(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1376(.a(s_118), .O(gate505inter3));
  inv1  gate1377(.a(s_119), .O(gate505inter4));
  nand2 gate1378(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1379(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1380(.a(G1272), .O(gate505inter7));
  inv1  gate1381(.a(G1273), .O(gate505inter8));
  nand2 gate1382(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1383(.a(s_119), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1384(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1385(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1386(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1079(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1080(.a(gate511inter0), .b(s_76), .O(gate511inter1));
  and2  gate1081(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1082(.a(s_76), .O(gate511inter3));
  inv1  gate1083(.a(s_77), .O(gate511inter4));
  nand2 gate1084(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1085(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1086(.a(G1284), .O(gate511inter7));
  inv1  gate1087(.a(G1285), .O(gate511inter8));
  nand2 gate1088(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1089(.a(s_77), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1090(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1091(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1092(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1457(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1458(.a(gate512inter0), .b(s_130), .O(gate512inter1));
  and2  gate1459(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1460(.a(s_130), .O(gate512inter3));
  inv1  gate1461(.a(s_131), .O(gate512inter4));
  nand2 gate1462(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1463(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1464(.a(G1286), .O(gate512inter7));
  inv1  gate1465(.a(G1287), .O(gate512inter8));
  nand2 gate1466(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1467(.a(s_131), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1468(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1469(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1470(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1513(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1514(.a(gate513inter0), .b(s_138), .O(gate513inter1));
  and2  gate1515(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1516(.a(s_138), .O(gate513inter3));
  inv1  gate1517(.a(s_139), .O(gate513inter4));
  nand2 gate1518(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1519(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1520(.a(G1288), .O(gate513inter7));
  inv1  gate1521(.a(G1289), .O(gate513inter8));
  nand2 gate1522(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1523(.a(s_139), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1524(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1525(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1526(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule