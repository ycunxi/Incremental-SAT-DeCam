module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate7inter0, gate7inter1, gate7inter2, gate7inter3, gate7inter4, gate7inter5, gate7inter6, gate7inter7, gate7inter8, gate7inter9, gate7inter10, gate7inter11, gate7inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate357(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate358(.a(gate4inter0), .b(s_22), .O(gate4inter1));
  and2  gate359(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate360(.a(s_22), .O(gate4inter3));
  inv1  gate361(.a(s_23), .O(gate4inter4));
  nand2 gate362(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate363(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate364(.a(N25), .O(gate4inter7));
  inv1  gate365(.a(N29), .O(gate4inter8));
  nand2 gate366(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate367(.a(s_23), .b(gate4inter3), .O(gate4inter10));
  nor2  gate368(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate369(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate370(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );

  xor2  gate273(.a(N53), .b(N49), .O(gate7inter0));
  nand2 gate274(.a(gate7inter0), .b(s_10), .O(gate7inter1));
  and2  gate275(.a(N53), .b(N49), .O(gate7inter2));
  inv1  gate276(.a(s_10), .O(gate7inter3));
  inv1  gate277(.a(s_11), .O(gate7inter4));
  nand2 gate278(.a(gate7inter4), .b(gate7inter3), .O(gate7inter5));
  nor2  gate279(.a(gate7inter5), .b(gate7inter2), .O(gate7inter6));
  inv1  gate280(.a(N49), .O(gate7inter7));
  inv1  gate281(.a(N53), .O(gate7inter8));
  nand2 gate282(.a(gate7inter8), .b(gate7inter7), .O(gate7inter9));
  nand2 gate283(.a(s_11), .b(gate7inter3), .O(gate7inter10));
  nor2  gate284(.a(gate7inter10), .b(gate7inter9), .O(gate7inter11));
  nor2  gate285(.a(gate7inter11), .b(gate7inter6), .O(gate7inter12));
  nand2 gate286(.a(gate7inter12), .b(gate7inter1), .O(N256));

  xor2  gate371(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate372(.a(gate8inter0), .b(s_24), .O(gate8inter1));
  and2  gate373(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate374(.a(s_24), .O(gate8inter3));
  inv1  gate375(.a(s_25), .O(gate8inter4));
  nand2 gate376(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate377(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate378(.a(N57), .O(gate8inter7));
  inv1  gate379(.a(N61), .O(gate8inter8));
  nand2 gate380(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate381(.a(s_25), .b(gate8inter3), .O(gate8inter10));
  nor2  gate382(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate383(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate384(.a(gate8inter12), .b(gate8inter1), .O(N257));
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );

  xor2  gate301(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate302(.a(gate13inter0), .b(s_14), .O(gate13inter1));
  and2  gate303(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate304(.a(s_14), .O(gate13inter3));
  inv1  gate305(.a(s_15), .O(gate13inter4));
  nand2 gate306(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate307(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate308(.a(N97), .O(gate13inter7));
  inv1  gate309(.a(N101), .O(gate13inter8));
  nand2 gate310(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate311(.a(s_15), .b(gate13inter3), .O(gate13inter10));
  nor2  gate312(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate313(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate314(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate203(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate204(.a(gate25inter0), .b(s_0), .O(gate25inter1));
  and2  gate205(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate206(.a(s_0), .O(gate25inter3));
  inv1  gate207(.a(s_1), .O(gate25inter4));
  nand2 gate208(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate209(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate210(.a(N1), .O(gate25inter7));
  inv1  gate211(.a(N17), .O(gate25inter8));
  nand2 gate212(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate213(.a(s_1), .b(gate25inter3), .O(gate25inter10));
  nor2  gate214(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate215(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate216(.a(gate25inter12), .b(gate25inter1), .O(N274));
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );

  xor2  gate245(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate246(.a(gate28inter0), .b(s_6), .O(gate28inter1));
  and2  gate247(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate248(.a(s_6), .O(gate28inter3));
  inv1  gate249(.a(s_7), .O(gate28inter4));
  nand2 gate250(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate251(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate252(.a(N37), .O(gate28inter7));
  inv1  gate253(.a(N53), .O(gate28inter8));
  nand2 gate254(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate255(.a(s_7), .b(gate28inter3), .O(gate28inter10));
  nor2  gate256(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate257(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate258(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );

  xor2  gate231(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate232(.a(gate31inter0), .b(s_4), .O(gate31inter1));
  and2  gate233(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate234(.a(s_4), .O(gate31inter3));
  inv1  gate235(.a(s_5), .O(gate31inter4));
  nand2 gate236(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate237(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate238(.a(N13), .O(gate31inter7));
  inv1  gate239(.a(N29), .O(gate31inter8));
  nand2 gate240(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate241(.a(s_5), .b(gate31inter3), .O(gate31inter10));
  nor2  gate242(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate243(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate244(.a(gate31inter12), .b(gate31inter1), .O(N280));
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );

  xor2  gate427(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate428(.a(gate43inter0), .b(s_32), .O(gate43inter1));
  and2  gate429(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate430(.a(s_32), .O(gate43inter3));
  inv1  gate431(.a(s_33), .O(gate43inter4));
  nand2 gate432(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate433(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate434(.a(N254), .O(gate43inter7));
  inv1  gate435(.a(N255), .O(gate43inter8));
  nand2 gate436(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate437(.a(s_33), .b(gate43inter3), .O(gate43inter10));
  nor2  gate438(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate439(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate440(.a(gate43inter12), .b(gate43inter1), .O(N296));
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );

  xor2  gate483(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate484(.a(gate48inter0), .b(s_40), .O(gate48inter1));
  and2  gate485(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate486(.a(s_40), .O(gate48inter3));
  inv1  gate487(.a(s_41), .O(gate48inter4));
  nand2 gate488(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate489(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate490(.a(N264), .O(gate48inter7));
  inv1  gate491(.a(N265), .O(gate48inter8));
  nand2 gate492(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate493(.a(s_41), .b(gate48inter3), .O(gate48inter10));
  nor2  gate494(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate495(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate496(.a(gate48inter12), .b(gate48inter1), .O(N311));

  xor2  gate259(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate260(.a(gate49inter0), .b(s_8), .O(gate49inter1));
  and2  gate261(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate262(.a(s_8), .O(gate49inter3));
  inv1  gate263(.a(s_9), .O(gate49inter4));
  nand2 gate264(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate265(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate266(.a(N274), .O(gate49inter7));
  inv1  gate267(.a(N275), .O(gate49inter8));
  nand2 gate268(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate269(.a(s_9), .b(gate49inter3), .O(gate49inter10));
  nor2  gate270(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate271(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate272(.a(gate49inter12), .b(gate49inter1), .O(N314));
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );

  xor2  gate287(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate288(.a(gate57inter0), .b(s_12), .O(gate57inter1));
  and2  gate289(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate290(.a(s_12), .O(gate57inter3));
  inv1  gate291(.a(s_13), .O(gate57inter4));
  nand2 gate292(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate293(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate294(.a(N290), .O(gate57inter7));
  inv1  gate295(.a(N293), .O(gate57inter8));
  nand2 gate296(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate297(.a(s_13), .b(gate57inter3), .O(gate57inter10));
  nor2  gate298(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate299(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate300(.a(gate57inter12), .b(gate57inter1), .O(N338));
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate413(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate414(.a(gate75inter0), .b(s_30), .O(gate75inter1));
  and2  gate415(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate416(.a(s_30), .O(gate75inter3));
  inv1  gate417(.a(s_31), .O(gate75inter4));
  nand2 gate418(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate419(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate420(.a(N316), .O(gate75inter7));
  inv1  gate421(.a(N348), .O(gate75inter8));
  nand2 gate422(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate423(.a(s_31), .b(gate75inter3), .O(gate75inter10));
  nor2  gate424(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate425(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate426(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate385(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate386(.a(gate172inter0), .b(s_26), .O(gate172inter1));
  and2  gate387(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate388(.a(s_26), .O(gate172inter3));
  inv1  gate389(.a(s_27), .O(gate172inter4));
  nand2 gate390(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate391(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate392(.a(N5), .O(gate172inter7));
  inv1  gate393(.a(N693), .O(gate172inter8));
  nand2 gate394(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate395(.a(s_27), .b(gate172inter3), .O(gate172inter10));
  nor2  gate396(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate397(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate398(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate343(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate344(.a(gate176inter0), .b(s_20), .O(gate176inter1));
  and2  gate345(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate346(.a(s_20), .O(gate176inter3));
  inv1  gate347(.a(s_21), .O(gate176inter4));
  nand2 gate348(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate349(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate350(.a(N21), .O(gate176inter7));
  inv1  gate351(.a(N697), .O(gate176inter8));
  nand2 gate352(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate353(.a(s_21), .b(gate176inter3), .O(gate176inter10));
  nor2  gate354(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate355(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate356(.a(gate176inter12), .b(gate176inter1), .O(N729));

  xor2  gate315(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate316(.a(gate177inter0), .b(s_16), .O(gate177inter1));
  and2  gate317(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate318(.a(s_16), .O(gate177inter3));
  inv1  gate319(.a(s_17), .O(gate177inter4));
  nand2 gate320(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate321(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate322(.a(N25), .O(gate177inter7));
  inv1  gate323(.a(N698), .O(gate177inter8));
  nand2 gate324(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate325(.a(s_17), .b(gate177inter3), .O(gate177inter10));
  nor2  gate326(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate327(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate328(.a(gate177inter12), .b(gate177inter1), .O(N730));

  xor2  gate441(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate442(.a(gate178inter0), .b(s_34), .O(gate178inter1));
  and2  gate443(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate444(.a(s_34), .O(gate178inter3));
  inv1  gate445(.a(s_35), .O(gate178inter4));
  nand2 gate446(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate447(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate448(.a(N29), .O(gate178inter7));
  inv1  gate449(.a(N699), .O(gate178inter8));
  nand2 gate450(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate451(.a(s_35), .b(gate178inter3), .O(gate178inter10));
  nor2  gate452(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate453(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate454(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );

  xor2  gate329(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate330(.a(gate183inter0), .b(s_18), .O(gate183inter1));
  and2  gate331(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate332(.a(s_18), .O(gate183inter3));
  inv1  gate333(.a(s_19), .O(gate183inter4));
  nand2 gate334(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate335(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate336(.a(N49), .O(gate183inter7));
  inv1  gate337(.a(N704), .O(gate183inter8));
  nand2 gate338(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate339(.a(s_19), .b(gate183inter3), .O(gate183inter10));
  nor2  gate340(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate341(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate342(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate455(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate456(.a(gate186inter0), .b(s_36), .O(gate186inter1));
  and2  gate457(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate458(.a(s_36), .O(gate186inter3));
  inv1  gate459(.a(s_37), .O(gate186inter4));
  nand2 gate460(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate461(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate462(.a(N61), .O(gate186inter7));
  inv1  gate463(.a(N707), .O(gate186inter8));
  nand2 gate464(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate465(.a(s_37), .b(gate186inter3), .O(gate186inter10));
  nor2  gate466(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate467(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate468(.a(gate186inter12), .b(gate186inter1), .O(N739));
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );

  xor2  gate399(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate400(.a(gate195inter0), .b(s_28), .O(gate195inter1));
  and2  gate401(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate402(.a(s_28), .O(gate195inter3));
  inv1  gate403(.a(s_29), .O(gate195inter4));
  nand2 gate404(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate405(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate406(.a(N97), .O(gate195inter7));
  inv1  gate407(.a(N716), .O(gate195inter8));
  nand2 gate408(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate409(.a(s_29), .b(gate195inter3), .O(gate195inter10));
  nor2  gate410(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate411(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate412(.a(gate195inter12), .b(gate195inter1), .O(N748));
xor2 gate196( .a(N101), .b(N717), .O(N749) );

  xor2  gate217(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate218(.a(gate197inter0), .b(s_2), .O(gate197inter1));
  and2  gate219(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate220(.a(s_2), .O(gate197inter3));
  inv1  gate221(.a(s_3), .O(gate197inter4));
  nand2 gate222(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate223(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate224(.a(N105), .O(gate197inter7));
  inv1  gate225(.a(N718), .O(gate197inter8));
  nand2 gate226(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate227(.a(s_3), .b(gate197inter3), .O(gate197inter10));
  nor2  gate228(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate229(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate230(.a(gate197inter12), .b(gate197inter1), .O(N750));

  xor2  gate469(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate470(.a(gate198inter0), .b(s_38), .O(gate198inter1));
  and2  gate471(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate472(.a(s_38), .O(gate198inter3));
  inv1  gate473(.a(s_39), .O(gate198inter4));
  nand2 gate474(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate475(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate476(.a(N109), .O(gate198inter7));
  inv1  gate477(.a(N719), .O(gate198inter8));
  nand2 gate478(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate479(.a(s_39), .b(gate198inter3), .O(gate198inter10));
  nor2  gate480(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate481(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate482(.a(gate198inter12), .b(gate198inter1), .O(N751));
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule