module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate259(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate260(.a(gate29inter0), .b(s_14), .O(gate29inter1));
  and2  gate261(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate262(.a(s_14), .O(gate29inter3));
  inv1  gate263(.a(s_15), .O(gate29inter4));
  nand2 gate264(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate265(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate266(.a(N150), .O(gate29inter7));
  inv1  gate267(.a(N108), .O(gate29inter8));
  nand2 gate268(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate269(.a(s_15), .b(gate29inter3), .O(gate29inter10));
  nor2  gate270(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate271(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate272(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );

  xor2  gate273(.a(N127), .b(N40), .O(gate33inter0));
  nand2 gate274(.a(gate33inter0), .b(s_16), .O(gate33inter1));
  and2  gate275(.a(N127), .b(N40), .O(gate33inter2));
  inv1  gate276(.a(s_16), .O(gate33inter3));
  inv1  gate277(.a(s_17), .O(gate33inter4));
  nand2 gate278(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate279(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate280(.a(N40), .O(gate33inter7));
  inv1  gate281(.a(N127), .O(gate33inter8));
  nand2 gate282(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate283(.a(s_17), .b(gate33inter3), .O(gate33inter10));
  nor2  gate284(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate285(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate286(.a(gate33inter12), .b(gate33inter1), .O(N186));
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );

  xor2  gate217(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate218(.a(gate39inter0), .b(s_8), .O(gate39inter1));
  and2  gate219(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate220(.a(s_8), .O(gate39inter3));
  inv1  gate221(.a(s_9), .O(gate39inter4));
  nand2 gate222(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate223(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate224(.a(N79), .O(gate39inter7));
  inv1  gate225(.a(N139), .O(gate39inter8));
  nand2 gate226(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate227(.a(s_9), .b(gate39inter3), .O(gate39inter10));
  nor2  gate228(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate229(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate230(.a(gate39inter12), .b(gate39inter1), .O(N192));
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );

  xor2  gate343(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate344(.a(gate42inter0), .b(s_26), .O(gate42inter1));
  and2  gate345(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate346(.a(s_26), .O(gate42inter3));
  inv1  gate347(.a(s_27), .O(gate42inter4));
  nand2 gate348(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate349(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate350(.a(N99), .O(gate42inter7));
  inv1  gate351(.a(N147), .O(gate42inter8));
  nand2 gate352(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate353(.a(s_27), .b(gate42inter3), .O(gate42inter10));
  nor2  gate354(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate355(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate356(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );

  xor2  gate175(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate176(.a(gate51inter0), .b(s_2), .O(gate51inter1));
  and2  gate177(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate178(.a(s_2), .O(gate51inter3));
  inv1  gate179(.a(s_3), .O(gate51inter4));
  nand2 gate180(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate181(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate182(.a(N203), .O(gate51inter7));
  inv1  gate183(.a(N159), .O(gate51inter8));
  nand2 gate184(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate185(.a(s_3), .b(gate51inter3), .O(gate51inter10));
  nor2  gate186(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate187(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate188(.a(gate51inter12), .b(gate51inter1), .O(N227));

  xor2  gate189(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate190(.a(gate52inter0), .b(s_4), .O(gate52inter1));
  and2  gate191(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate192(.a(s_4), .O(gate52inter3));
  inv1  gate193(.a(s_5), .O(gate52inter4));
  nand2 gate194(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate195(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate196(.a(N203), .O(gate52inter7));
  inv1  gate197(.a(N162), .O(gate52inter8));
  nand2 gate198(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate199(.a(s_5), .b(gate52inter3), .O(gate52inter10));
  nor2  gate200(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate201(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate202(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate161(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate162(.a(gate59inter0), .b(s_0), .O(gate59inter1));
  and2  gate163(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate164(.a(s_0), .O(gate59inter3));
  inv1  gate165(.a(s_1), .O(gate59inter4));
  nand2 gate166(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate167(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate168(.a(N203), .O(gate59inter7));
  inv1  gate169(.a(N177), .O(gate59inter8));
  nand2 gate170(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate171(.a(s_1), .b(gate59inter3), .O(gate59inter10));
  nor2  gate172(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate173(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate174(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );

  xor2  gate203(.a(N180), .b(N203), .O(gate61inter0));
  nand2 gate204(.a(gate61inter0), .b(s_6), .O(gate61inter1));
  and2  gate205(.a(N180), .b(N203), .O(gate61inter2));
  inv1  gate206(.a(s_6), .O(gate61inter3));
  inv1  gate207(.a(s_7), .O(gate61inter4));
  nand2 gate208(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate209(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate210(.a(N203), .O(gate61inter7));
  inv1  gate211(.a(N180), .O(gate61inter8));
  nand2 gate212(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate213(.a(s_7), .b(gate61inter3), .O(gate61inter10));
  nor2  gate214(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate215(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate216(.a(gate61inter12), .b(gate61inter1), .O(N251));
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate357(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate358(.a(gate65inter0), .b(s_28), .O(gate65inter1));
  and2  gate359(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate360(.a(s_28), .O(gate65inter3));
  inv1  gate361(.a(s_29), .O(gate65inter4));
  nand2 gate362(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate363(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate364(.a(N213), .O(gate65inter7));
  inv1  gate365(.a(N76), .O(gate65inter8));
  nand2 gate366(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate367(.a(s_29), .b(gate65inter3), .O(gate65inter10));
  nor2  gate368(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate369(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate370(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate245(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate246(.a(gate68inter0), .b(s_12), .O(gate68inter1));
  and2  gate247(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate248(.a(s_12), .O(gate68inter3));
  inv1  gate249(.a(s_13), .O(gate68inter4));
  nand2 gate250(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate251(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate252(.a(N224), .O(gate68inter7));
  inv1  gate253(.a(N157), .O(gate68inter8));
  nand2 gate254(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate255(.a(s_13), .b(gate68inter3), .O(gate68inter10));
  nor2  gate256(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate257(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate258(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate287(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate288(.a(gate75inter0), .b(s_18), .O(gate75inter1));
  and2  gate289(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate290(.a(s_18), .O(gate75inter3));
  inv1  gate291(.a(s_19), .O(gate75inter4));
  nand2 gate292(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate293(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate294(.a(N243), .O(gate75inter7));
  inv1  gate295(.a(N193), .O(gate75inter8));
  nand2 gate296(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate297(.a(s_19), .b(gate75inter3), .O(gate75inter10));
  nor2  gate298(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate299(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate300(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate231(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate232(.a(gate105inter0), .b(s_10), .O(gate105inter1));
  and2  gate233(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate234(.a(s_10), .O(gate105inter3));
  inv1  gate235(.a(s_11), .O(gate105inter4));
  nand2 gate236(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate237(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate238(.a(N319), .O(gate105inter7));
  inv1  gate239(.a(N21), .O(gate105inter8));
  nand2 gate240(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate241(.a(s_11), .b(gate105inter3), .O(gate105inter10));
  nor2  gate242(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate243(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate244(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate301(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate302(.a(gate113inter0), .b(s_20), .O(gate113inter1));
  and2  gate303(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate304(.a(s_20), .O(gate113inter3));
  inv1  gate305(.a(s_21), .O(gate113inter4));
  nand2 gate306(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate307(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate308(.a(N319), .O(gate113inter7));
  inv1  gate309(.a(N73), .O(gate113inter8));
  nand2 gate310(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate311(.a(s_21), .b(gate113inter3), .O(gate113inter10));
  nor2  gate312(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate313(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate314(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate315(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate316(.a(gate119inter0), .b(s_22), .O(gate119inter1));
  and2  gate317(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate318(.a(s_22), .O(gate119inter3));
  inv1  gate319(.a(s_23), .O(gate119inter4));
  nand2 gate320(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate321(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate322(.a(N332), .O(gate119inter7));
  inv1  gate323(.a(N302), .O(gate119inter8));
  nand2 gate324(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate325(.a(s_23), .b(gate119inter3), .O(gate119inter10));
  nor2  gate326(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate327(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate328(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );

  xor2  gate329(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate330(.a(gate130inter0), .b(s_24), .O(gate130inter1));
  and2  gate331(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate332(.a(s_24), .O(gate130inter3));
  inv1  gate333(.a(s_25), .O(gate130inter4));
  nand2 gate334(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate335(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate336(.a(N360), .O(gate130inter7));
  inv1  gate337(.a(N27), .O(gate130inter8));
  nand2 gate338(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate339(.a(s_25), .b(gate130inter3), .O(gate130inter10));
  nor2  gate340(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate341(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate342(.a(gate130inter12), .b(gate130inter1), .O(N372));
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );

  xor2  gate371(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate372(.a(gate137inter0), .b(s_30), .O(gate137inter1));
  and2  gate373(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate374(.a(s_30), .O(gate137inter3));
  inv1  gate375(.a(s_31), .O(gate137inter4));
  nand2 gate376(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate377(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate378(.a(N360), .O(gate137inter7));
  inv1  gate379(.a(N115), .O(gate137inter8));
  nand2 gate380(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate381(.a(s_31), .b(gate137inter3), .O(gate137inter10));
  nor2  gate382(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate383(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate384(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule