module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1303(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1304(.a(gate11inter0), .b(s_108), .O(gate11inter1));
  and2  gate1305(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1306(.a(s_108), .O(gate11inter3));
  inv1  gate1307(.a(s_109), .O(gate11inter4));
  nand2 gate1308(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1309(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1310(.a(G5), .O(gate11inter7));
  inv1  gate1311(.a(G6), .O(gate11inter8));
  nand2 gate1312(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1313(.a(s_109), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1314(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1315(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1316(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1723(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1724(.a(gate12inter0), .b(s_168), .O(gate12inter1));
  and2  gate1725(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1726(.a(s_168), .O(gate12inter3));
  inv1  gate1727(.a(s_169), .O(gate12inter4));
  nand2 gate1728(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1729(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1730(.a(G7), .O(gate12inter7));
  inv1  gate1731(.a(G8), .O(gate12inter8));
  nand2 gate1732(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1733(.a(s_169), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1734(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1735(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1736(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1541(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1542(.a(gate17inter0), .b(s_142), .O(gate17inter1));
  and2  gate1543(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1544(.a(s_142), .O(gate17inter3));
  inv1  gate1545(.a(s_143), .O(gate17inter4));
  nand2 gate1546(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1547(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1548(.a(G17), .O(gate17inter7));
  inv1  gate1549(.a(G18), .O(gate17inter8));
  nand2 gate1550(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1551(.a(s_143), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1552(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1553(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1554(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1499(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1500(.a(gate33inter0), .b(s_136), .O(gate33inter1));
  and2  gate1501(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1502(.a(s_136), .O(gate33inter3));
  inv1  gate1503(.a(s_137), .O(gate33inter4));
  nand2 gate1504(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1505(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1506(.a(G17), .O(gate33inter7));
  inv1  gate1507(.a(G21), .O(gate33inter8));
  nand2 gate1508(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1509(.a(s_137), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1510(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1511(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1512(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1051(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1052(.a(gate45inter0), .b(s_72), .O(gate45inter1));
  and2  gate1053(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1054(.a(s_72), .O(gate45inter3));
  inv1  gate1055(.a(s_73), .O(gate45inter4));
  nand2 gate1056(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1057(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1058(.a(G5), .O(gate45inter7));
  inv1  gate1059(.a(G272), .O(gate45inter8));
  nand2 gate1060(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1061(.a(s_73), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1062(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1063(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1064(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1709(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1710(.a(gate47inter0), .b(s_166), .O(gate47inter1));
  and2  gate1711(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1712(.a(s_166), .O(gate47inter3));
  inv1  gate1713(.a(s_167), .O(gate47inter4));
  nand2 gate1714(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1715(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1716(.a(G7), .O(gate47inter7));
  inv1  gate1717(.a(G275), .O(gate47inter8));
  nand2 gate1718(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1719(.a(s_167), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1720(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1721(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1722(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate659(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate660(.a(gate52inter0), .b(s_16), .O(gate52inter1));
  and2  gate661(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate662(.a(s_16), .O(gate52inter3));
  inv1  gate663(.a(s_17), .O(gate52inter4));
  nand2 gate664(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate665(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate666(.a(G12), .O(gate52inter7));
  inv1  gate667(.a(G281), .O(gate52inter8));
  nand2 gate668(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate669(.a(s_17), .b(gate52inter3), .O(gate52inter10));
  nor2  gate670(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate671(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate672(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate897(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate898(.a(gate55inter0), .b(s_50), .O(gate55inter1));
  and2  gate899(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate900(.a(s_50), .O(gate55inter3));
  inv1  gate901(.a(s_51), .O(gate55inter4));
  nand2 gate902(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate903(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate904(.a(G15), .O(gate55inter7));
  inv1  gate905(.a(G287), .O(gate55inter8));
  nand2 gate906(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate907(.a(s_51), .b(gate55inter3), .O(gate55inter10));
  nor2  gate908(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate909(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate910(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate813(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate814(.a(gate56inter0), .b(s_38), .O(gate56inter1));
  and2  gate815(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate816(.a(s_38), .O(gate56inter3));
  inv1  gate817(.a(s_39), .O(gate56inter4));
  nand2 gate818(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate819(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate820(.a(G16), .O(gate56inter7));
  inv1  gate821(.a(G287), .O(gate56inter8));
  nand2 gate822(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate823(.a(s_39), .b(gate56inter3), .O(gate56inter10));
  nor2  gate824(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate825(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate826(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate785(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate786(.a(gate60inter0), .b(s_34), .O(gate60inter1));
  and2  gate787(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate788(.a(s_34), .O(gate60inter3));
  inv1  gate789(.a(s_35), .O(gate60inter4));
  nand2 gate790(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate791(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate792(.a(G20), .O(gate60inter7));
  inv1  gate793(.a(G293), .O(gate60inter8));
  nand2 gate794(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate795(.a(s_35), .b(gate60inter3), .O(gate60inter10));
  nor2  gate796(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate797(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate798(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1079(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1080(.a(gate79inter0), .b(s_76), .O(gate79inter1));
  and2  gate1081(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1082(.a(s_76), .O(gate79inter3));
  inv1  gate1083(.a(s_77), .O(gate79inter4));
  nand2 gate1084(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1085(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1086(.a(G10), .O(gate79inter7));
  inv1  gate1087(.a(G323), .O(gate79inter8));
  nand2 gate1088(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1089(.a(s_77), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1090(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1091(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1092(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1093(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1094(.a(gate81inter0), .b(s_78), .O(gate81inter1));
  and2  gate1095(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1096(.a(s_78), .O(gate81inter3));
  inv1  gate1097(.a(s_79), .O(gate81inter4));
  nand2 gate1098(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1099(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1100(.a(G3), .O(gate81inter7));
  inv1  gate1101(.a(G326), .O(gate81inter8));
  nand2 gate1102(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1103(.a(s_79), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1104(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1105(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1106(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1569(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1570(.a(gate83inter0), .b(s_146), .O(gate83inter1));
  and2  gate1571(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1572(.a(s_146), .O(gate83inter3));
  inv1  gate1573(.a(s_147), .O(gate83inter4));
  nand2 gate1574(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1575(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1576(.a(G11), .O(gate83inter7));
  inv1  gate1577(.a(G329), .O(gate83inter8));
  nand2 gate1578(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1579(.a(s_147), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1580(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1581(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1582(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1135(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1136(.a(gate94inter0), .b(s_84), .O(gate94inter1));
  and2  gate1137(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1138(.a(s_84), .O(gate94inter3));
  inv1  gate1139(.a(s_85), .O(gate94inter4));
  nand2 gate1140(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1141(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1142(.a(G22), .O(gate94inter7));
  inv1  gate1143(.a(G344), .O(gate94inter8));
  nand2 gate1144(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1145(.a(s_85), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1146(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1147(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1148(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1373(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1374(.a(gate95inter0), .b(s_118), .O(gate95inter1));
  and2  gate1375(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1376(.a(s_118), .O(gate95inter3));
  inv1  gate1377(.a(s_119), .O(gate95inter4));
  nand2 gate1378(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1379(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1380(.a(G26), .O(gate95inter7));
  inv1  gate1381(.a(G347), .O(gate95inter8));
  nand2 gate1382(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1383(.a(s_119), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1384(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1385(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1386(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate841(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate842(.a(gate99inter0), .b(s_42), .O(gate99inter1));
  and2  gate843(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate844(.a(s_42), .O(gate99inter3));
  inv1  gate845(.a(s_43), .O(gate99inter4));
  nand2 gate846(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate847(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate848(.a(G27), .O(gate99inter7));
  inv1  gate849(.a(G353), .O(gate99inter8));
  nand2 gate850(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate851(.a(s_43), .b(gate99inter3), .O(gate99inter10));
  nor2  gate852(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate853(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate854(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1177(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1178(.a(gate104inter0), .b(s_90), .O(gate104inter1));
  and2  gate1179(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1180(.a(s_90), .O(gate104inter3));
  inv1  gate1181(.a(s_91), .O(gate104inter4));
  nand2 gate1182(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1183(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1184(.a(G32), .O(gate104inter7));
  inv1  gate1185(.a(G359), .O(gate104inter8));
  nand2 gate1186(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1187(.a(s_91), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1188(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1189(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1190(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1555(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1556(.a(gate106inter0), .b(s_144), .O(gate106inter1));
  and2  gate1557(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1558(.a(s_144), .O(gate106inter3));
  inv1  gate1559(.a(s_145), .O(gate106inter4));
  nand2 gate1560(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1561(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1562(.a(G364), .O(gate106inter7));
  inv1  gate1563(.a(G365), .O(gate106inter8));
  nand2 gate1564(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1565(.a(s_145), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1566(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1567(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1568(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1415(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1416(.a(gate107inter0), .b(s_124), .O(gate107inter1));
  and2  gate1417(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1418(.a(s_124), .O(gate107inter3));
  inv1  gate1419(.a(s_125), .O(gate107inter4));
  nand2 gate1420(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1421(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1422(.a(G366), .O(gate107inter7));
  inv1  gate1423(.a(G367), .O(gate107inter8));
  nand2 gate1424(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1425(.a(s_125), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1426(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1427(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1428(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate631(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate632(.a(gate108inter0), .b(s_12), .O(gate108inter1));
  and2  gate633(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate634(.a(s_12), .O(gate108inter3));
  inv1  gate635(.a(s_13), .O(gate108inter4));
  nand2 gate636(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate637(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate638(.a(G368), .O(gate108inter7));
  inv1  gate639(.a(G369), .O(gate108inter8));
  nand2 gate640(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate641(.a(s_13), .b(gate108inter3), .O(gate108inter10));
  nor2  gate642(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate643(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate644(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate547(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate548(.a(gate109inter0), .b(s_0), .O(gate109inter1));
  and2  gate549(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate550(.a(s_0), .O(gate109inter3));
  inv1  gate551(.a(s_1), .O(gate109inter4));
  nand2 gate552(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate553(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate554(.a(G370), .O(gate109inter7));
  inv1  gate555(.a(G371), .O(gate109inter8));
  nand2 gate556(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate557(.a(s_1), .b(gate109inter3), .O(gate109inter10));
  nor2  gate558(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate559(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate560(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate603(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate604(.a(gate116inter0), .b(s_8), .O(gate116inter1));
  and2  gate605(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate606(.a(s_8), .O(gate116inter3));
  inv1  gate607(.a(s_9), .O(gate116inter4));
  nand2 gate608(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate609(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate610(.a(G384), .O(gate116inter7));
  inv1  gate611(.a(G385), .O(gate116inter8));
  nand2 gate612(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate613(.a(s_9), .b(gate116inter3), .O(gate116inter10));
  nor2  gate614(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate615(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate616(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate883(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate884(.a(gate118inter0), .b(s_48), .O(gate118inter1));
  and2  gate885(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate886(.a(s_48), .O(gate118inter3));
  inv1  gate887(.a(s_49), .O(gate118inter4));
  nand2 gate888(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate889(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate890(.a(G388), .O(gate118inter7));
  inv1  gate891(.a(G389), .O(gate118inter8));
  nand2 gate892(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate893(.a(s_49), .b(gate118inter3), .O(gate118inter10));
  nor2  gate894(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate895(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate896(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1023(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1024(.a(gate119inter0), .b(s_68), .O(gate119inter1));
  and2  gate1025(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1026(.a(s_68), .O(gate119inter3));
  inv1  gate1027(.a(s_69), .O(gate119inter4));
  nand2 gate1028(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1029(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1030(.a(G390), .O(gate119inter7));
  inv1  gate1031(.a(G391), .O(gate119inter8));
  nand2 gate1032(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1033(.a(s_69), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1034(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1035(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1036(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate827(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate828(.a(gate128inter0), .b(s_40), .O(gate128inter1));
  and2  gate829(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate830(.a(s_40), .O(gate128inter3));
  inv1  gate831(.a(s_41), .O(gate128inter4));
  nand2 gate832(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate833(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate834(.a(G408), .O(gate128inter7));
  inv1  gate835(.a(G409), .O(gate128inter8));
  nand2 gate836(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate837(.a(s_41), .b(gate128inter3), .O(gate128inter10));
  nor2  gate838(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate839(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate840(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1471(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1472(.a(gate130inter0), .b(s_132), .O(gate130inter1));
  and2  gate1473(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1474(.a(s_132), .O(gate130inter3));
  inv1  gate1475(.a(s_133), .O(gate130inter4));
  nand2 gate1476(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1477(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1478(.a(G412), .O(gate130inter7));
  inv1  gate1479(.a(G413), .O(gate130inter8));
  nand2 gate1480(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1481(.a(s_133), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1482(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1483(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1484(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1625(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1626(.a(gate136inter0), .b(s_154), .O(gate136inter1));
  and2  gate1627(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1628(.a(s_154), .O(gate136inter3));
  inv1  gate1629(.a(s_155), .O(gate136inter4));
  nand2 gate1630(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1631(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1632(.a(G424), .O(gate136inter7));
  inv1  gate1633(.a(G425), .O(gate136inter8));
  nand2 gate1634(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1635(.a(s_155), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1636(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1637(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1638(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1387(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1388(.a(gate143inter0), .b(s_120), .O(gate143inter1));
  and2  gate1389(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1390(.a(s_120), .O(gate143inter3));
  inv1  gate1391(.a(s_121), .O(gate143inter4));
  nand2 gate1392(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1393(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1394(.a(G462), .O(gate143inter7));
  inv1  gate1395(.a(G465), .O(gate143inter8));
  nand2 gate1396(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1397(.a(s_121), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1398(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1399(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1400(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1275(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1276(.a(gate147inter0), .b(s_104), .O(gate147inter1));
  and2  gate1277(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1278(.a(s_104), .O(gate147inter3));
  inv1  gate1279(.a(s_105), .O(gate147inter4));
  nand2 gate1280(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1281(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1282(.a(G486), .O(gate147inter7));
  inv1  gate1283(.a(G489), .O(gate147inter8));
  nand2 gate1284(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1285(.a(s_105), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1286(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1287(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1288(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1289(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1290(.a(gate152inter0), .b(s_106), .O(gate152inter1));
  and2  gate1291(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1292(.a(s_106), .O(gate152inter3));
  inv1  gate1293(.a(s_107), .O(gate152inter4));
  nand2 gate1294(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1295(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1296(.a(G516), .O(gate152inter7));
  inv1  gate1297(.a(G519), .O(gate152inter8));
  nand2 gate1298(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1299(.a(s_107), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1300(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1301(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1302(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate743(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate744(.a(gate159inter0), .b(s_28), .O(gate159inter1));
  and2  gate745(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate746(.a(s_28), .O(gate159inter3));
  inv1  gate747(.a(s_29), .O(gate159inter4));
  nand2 gate748(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate749(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate750(.a(G444), .O(gate159inter7));
  inv1  gate751(.a(G531), .O(gate159inter8));
  nand2 gate752(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate753(.a(s_29), .b(gate159inter3), .O(gate159inter10));
  nor2  gate754(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate755(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate756(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1653(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1654(.a(gate170inter0), .b(s_158), .O(gate170inter1));
  and2  gate1655(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1656(.a(s_158), .O(gate170inter3));
  inv1  gate1657(.a(s_159), .O(gate170inter4));
  nand2 gate1658(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1659(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1660(.a(G477), .O(gate170inter7));
  inv1  gate1661(.a(G546), .O(gate170inter8));
  nand2 gate1662(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1663(.a(s_159), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1664(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1665(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1666(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1695(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1696(.a(gate171inter0), .b(s_164), .O(gate171inter1));
  and2  gate1697(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1698(.a(s_164), .O(gate171inter3));
  inv1  gate1699(.a(s_165), .O(gate171inter4));
  nand2 gate1700(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1701(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1702(.a(G480), .O(gate171inter7));
  inv1  gate1703(.a(G549), .O(gate171inter8));
  nand2 gate1704(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1705(.a(s_165), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1706(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1707(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1708(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1107(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1108(.a(gate172inter0), .b(s_80), .O(gate172inter1));
  and2  gate1109(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1110(.a(s_80), .O(gate172inter3));
  inv1  gate1111(.a(s_81), .O(gate172inter4));
  nand2 gate1112(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1113(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1114(.a(G483), .O(gate172inter7));
  inv1  gate1115(.a(G549), .O(gate172inter8));
  nand2 gate1116(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1117(.a(s_81), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1118(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1119(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1120(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1121(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1122(.a(gate174inter0), .b(s_82), .O(gate174inter1));
  and2  gate1123(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1124(.a(s_82), .O(gate174inter3));
  inv1  gate1125(.a(s_83), .O(gate174inter4));
  nand2 gate1126(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1127(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1128(.a(G489), .O(gate174inter7));
  inv1  gate1129(.a(G552), .O(gate174inter8));
  nand2 gate1130(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1131(.a(s_83), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1132(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1133(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1134(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1597(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1598(.a(gate175inter0), .b(s_150), .O(gate175inter1));
  and2  gate1599(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1600(.a(s_150), .O(gate175inter3));
  inv1  gate1601(.a(s_151), .O(gate175inter4));
  nand2 gate1602(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1603(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1604(.a(G492), .O(gate175inter7));
  inv1  gate1605(.a(G555), .O(gate175inter8));
  nand2 gate1606(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1607(.a(s_151), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1608(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1609(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1610(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate575(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate576(.a(gate178inter0), .b(s_4), .O(gate178inter1));
  and2  gate577(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate578(.a(s_4), .O(gate178inter3));
  inv1  gate579(.a(s_5), .O(gate178inter4));
  nand2 gate580(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate581(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate582(.a(G501), .O(gate178inter7));
  inv1  gate583(.a(G558), .O(gate178inter8));
  nand2 gate584(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate585(.a(s_5), .b(gate178inter3), .O(gate178inter10));
  nor2  gate586(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate587(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate588(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate939(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate940(.a(gate179inter0), .b(s_56), .O(gate179inter1));
  and2  gate941(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate942(.a(s_56), .O(gate179inter3));
  inv1  gate943(.a(s_57), .O(gate179inter4));
  nand2 gate944(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate945(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate946(.a(G504), .O(gate179inter7));
  inv1  gate947(.a(G561), .O(gate179inter8));
  nand2 gate948(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate949(.a(s_57), .b(gate179inter3), .O(gate179inter10));
  nor2  gate950(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate951(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate952(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1737(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1738(.a(gate182inter0), .b(s_170), .O(gate182inter1));
  and2  gate1739(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1740(.a(s_170), .O(gate182inter3));
  inv1  gate1741(.a(s_171), .O(gate182inter4));
  nand2 gate1742(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1743(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1744(.a(G513), .O(gate182inter7));
  inv1  gate1745(.a(G564), .O(gate182inter8));
  nand2 gate1746(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1747(.a(s_171), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1748(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1749(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1750(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1331(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1332(.a(gate191inter0), .b(s_112), .O(gate191inter1));
  and2  gate1333(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1334(.a(s_112), .O(gate191inter3));
  inv1  gate1335(.a(s_113), .O(gate191inter4));
  nand2 gate1336(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1337(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1338(.a(G582), .O(gate191inter7));
  inv1  gate1339(.a(G583), .O(gate191inter8));
  nand2 gate1340(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1341(.a(s_113), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1342(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1343(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1344(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1457(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1458(.a(gate202inter0), .b(s_130), .O(gate202inter1));
  and2  gate1459(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1460(.a(s_130), .O(gate202inter3));
  inv1  gate1461(.a(s_131), .O(gate202inter4));
  nand2 gate1462(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1463(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1464(.a(G612), .O(gate202inter7));
  inv1  gate1465(.a(G617), .O(gate202inter8));
  nand2 gate1466(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1467(.a(s_131), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1468(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1469(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1470(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate869(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate870(.a(gate214inter0), .b(s_46), .O(gate214inter1));
  and2  gate871(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate872(.a(s_46), .O(gate214inter3));
  inv1  gate873(.a(s_47), .O(gate214inter4));
  nand2 gate874(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate875(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate876(.a(G612), .O(gate214inter7));
  inv1  gate877(.a(G672), .O(gate214inter8));
  nand2 gate878(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate879(.a(s_47), .b(gate214inter3), .O(gate214inter10));
  nor2  gate880(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate881(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate882(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate995(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate996(.a(gate218inter0), .b(s_64), .O(gate218inter1));
  and2  gate997(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate998(.a(s_64), .O(gate218inter3));
  inv1  gate999(.a(s_65), .O(gate218inter4));
  nand2 gate1000(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1001(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1002(.a(G627), .O(gate218inter7));
  inv1  gate1003(.a(G678), .O(gate218inter8));
  nand2 gate1004(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1005(.a(s_65), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1006(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1007(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1008(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate715(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate716(.a(gate230inter0), .b(s_24), .O(gate230inter1));
  and2  gate717(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate718(.a(s_24), .O(gate230inter3));
  inv1  gate719(.a(s_25), .O(gate230inter4));
  nand2 gate720(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate721(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate722(.a(G700), .O(gate230inter7));
  inv1  gate723(.a(G701), .O(gate230inter8));
  nand2 gate724(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate725(.a(s_25), .b(gate230inter3), .O(gate230inter10));
  nor2  gate726(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate727(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate728(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1401(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1402(.a(gate233inter0), .b(s_122), .O(gate233inter1));
  and2  gate1403(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1404(.a(s_122), .O(gate233inter3));
  inv1  gate1405(.a(s_123), .O(gate233inter4));
  nand2 gate1406(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1407(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1408(.a(G242), .O(gate233inter7));
  inv1  gate1409(.a(G718), .O(gate233inter8));
  nand2 gate1410(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1411(.a(s_123), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1412(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1413(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1414(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate855(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate856(.a(gate238inter0), .b(s_44), .O(gate238inter1));
  and2  gate857(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate858(.a(s_44), .O(gate238inter3));
  inv1  gate859(.a(s_45), .O(gate238inter4));
  nand2 gate860(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate861(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate862(.a(G257), .O(gate238inter7));
  inv1  gate863(.a(G709), .O(gate238inter8));
  nand2 gate864(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate865(.a(s_45), .b(gate238inter3), .O(gate238inter10));
  nor2  gate866(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate867(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate868(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1429(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1430(.a(gate240inter0), .b(s_126), .O(gate240inter1));
  and2  gate1431(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1432(.a(s_126), .O(gate240inter3));
  inv1  gate1433(.a(s_127), .O(gate240inter4));
  nand2 gate1434(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1435(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1436(.a(G263), .O(gate240inter7));
  inv1  gate1437(.a(G715), .O(gate240inter8));
  nand2 gate1438(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1439(.a(s_127), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1440(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1441(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1442(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1065(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1066(.a(gate243inter0), .b(s_74), .O(gate243inter1));
  and2  gate1067(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1068(.a(s_74), .O(gate243inter3));
  inv1  gate1069(.a(s_75), .O(gate243inter4));
  nand2 gate1070(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1071(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1072(.a(G245), .O(gate243inter7));
  inv1  gate1073(.a(G733), .O(gate243inter8));
  nand2 gate1074(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1075(.a(s_75), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1076(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1077(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1078(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate925(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate926(.a(gate250inter0), .b(s_54), .O(gate250inter1));
  and2  gate927(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate928(.a(s_54), .O(gate250inter3));
  inv1  gate929(.a(s_55), .O(gate250inter4));
  nand2 gate930(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate931(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate932(.a(G706), .O(gate250inter7));
  inv1  gate933(.a(G742), .O(gate250inter8));
  nand2 gate934(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate935(.a(s_55), .b(gate250inter3), .O(gate250inter10));
  nor2  gate936(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate937(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate938(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate687(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate688(.a(gate252inter0), .b(s_20), .O(gate252inter1));
  and2  gate689(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate690(.a(s_20), .O(gate252inter3));
  inv1  gate691(.a(s_21), .O(gate252inter4));
  nand2 gate692(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate693(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate694(.a(G709), .O(gate252inter7));
  inv1  gate695(.a(G745), .O(gate252inter8));
  nand2 gate696(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate697(.a(s_21), .b(gate252inter3), .O(gate252inter10));
  nor2  gate698(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate699(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate700(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate701(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate702(.a(gate258inter0), .b(s_22), .O(gate258inter1));
  and2  gate703(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate704(.a(s_22), .O(gate258inter3));
  inv1  gate705(.a(s_23), .O(gate258inter4));
  nand2 gate706(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate707(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate708(.a(G756), .O(gate258inter7));
  inv1  gate709(.a(G757), .O(gate258inter8));
  nand2 gate710(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate711(.a(s_23), .b(gate258inter3), .O(gate258inter10));
  nor2  gate712(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate713(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate714(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1345(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1346(.a(gate261inter0), .b(s_114), .O(gate261inter1));
  and2  gate1347(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1348(.a(s_114), .O(gate261inter3));
  inv1  gate1349(.a(s_115), .O(gate261inter4));
  nand2 gate1350(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1351(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1352(.a(G762), .O(gate261inter7));
  inv1  gate1353(.a(G763), .O(gate261inter8));
  nand2 gate1354(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1355(.a(s_115), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1356(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1357(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1358(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate981(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate982(.a(gate262inter0), .b(s_62), .O(gate262inter1));
  and2  gate983(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate984(.a(s_62), .O(gate262inter3));
  inv1  gate985(.a(s_63), .O(gate262inter4));
  nand2 gate986(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate987(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate988(.a(G764), .O(gate262inter7));
  inv1  gate989(.a(G765), .O(gate262inter8));
  nand2 gate990(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate991(.a(s_63), .b(gate262inter3), .O(gate262inter10));
  nor2  gate992(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate993(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate994(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1667(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1668(.a(gate266inter0), .b(s_160), .O(gate266inter1));
  and2  gate1669(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1670(.a(s_160), .O(gate266inter3));
  inv1  gate1671(.a(s_161), .O(gate266inter4));
  nand2 gate1672(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1673(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1674(.a(G645), .O(gate266inter7));
  inv1  gate1675(.a(G773), .O(gate266inter8));
  nand2 gate1676(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1677(.a(s_161), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1678(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1679(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1680(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1681(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1682(.a(gate268inter0), .b(s_162), .O(gate268inter1));
  and2  gate1683(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1684(.a(s_162), .O(gate268inter3));
  inv1  gate1685(.a(s_163), .O(gate268inter4));
  nand2 gate1686(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1687(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1688(.a(G651), .O(gate268inter7));
  inv1  gate1689(.a(G779), .O(gate268inter8));
  nand2 gate1690(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1691(.a(s_163), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1692(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1693(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1694(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1639(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1640(.a(gate271inter0), .b(s_156), .O(gate271inter1));
  and2  gate1641(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1642(.a(s_156), .O(gate271inter3));
  inv1  gate1643(.a(s_157), .O(gate271inter4));
  nand2 gate1644(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1645(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1646(.a(G660), .O(gate271inter7));
  inv1  gate1647(.a(G788), .O(gate271inter8));
  nand2 gate1648(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1649(.a(s_157), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1650(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1651(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1652(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1261(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1262(.a(gate275inter0), .b(s_102), .O(gate275inter1));
  and2  gate1263(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1264(.a(s_102), .O(gate275inter3));
  inv1  gate1265(.a(s_103), .O(gate275inter4));
  nand2 gate1266(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1267(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1268(.a(G645), .O(gate275inter7));
  inv1  gate1269(.a(G797), .O(gate275inter8));
  nand2 gate1270(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1271(.a(s_103), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1272(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1273(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1274(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1513(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1514(.a(gate279inter0), .b(s_138), .O(gate279inter1));
  and2  gate1515(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1516(.a(s_138), .O(gate279inter3));
  inv1  gate1517(.a(s_139), .O(gate279inter4));
  nand2 gate1518(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1519(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1520(.a(G651), .O(gate279inter7));
  inv1  gate1521(.a(G803), .O(gate279inter8));
  nand2 gate1522(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1523(.a(s_139), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1524(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1525(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1526(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1583(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1584(.a(gate282inter0), .b(s_148), .O(gate282inter1));
  and2  gate1585(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1586(.a(s_148), .O(gate282inter3));
  inv1  gate1587(.a(s_149), .O(gate282inter4));
  nand2 gate1588(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1589(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1590(.a(G782), .O(gate282inter7));
  inv1  gate1591(.a(G806), .O(gate282inter8));
  nand2 gate1592(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1593(.a(s_149), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1594(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1595(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1596(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate617(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate618(.a(gate289inter0), .b(s_10), .O(gate289inter1));
  and2  gate619(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate620(.a(s_10), .O(gate289inter3));
  inv1  gate621(.a(s_11), .O(gate289inter4));
  nand2 gate622(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate623(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate624(.a(G818), .O(gate289inter7));
  inv1  gate625(.a(G819), .O(gate289inter8));
  nand2 gate626(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate627(.a(s_11), .b(gate289inter3), .O(gate289inter10));
  nor2  gate628(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate629(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate630(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate953(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate954(.a(gate388inter0), .b(s_58), .O(gate388inter1));
  and2  gate955(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate956(.a(s_58), .O(gate388inter3));
  inv1  gate957(.a(s_59), .O(gate388inter4));
  nand2 gate958(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate959(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate960(.a(G2), .O(gate388inter7));
  inv1  gate961(.a(G1039), .O(gate388inter8));
  nand2 gate962(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate963(.a(s_59), .b(gate388inter3), .O(gate388inter10));
  nor2  gate964(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate965(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate966(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1163(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1164(.a(gate390inter0), .b(s_88), .O(gate390inter1));
  and2  gate1165(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1166(.a(s_88), .O(gate390inter3));
  inv1  gate1167(.a(s_89), .O(gate390inter4));
  nand2 gate1168(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1169(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1170(.a(G4), .O(gate390inter7));
  inv1  gate1171(.a(G1045), .O(gate390inter8));
  nand2 gate1172(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1173(.a(s_89), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1174(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1175(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1176(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1009(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1010(.a(gate402inter0), .b(s_66), .O(gate402inter1));
  and2  gate1011(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1012(.a(s_66), .O(gate402inter3));
  inv1  gate1013(.a(s_67), .O(gate402inter4));
  nand2 gate1014(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1015(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1016(.a(G16), .O(gate402inter7));
  inv1  gate1017(.a(G1081), .O(gate402inter8));
  nand2 gate1018(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1019(.a(s_67), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1020(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1021(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1022(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1219(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1220(.a(gate409inter0), .b(s_96), .O(gate409inter1));
  and2  gate1221(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1222(.a(s_96), .O(gate409inter3));
  inv1  gate1223(.a(s_97), .O(gate409inter4));
  nand2 gate1224(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1225(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1226(.a(G23), .O(gate409inter7));
  inv1  gate1227(.a(G1102), .O(gate409inter8));
  nand2 gate1228(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1229(.a(s_97), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1230(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1231(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1232(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1359(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1360(.a(gate417inter0), .b(s_116), .O(gate417inter1));
  and2  gate1361(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1362(.a(s_116), .O(gate417inter3));
  inv1  gate1363(.a(s_117), .O(gate417inter4));
  nand2 gate1364(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1365(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1366(.a(G31), .O(gate417inter7));
  inv1  gate1367(.a(G1126), .O(gate417inter8));
  nand2 gate1368(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1369(.a(s_117), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1370(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1371(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1372(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1149(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1150(.a(gate420inter0), .b(s_86), .O(gate420inter1));
  and2  gate1151(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1152(.a(s_86), .O(gate420inter3));
  inv1  gate1153(.a(s_87), .O(gate420inter4));
  nand2 gate1154(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1155(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1156(.a(G1036), .O(gate420inter7));
  inv1  gate1157(.a(G1132), .O(gate420inter8));
  nand2 gate1158(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1159(.a(s_87), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1160(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1161(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1162(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1205(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1206(.a(gate425inter0), .b(s_94), .O(gate425inter1));
  and2  gate1207(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1208(.a(s_94), .O(gate425inter3));
  inv1  gate1209(.a(s_95), .O(gate425inter4));
  nand2 gate1210(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1211(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1212(.a(G4), .O(gate425inter7));
  inv1  gate1213(.a(G1141), .O(gate425inter8));
  nand2 gate1214(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1215(.a(s_95), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1216(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1217(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1218(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1443(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1444(.a(gate428inter0), .b(s_128), .O(gate428inter1));
  and2  gate1445(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1446(.a(s_128), .O(gate428inter3));
  inv1  gate1447(.a(s_129), .O(gate428inter4));
  nand2 gate1448(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1449(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1450(.a(G1048), .O(gate428inter7));
  inv1  gate1451(.a(G1144), .O(gate428inter8));
  nand2 gate1452(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1453(.a(s_129), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1454(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1455(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1456(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate729(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate730(.a(gate431inter0), .b(s_26), .O(gate431inter1));
  and2  gate731(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate732(.a(s_26), .O(gate431inter3));
  inv1  gate733(.a(s_27), .O(gate431inter4));
  nand2 gate734(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate735(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate736(.a(G7), .O(gate431inter7));
  inv1  gate737(.a(G1150), .O(gate431inter8));
  nand2 gate738(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate739(.a(s_27), .b(gate431inter3), .O(gate431inter10));
  nor2  gate740(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate741(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate742(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1037(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1038(.a(gate435inter0), .b(s_70), .O(gate435inter1));
  and2  gate1039(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1040(.a(s_70), .O(gate435inter3));
  inv1  gate1041(.a(s_71), .O(gate435inter4));
  nand2 gate1042(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1043(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1044(.a(G9), .O(gate435inter7));
  inv1  gate1045(.a(G1156), .O(gate435inter8));
  nand2 gate1046(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1047(.a(s_71), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1048(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1049(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1050(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate757(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate758(.a(gate445inter0), .b(s_30), .O(gate445inter1));
  and2  gate759(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate760(.a(s_30), .O(gate445inter3));
  inv1  gate761(.a(s_31), .O(gate445inter4));
  nand2 gate762(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate763(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate764(.a(G14), .O(gate445inter7));
  inv1  gate765(.a(G1171), .O(gate445inter8));
  nand2 gate766(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate767(.a(s_31), .b(gate445inter3), .O(gate445inter10));
  nor2  gate768(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate769(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate770(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1527(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1528(.a(gate448inter0), .b(s_140), .O(gate448inter1));
  and2  gate1529(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1530(.a(s_140), .O(gate448inter3));
  inv1  gate1531(.a(s_141), .O(gate448inter4));
  nand2 gate1532(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1533(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1534(.a(G1078), .O(gate448inter7));
  inv1  gate1535(.a(G1174), .O(gate448inter8));
  nand2 gate1536(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1537(.a(s_141), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1538(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1539(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1540(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1611(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1612(.a(gate458inter0), .b(s_152), .O(gate458inter1));
  and2  gate1613(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1614(.a(s_152), .O(gate458inter3));
  inv1  gate1615(.a(s_153), .O(gate458inter4));
  nand2 gate1616(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1617(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1618(.a(G1093), .O(gate458inter7));
  inv1  gate1619(.a(G1189), .O(gate458inter8));
  nand2 gate1620(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1621(.a(s_153), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1622(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1623(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1624(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate799(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate800(.a(gate471inter0), .b(s_36), .O(gate471inter1));
  and2  gate801(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate802(.a(s_36), .O(gate471inter3));
  inv1  gate803(.a(s_37), .O(gate471inter4));
  nand2 gate804(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate805(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate806(.a(G27), .O(gate471inter7));
  inv1  gate807(.a(G1210), .O(gate471inter8));
  nand2 gate808(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate809(.a(s_37), .b(gate471inter3), .O(gate471inter10));
  nor2  gate810(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate811(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate812(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate589(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate590(.a(gate473inter0), .b(s_6), .O(gate473inter1));
  and2  gate591(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate592(.a(s_6), .O(gate473inter3));
  inv1  gate593(.a(s_7), .O(gate473inter4));
  nand2 gate594(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate595(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate596(.a(G28), .O(gate473inter7));
  inv1  gate597(.a(G1213), .O(gate473inter8));
  nand2 gate598(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate599(.a(s_7), .b(gate473inter3), .O(gate473inter10));
  nor2  gate600(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate601(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate602(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate645(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate646(.a(gate477inter0), .b(s_14), .O(gate477inter1));
  and2  gate647(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate648(.a(s_14), .O(gate477inter3));
  inv1  gate649(.a(s_15), .O(gate477inter4));
  nand2 gate650(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate651(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate652(.a(G30), .O(gate477inter7));
  inv1  gate653(.a(G1219), .O(gate477inter8));
  nand2 gate654(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate655(.a(s_15), .b(gate477inter3), .O(gate477inter10));
  nor2  gate656(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate657(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate658(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1247(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1248(.a(gate479inter0), .b(s_100), .O(gate479inter1));
  and2  gate1249(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1250(.a(s_100), .O(gate479inter3));
  inv1  gate1251(.a(s_101), .O(gate479inter4));
  nand2 gate1252(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1253(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1254(.a(G31), .O(gate479inter7));
  inv1  gate1255(.a(G1222), .O(gate479inter8));
  nand2 gate1256(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1257(.a(s_101), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1258(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1259(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1260(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1317(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1318(.a(gate481inter0), .b(s_110), .O(gate481inter1));
  and2  gate1319(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1320(.a(s_110), .O(gate481inter3));
  inv1  gate1321(.a(s_111), .O(gate481inter4));
  nand2 gate1322(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1323(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1324(.a(G32), .O(gate481inter7));
  inv1  gate1325(.a(G1225), .O(gate481inter8));
  nand2 gate1326(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1327(.a(s_111), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1328(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1329(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1330(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate771(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate772(.a(gate484inter0), .b(s_32), .O(gate484inter1));
  and2  gate773(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate774(.a(s_32), .O(gate484inter3));
  inv1  gate775(.a(s_33), .O(gate484inter4));
  nand2 gate776(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate777(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate778(.a(G1230), .O(gate484inter7));
  inv1  gate779(.a(G1231), .O(gate484inter8));
  nand2 gate780(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate781(.a(s_33), .b(gate484inter3), .O(gate484inter10));
  nor2  gate782(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate783(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate784(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1191(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1192(.a(gate490inter0), .b(s_92), .O(gate490inter1));
  and2  gate1193(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1194(.a(s_92), .O(gate490inter3));
  inv1  gate1195(.a(s_93), .O(gate490inter4));
  nand2 gate1196(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1197(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1198(.a(G1242), .O(gate490inter7));
  inv1  gate1199(.a(G1243), .O(gate490inter8));
  nand2 gate1200(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1201(.a(s_93), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1202(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1203(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1204(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate673(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate674(.a(gate491inter0), .b(s_18), .O(gate491inter1));
  and2  gate675(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate676(.a(s_18), .O(gate491inter3));
  inv1  gate677(.a(s_19), .O(gate491inter4));
  nand2 gate678(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate679(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate680(.a(G1244), .O(gate491inter7));
  inv1  gate681(.a(G1245), .O(gate491inter8));
  nand2 gate682(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate683(.a(s_19), .b(gate491inter3), .O(gate491inter10));
  nor2  gate684(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate685(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate686(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate967(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate968(.a(gate496inter0), .b(s_60), .O(gate496inter1));
  and2  gate969(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate970(.a(s_60), .O(gate496inter3));
  inv1  gate971(.a(s_61), .O(gate496inter4));
  nand2 gate972(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate973(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate974(.a(G1254), .O(gate496inter7));
  inv1  gate975(.a(G1255), .O(gate496inter8));
  nand2 gate976(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate977(.a(s_61), .b(gate496inter3), .O(gate496inter10));
  nor2  gate978(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate979(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate980(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1233(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1234(.a(gate497inter0), .b(s_98), .O(gate497inter1));
  and2  gate1235(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1236(.a(s_98), .O(gate497inter3));
  inv1  gate1237(.a(s_99), .O(gate497inter4));
  nand2 gate1238(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1239(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1240(.a(G1256), .O(gate497inter7));
  inv1  gate1241(.a(G1257), .O(gate497inter8));
  nand2 gate1242(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1243(.a(s_99), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1244(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1245(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1246(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate561(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate562(.a(gate500inter0), .b(s_2), .O(gate500inter1));
  and2  gate563(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate564(.a(s_2), .O(gate500inter3));
  inv1  gate565(.a(s_3), .O(gate500inter4));
  nand2 gate566(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate567(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate568(.a(G1262), .O(gate500inter7));
  inv1  gate569(.a(G1263), .O(gate500inter8));
  nand2 gate570(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate571(.a(s_3), .b(gate500inter3), .O(gate500inter10));
  nor2  gate572(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate573(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate574(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1485(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1486(.a(gate502inter0), .b(s_134), .O(gate502inter1));
  and2  gate1487(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1488(.a(s_134), .O(gate502inter3));
  inv1  gate1489(.a(s_135), .O(gate502inter4));
  nand2 gate1490(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1491(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1492(.a(G1266), .O(gate502inter7));
  inv1  gate1493(.a(G1267), .O(gate502inter8));
  nand2 gate1494(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1495(.a(s_135), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1496(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1497(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1498(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate911(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate912(.a(gate509inter0), .b(s_52), .O(gate509inter1));
  and2  gate913(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate914(.a(s_52), .O(gate509inter3));
  inv1  gate915(.a(s_53), .O(gate509inter4));
  nand2 gate916(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate917(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate918(.a(G1280), .O(gate509inter7));
  inv1  gate919(.a(G1281), .O(gate509inter8));
  nand2 gate920(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate921(.a(s_53), .b(gate509inter3), .O(gate509inter10));
  nor2  gate922(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate923(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate924(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule