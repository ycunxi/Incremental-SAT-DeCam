module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate855(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate856(.a(gate16inter0), .b(s_44), .O(gate16inter1));
  and2  gate857(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate858(.a(s_44), .O(gate16inter3));
  inv1  gate859(.a(s_45), .O(gate16inter4));
  nand2 gate860(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate861(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate862(.a(G15), .O(gate16inter7));
  inv1  gate863(.a(G16), .O(gate16inter8));
  nand2 gate864(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate865(.a(s_45), .b(gate16inter3), .O(gate16inter10));
  nor2  gate866(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate867(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate868(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1821(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1822(.a(gate19inter0), .b(s_182), .O(gate19inter1));
  and2  gate1823(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1824(.a(s_182), .O(gate19inter3));
  inv1  gate1825(.a(s_183), .O(gate19inter4));
  nand2 gate1826(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1827(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1828(.a(G21), .O(gate19inter7));
  inv1  gate1829(.a(G22), .O(gate19inter8));
  nand2 gate1830(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1831(.a(s_183), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1832(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1833(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1834(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2423(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2424(.a(gate23inter0), .b(s_268), .O(gate23inter1));
  and2  gate2425(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2426(.a(s_268), .O(gate23inter3));
  inv1  gate2427(.a(s_269), .O(gate23inter4));
  nand2 gate2428(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2429(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2430(.a(G29), .O(gate23inter7));
  inv1  gate2431(.a(G30), .O(gate23inter8));
  nand2 gate2432(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2433(.a(s_269), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2434(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2435(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2436(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate799(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate800(.a(gate25inter0), .b(s_36), .O(gate25inter1));
  and2  gate801(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate802(.a(s_36), .O(gate25inter3));
  inv1  gate803(.a(s_37), .O(gate25inter4));
  nand2 gate804(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate805(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate806(.a(G1), .O(gate25inter7));
  inv1  gate807(.a(G5), .O(gate25inter8));
  nand2 gate808(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate809(.a(s_37), .b(gate25inter3), .O(gate25inter10));
  nor2  gate810(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate811(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate812(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1877(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1878(.a(gate29inter0), .b(s_190), .O(gate29inter1));
  and2  gate1879(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1880(.a(s_190), .O(gate29inter3));
  inv1  gate1881(.a(s_191), .O(gate29inter4));
  nand2 gate1882(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1883(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1884(.a(G3), .O(gate29inter7));
  inv1  gate1885(.a(G7), .O(gate29inter8));
  nand2 gate1886(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1887(.a(s_191), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1888(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1889(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1890(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1457(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1458(.a(gate31inter0), .b(s_130), .O(gate31inter1));
  and2  gate1459(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1460(.a(s_130), .O(gate31inter3));
  inv1  gate1461(.a(s_131), .O(gate31inter4));
  nand2 gate1462(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1463(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1464(.a(G4), .O(gate31inter7));
  inv1  gate1465(.a(G8), .O(gate31inter8));
  nand2 gate1466(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1467(.a(s_131), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1468(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1469(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1470(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1261(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1262(.a(gate32inter0), .b(s_102), .O(gate32inter1));
  and2  gate1263(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1264(.a(s_102), .O(gate32inter3));
  inv1  gate1265(.a(s_103), .O(gate32inter4));
  nand2 gate1266(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1267(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1268(.a(G12), .O(gate32inter7));
  inv1  gate1269(.a(G16), .O(gate32inter8));
  nand2 gate1270(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1271(.a(s_103), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1272(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1273(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1274(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1583(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1584(.a(gate33inter0), .b(s_148), .O(gate33inter1));
  and2  gate1585(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1586(.a(s_148), .O(gate33inter3));
  inv1  gate1587(.a(s_149), .O(gate33inter4));
  nand2 gate1588(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1589(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1590(.a(G17), .O(gate33inter7));
  inv1  gate1591(.a(G21), .O(gate33inter8));
  nand2 gate1592(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1593(.a(s_149), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1594(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1595(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1596(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2339(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2340(.a(gate36inter0), .b(s_256), .O(gate36inter1));
  and2  gate2341(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2342(.a(s_256), .O(gate36inter3));
  inv1  gate2343(.a(s_257), .O(gate36inter4));
  nand2 gate2344(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2345(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2346(.a(G26), .O(gate36inter7));
  inv1  gate2347(.a(G30), .O(gate36inter8));
  nand2 gate2348(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2349(.a(s_257), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2350(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2351(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2352(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1933(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1934(.a(gate38inter0), .b(s_198), .O(gate38inter1));
  and2  gate1935(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1936(.a(s_198), .O(gate38inter3));
  inv1  gate1937(.a(s_199), .O(gate38inter4));
  nand2 gate1938(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1939(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1940(.a(G27), .O(gate38inter7));
  inv1  gate1941(.a(G31), .O(gate38inter8));
  nand2 gate1942(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1943(.a(s_199), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1944(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1945(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1946(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate561(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate562(.a(gate40inter0), .b(s_2), .O(gate40inter1));
  and2  gate563(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate564(.a(s_2), .O(gate40inter3));
  inv1  gate565(.a(s_3), .O(gate40inter4));
  nand2 gate566(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate567(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate568(.a(G28), .O(gate40inter7));
  inv1  gate569(.a(G32), .O(gate40inter8));
  nand2 gate570(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate571(.a(s_3), .b(gate40inter3), .O(gate40inter10));
  nor2  gate572(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate573(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate574(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1569(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1570(.a(gate41inter0), .b(s_146), .O(gate41inter1));
  and2  gate1571(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1572(.a(s_146), .O(gate41inter3));
  inv1  gate1573(.a(s_147), .O(gate41inter4));
  nand2 gate1574(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1575(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1576(.a(G1), .O(gate41inter7));
  inv1  gate1577(.a(G266), .O(gate41inter8));
  nand2 gate1578(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1579(.a(s_147), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1580(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1581(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1582(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1275(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1276(.a(gate44inter0), .b(s_104), .O(gate44inter1));
  and2  gate1277(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1278(.a(s_104), .O(gate44inter3));
  inv1  gate1279(.a(s_105), .O(gate44inter4));
  nand2 gate1280(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1281(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1282(.a(G4), .O(gate44inter7));
  inv1  gate1283(.a(G269), .O(gate44inter8));
  nand2 gate1284(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1285(.a(s_105), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1286(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1287(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1288(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate659(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate660(.a(gate45inter0), .b(s_16), .O(gate45inter1));
  and2  gate661(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate662(.a(s_16), .O(gate45inter3));
  inv1  gate663(.a(s_17), .O(gate45inter4));
  nand2 gate664(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate665(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate666(.a(G5), .O(gate45inter7));
  inv1  gate667(.a(G272), .O(gate45inter8));
  nand2 gate668(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate669(.a(s_17), .b(gate45inter3), .O(gate45inter10));
  nor2  gate670(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate671(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate672(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate827(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate828(.a(gate48inter0), .b(s_40), .O(gate48inter1));
  and2  gate829(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate830(.a(s_40), .O(gate48inter3));
  inv1  gate831(.a(s_41), .O(gate48inter4));
  nand2 gate832(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate833(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate834(.a(G8), .O(gate48inter7));
  inv1  gate835(.a(G275), .O(gate48inter8));
  nand2 gate836(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate837(.a(s_41), .b(gate48inter3), .O(gate48inter10));
  nor2  gate838(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate839(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate840(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1863(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1864(.a(gate49inter0), .b(s_188), .O(gate49inter1));
  and2  gate1865(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1866(.a(s_188), .O(gate49inter3));
  inv1  gate1867(.a(s_189), .O(gate49inter4));
  nand2 gate1868(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1869(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1870(.a(G9), .O(gate49inter7));
  inv1  gate1871(.a(G278), .O(gate49inter8));
  nand2 gate1872(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1873(.a(s_189), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1874(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1875(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1876(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2493(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2494(.a(gate50inter0), .b(s_278), .O(gate50inter1));
  and2  gate2495(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2496(.a(s_278), .O(gate50inter3));
  inv1  gate2497(.a(s_279), .O(gate50inter4));
  nand2 gate2498(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2499(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2500(.a(G10), .O(gate50inter7));
  inv1  gate2501(.a(G278), .O(gate50inter8));
  nand2 gate2502(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2503(.a(s_279), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2504(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2505(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2506(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2507(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2508(.a(gate53inter0), .b(s_280), .O(gate53inter1));
  and2  gate2509(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2510(.a(s_280), .O(gate53inter3));
  inv1  gate2511(.a(s_281), .O(gate53inter4));
  nand2 gate2512(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2513(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2514(.a(G13), .O(gate53inter7));
  inv1  gate2515(.a(G284), .O(gate53inter8));
  nand2 gate2516(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2517(.a(s_281), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2518(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2519(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2520(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1065(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1066(.a(gate54inter0), .b(s_74), .O(gate54inter1));
  and2  gate1067(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1068(.a(s_74), .O(gate54inter3));
  inv1  gate1069(.a(s_75), .O(gate54inter4));
  nand2 gate1070(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1071(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1072(.a(G14), .O(gate54inter7));
  inv1  gate1073(.a(G284), .O(gate54inter8));
  nand2 gate1074(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1075(.a(s_75), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1076(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1077(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1078(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1401(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1402(.a(gate55inter0), .b(s_122), .O(gate55inter1));
  and2  gate1403(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1404(.a(s_122), .O(gate55inter3));
  inv1  gate1405(.a(s_123), .O(gate55inter4));
  nand2 gate1406(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1407(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1408(.a(G15), .O(gate55inter7));
  inv1  gate1409(.a(G287), .O(gate55inter8));
  nand2 gate1410(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1411(.a(s_123), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1412(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1413(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1414(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1961(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1962(.a(gate59inter0), .b(s_202), .O(gate59inter1));
  and2  gate1963(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1964(.a(s_202), .O(gate59inter3));
  inv1  gate1965(.a(s_203), .O(gate59inter4));
  nand2 gate1966(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1967(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1968(.a(G19), .O(gate59inter7));
  inv1  gate1969(.a(G293), .O(gate59inter8));
  nand2 gate1970(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1971(.a(s_203), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1972(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1973(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1974(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate981(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate982(.a(gate61inter0), .b(s_62), .O(gate61inter1));
  and2  gate983(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate984(.a(s_62), .O(gate61inter3));
  inv1  gate985(.a(s_63), .O(gate61inter4));
  nand2 gate986(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate987(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate988(.a(G21), .O(gate61inter7));
  inv1  gate989(.a(G296), .O(gate61inter8));
  nand2 gate990(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate991(.a(s_63), .b(gate61inter3), .O(gate61inter10));
  nor2  gate992(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate993(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate994(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2213(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2214(.a(gate62inter0), .b(s_238), .O(gate62inter1));
  and2  gate2215(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2216(.a(s_238), .O(gate62inter3));
  inv1  gate2217(.a(s_239), .O(gate62inter4));
  nand2 gate2218(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2219(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2220(.a(G22), .O(gate62inter7));
  inv1  gate2221(.a(G296), .O(gate62inter8));
  nand2 gate2222(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2223(.a(s_239), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2224(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2225(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2226(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2115(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2116(.a(gate63inter0), .b(s_224), .O(gate63inter1));
  and2  gate2117(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2118(.a(s_224), .O(gate63inter3));
  inv1  gate2119(.a(s_225), .O(gate63inter4));
  nand2 gate2120(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2121(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2122(.a(G23), .O(gate63inter7));
  inv1  gate2123(.a(G299), .O(gate63inter8));
  nand2 gate2124(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2125(.a(s_225), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2126(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2127(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2128(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate687(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate688(.a(gate66inter0), .b(s_20), .O(gate66inter1));
  and2  gate689(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate690(.a(s_20), .O(gate66inter3));
  inv1  gate691(.a(s_21), .O(gate66inter4));
  nand2 gate692(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate693(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate694(.a(G26), .O(gate66inter7));
  inv1  gate695(.a(G302), .O(gate66inter8));
  nand2 gate696(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate697(.a(s_21), .b(gate66inter3), .O(gate66inter10));
  nor2  gate698(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate699(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate700(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate2549(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2550(.a(gate67inter0), .b(s_286), .O(gate67inter1));
  and2  gate2551(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2552(.a(s_286), .O(gate67inter3));
  inv1  gate2553(.a(s_287), .O(gate67inter4));
  nand2 gate2554(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2555(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2556(.a(G27), .O(gate67inter7));
  inv1  gate2557(.a(G305), .O(gate67inter8));
  nand2 gate2558(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2559(.a(s_287), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2560(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2561(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2562(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2255(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2256(.a(gate69inter0), .b(s_244), .O(gate69inter1));
  and2  gate2257(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2258(.a(s_244), .O(gate69inter3));
  inv1  gate2259(.a(s_245), .O(gate69inter4));
  nand2 gate2260(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2261(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2262(.a(G29), .O(gate69inter7));
  inv1  gate2263(.a(G308), .O(gate69inter8));
  nand2 gate2264(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2265(.a(s_245), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2266(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2267(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2268(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1891(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1892(.a(gate71inter0), .b(s_192), .O(gate71inter1));
  and2  gate1893(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1894(.a(s_192), .O(gate71inter3));
  inv1  gate1895(.a(s_193), .O(gate71inter4));
  nand2 gate1896(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1897(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1898(.a(G31), .O(gate71inter7));
  inv1  gate1899(.a(G311), .O(gate71inter8));
  nand2 gate1900(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1901(.a(s_193), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1902(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1903(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1904(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1807(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1808(.a(gate74inter0), .b(s_180), .O(gate74inter1));
  and2  gate1809(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1810(.a(s_180), .O(gate74inter3));
  inv1  gate1811(.a(s_181), .O(gate74inter4));
  nand2 gate1812(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1813(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1814(.a(G5), .O(gate74inter7));
  inv1  gate1815(.a(G314), .O(gate74inter8));
  nand2 gate1816(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1817(.a(s_181), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1818(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1819(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1820(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2535(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2536(.a(gate76inter0), .b(s_284), .O(gate76inter1));
  and2  gate2537(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2538(.a(s_284), .O(gate76inter3));
  inv1  gate2539(.a(s_285), .O(gate76inter4));
  nand2 gate2540(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2541(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2542(.a(G13), .O(gate76inter7));
  inv1  gate2543(.a(G317), .O(gate76inter8));
  nand2 gate2544(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2545(.a(s_285), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2546(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2547(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2548(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate729(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate730(.a(gate81inter0), .b(s_26), .O(gate81inter1));
  and2  gate731(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate732(.a(s_26), .O(gate81inter3));
  inv1  gate733(.a(s_27), .O(gate81inter4));
  nand2 gate734(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate735(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate736(.a(G3), .O(gate81inter7));
  inv1  gate737(.a(G326), .O(gate81inter8));
  nand2 gate738(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate739(.a(s_27), .b(gate81inter3), .O(gate81inter10));
  nor2  gate740(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate741(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate742(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate841(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate842(.a(gate83inter0), .b(s_42), .O(gate83inter1));
  and2  gate843(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate844(.a(s_42), .O(gate83inter3));
  inv1  gate845(.a(s_43), .O(gate83inter4));
  nand2 gate846(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate847(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate848(.a(G11), .O(gate83inter7));
  inv1  gate849(.a(G329), .O(gate83inter8));
  nand2 gate850(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate851(.a(s_43), .b(gate83inter3), .O(gate83inter10));
  nor2  gate852(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate853(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate854(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate715(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate716(.a(gate85inter0), .b(s_24), .O(gate85inter1));
  and2  gate717(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate718(.a(s_24), .O(gate85inter3));
  inv1  gate719(.a(s_25), .O(gate85inter4));
  nand2 gate720(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate721(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate722(.a(G4), .O(gate85inter7));
  inv1  gate723(.a(G332), .O(gate85inter8));
  nand2 gate724(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate725(.a(s_25), .b(gate85inter3), .O(gate85inter10));
  nor2  gate726(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate727(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate728(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1149(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1150(.a(gate86inter0), .b(s_86), .O(gate86inter1));
  and2  gate1151(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1152(.a(s_86), .O(gate86inter3));
  inv1  gate1153(.a(s_87), .O(gate86inter4));
  nand2 gate1154(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1155(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1156(.a(G8), .O(gate86inter7));
  inv1  gate1157(.a(G332), .O(gate86inter8));
  nand2 gate1158(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1159(.a(s_87), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1160(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1161(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1162(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate939(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate940(.a(gate91inter0), .b(s_56), .O(gate91inter1));
  and2  gate941(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate942(.a(s_56), .O(gate91inter3));
  inv1  gate943(.a(s_57), .O(gate91inter4));
  nand2 gate944(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate945(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate946(.a(G25), .O(gate91inter7));
  inv1  gate947(.a(G341), .O(gate91inter8));
  nand2 gate948(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate949(.a(s_57), .b(gate91inter3), .O(gate91inter10));
  nor2  gate950(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate951(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate952(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2171(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2172(.a(gate92inter0), .b(s_232), .O(gate92inter1));
  and2  gate2173(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2174(.a(s_232), .O(gate92inter3));
  inv1  gate2175(.a(s_233), .O(gate92inter4));
  nand2 gate2176(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2177(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2178(.a(G29), .O(gate92inter7));
  inv1  gate2179(.a(G341), .O(gate92inter8));
  nand2 gate2180(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2181(.a(s_233), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2182(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2183(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2184(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1191(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1192(.a(gate94inter0), .b(s_92), .O(gate94inter1));
  and2  gate1193(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1194(.a(s_92), .O(gate94inter3));
  inv1  gate1195(.a(s_93), .O(gate94inter4));
  nand2 gate1196(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1197(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1198(.a(G22), .O(gate94inter7));
  inv1  gate1199(.a(G344), .O(gate94inter8));
  nand2 gate1200(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1201(.a(s_93), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1202(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1203(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1204(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1121(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1122(.a(gate95inter0), .b(s_82), .O(gate95inter1));
  and2  gate1123(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1124(.a(s_82), .O(gate95inter3));
  inv1  gate1125(.a(s_83), .O(gate95inter4));
  nand2 gate1126(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1127(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1128(.a(G26), .O(gate95inter7));
  inv1  gate1129(.a(G347), .O(gate95inter8));
  nand2 gate1130(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1131(.a(s_83), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1132(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1133(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1134(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate995(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate996(.a(gate96inter0), .b(s_64), .O(gate96inter1));
  and2  gate997(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate998(.a(s_64), .O(gate96inter3));
  inv1  gate999(.a(s_65), .O(gate96inter4));
  nand2 gate1000(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1001(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1002(.a(G30), .O(gate96inter7));
  inv1  gate1003(.a(G347), .O(gate96inter8));
  nand2 gate1004(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1005(.a(s_65), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1006(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1007(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1008(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2325(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2326(.a(gate97inter0), .b(s_254), .O(gate97inter1));
  and2  gate2327(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2328(.a(s_254), .O(gate97inter3));
  inv1  gate2329(.a(s_255), .O(gate97inter4));
  nand2 gate2330(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2331(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2332(.a(G19), .O(gate97inter7));
  inv1  gate2333(.a(G350), .O(gate97inter8));
  nand2 gate2334(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2335(.a(s_255), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2336(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2337(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2338(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1051(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1052(.a(gate99inter0), .b(s_72), .O(gate99inter1));
  and2  gate1053(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1054(.a(s_72), .O(gate99inter3));
  inv1  gate1055(.a(s_73), .O(gate99inter4));
  nand2 gate1056(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1057(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1058(.a(G27), .O(gate99inter7));
  inv1  gate1059(.a(G353), .O(gate99inter8));
  nand2 gate1060(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1061(.a(s_73), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1062(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1063(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1064(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate645(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate646(.a(gate101inter0), .b(s_14), .O(gate101inter1));
  and2  gate647(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate648(.a(s_14), .O(gate101inter3));
  inv1  gate649(.a(s_15), .O(gate101inter4));
  nand2 gate650(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate651(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate652(.a(G20), .O(gate101inter7));
  inv1  gate653(.a(G356), .O(gate101inter8));
  nand2 gate654(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate655(.a(s_15), .b(gate101inter3), .O(gate101inter10));
  nor2  gate656(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate657(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate658(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate589(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate590(.a(gate104inter0), .b(s_6), .O(gate104inter1));
  and2  gate591(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate592(.a(s_6), .O(gate104inter3));
  inv1  gate593(.a(s_7), .O(gate104inter4));
  nand2 gate594(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate595(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate596(.a(G32), .O(gate104inter7));
  inv1  gate597(.a(G359), .O(gate104inter8));
  nand2 gate598(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate599(.a(s_7), .b(gate104inter3), .O(gate104inter10));
  nor2  gate600(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate601(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate602(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1625(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1626(.a(gate112inter0), .b(s_154), .O(gate112inter1));
  and2  gate1627(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1628(.a(s_154), .O(gate112inter3));
  inv1  gate1629(.a(s_155), .O(gate112inter4));
  nand2 gate1630(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1631(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1632(.a(G376), .O(gate112inter7));
  inv1  gate1633(.a(G377), .O(gate112inter8));
  nand2 gate1634(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1635(.a(s_155), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1636(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1637(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1638(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2101(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2102(.a(gate114inter0), .b(s_222), .O(gate114inter1));
  and2  gate2103(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2104(.a(s_222), .O(gate114inter3));
  inv1  gate2105(.a(s_223), .O(gate114inter4));
  nand2 gate2106(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2107(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2108(.a(G380), .O(gate114inter7));
  inv1  gate2109(.a(G381), .O(gate114inter8));
  nand2 gate2110(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2111(.a(s_223), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2112(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2113(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2114(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1303(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1304(.a(gate117inter0), .b(s_108), .O(gate117inter1));
  and2  gate1305(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1306(.a(s_108), .O(gate117inter3));
  inv1  gate1307(.a(s_109), .O(gate117inter4));
  nand2 gate1308(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1309(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1310(.a(G386), .O(gate117inter7));
  inv1  gate1311(.a(G387), .O(gate117inter8));
  nand2 gate1312(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1313(.a(s_109), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1314(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1315(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1316(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1317(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1318(.a(gate119inter0), .b(s_110), .O(gate119inter1));
  and2  gate1319(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1320(.a(s_110), .O(gate119inter3));
  inv1  gate1321(.a(s_111), .O(gate119inter4));
  nand2 gate1322(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1323(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1324(.a(G390), .O(gate119inter7));
  inv1  gate1325(.a(G391), .O(gate119inter8));
  nand2 gate1326(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1327(.a(s_111), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1328(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1329(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1330(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate2409(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2410(.a(gate120inter0), .b(s_266), .O(gate120inter1));
  and2  gate2411(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2412(.a(s_266), .O(gate120inter3));
  inv1  gate2413(.a(s_267), .O(gate120inter4));
  nand2 gate2414(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2415(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2416(.a(G392), .O(gate120inter7));
  inv1  gate2417(.a(G393), .O(gate120inter8));
  nand2 gate2418(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2419(.a(s_267), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2420(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2421(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2422(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1639(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1640(.a(gate121inter0), .b(s_156), .O(gate121inter1));
  and2  gate1641(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1642(.a(s_156), .O(gate121inter3));
  inv1  gate1643(.a(s_157), .O(gate121inter4));
  nand2 gate1644(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1645(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1646(.a(G394), .O(gate121inter7));
  inv1  gate1647(.a(G395), .O(gate121inter8));
  nand2 gate1648(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1649(.a(s_157), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1650(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1651(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1652(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2003(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2004(.a(gate122inter0), .b(s_208), .O(gate122inter1));
  and2  gate2005(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2006(.a(s_208), .O(gate122inter3));
  inv1  gate2007(.a(s_209), .O(gate122inter4));
  nand2 gate2008(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2009(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2010(.a(G396), .O(gate122inter7));
  inv1  gate2011(.a(G397), .O(gate122inter8));
  nand2 gate2012(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2013(.a(s_209), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2014(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2015(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2016(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1765(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1766(.a(gate123inter0), .b(s_174), .O(gate123inter1));
  and2  gate1767(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1768(.a(s_174), .O(gate123inter3));
  inv1  gate1769(.a(s_175), .O(gate123inter4));
  nand2 gate1770(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1771(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1772(.a(G398), .O(gate123inter7));
  inv1  gate1773(.a(G399), .O(gate123inter8));
  nand2 gate1774(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1775(.a(s_175), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1776(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1777(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1778(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1751(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1752(.a(gate127inter0), .b(s_172), .O(gate127inter1));
  and2  gate1753(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1754(.a(s_172), .O(gate127inter3));
  inv1  gate1755(.a(s_173), .O(gate127inter4));
  nand2 gate1756(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1757(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1758(.a(G406), .O(gate127inter7));
  inv1  gate1759(.a(G407), .O(gate127inter8));
  nand2 gate1760(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1761(.a(s_173), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1762(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1763(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1764(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate757(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate758(.a(gate133inter0), .b(s_30), .O(gate133inter1));
  and2  gate759(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate760(.a(s_30), .O(gate133inter3));
  inv1  gate761(.a(s_31), .O(gate133inter4));
  nand2 gate762(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate763(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate764(.a(G418), .O(gate133inter7));
  inv1  gate765(.a(G419), .O(gate133inter8));
  nand2 gate766(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate767(.a(s_31), .b(gate133inter3), .O(gate133inter10));
  nor2  gate768(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate769(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate770(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate2451(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2452(.a(gate134inter0), .b(s_272), .O(gate134inter1));
  and2  gate2453(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2454(.a(s_272), .O(gate134inter3));
  inv1  gate2455(.a(s_273), .O(gate134inter4));
  nand2 gate2456(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2457(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2458(.a(G420), .O(gate134inter7));
  inv1  gate2459(.a(G421), .O(gate134inter8));
  nand2 gate2460(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2461(.a(s_273), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2462(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2463(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2464(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2129(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2130(.a(gate137inter0), .b(s_226), .O(gate137inter1));
  and2  gate2131(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2132(.a(s_226), .O(gate137inter3));
  inv1  gate2133(.a(s_227), .O(gate137inter4));
  nand2 gate2134(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2135(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2136(.a(G426), .O(gate137inter7));
  inv1  gate2137(.a(G429), .O(gate137inter8));
  nand2 gate2138(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2139(.a(s_227), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2140(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2141(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2142(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2199(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2200(.a(gate139inter0), .b(s_236), .O(gate139inter1));
  and2  gate2201(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2202(.a(s_236), .O(gate139inter3));
  inv1  gate2203(.a(s_237), .O(gate139inter4));
  nand2 gate2204(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2205(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2206(.a(G438), .O(gate139inter7));
  inv1  gate2207(.a(G441), .O(gate139inter8));
  nand2 gate2208(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2209(.a(s_237), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2210(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2211(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2212(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1485(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1486(.a(gate140inter0), .b(s_134), .O(gate140inter1));
  and2  gate1487(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1488(.a(s_134), .O(gate140inter3));
  inv1  gate1489(.a(s_135), .O(gate140inter4));
  nand2 gate1490(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1491(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1492(.a(G444), .O(gate140inter7));
  inv1  gate1493(.a(G447), .O(gate140inter8));
  nand2 gate1494(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1495(.a(s_135), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1496(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1497(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1498(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate785(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate786(.a(gate143inter0), .b(s_34), .O(gate143inter1));
  and2  gate787(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate788(.a(s_34), .O(gate143inter3));
  inv1  gate789(.a(s_35), .O(gate143inter4));
  nand2 gate790(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate791(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate792(.a(G462), .O(gate143inter7));
  inv1  gate793(.a(G465), .O(gate143inter8));
  nand2 gate794(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate795(.a(s_35), .b(gate143inter3), .O(gate143inter10));
  nor2  gate796(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate797(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate798(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1709(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1710(.a(gate144inter0), .b(s_166), .O(gate144inter1));
  and2  gate1711(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1712(.a(s_166), .O(gate144inter3));
  inv1  gate1713(.a(s_167), .O(gate144inter4));
  nand2 gate1714(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1715(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1716(.a(G468), .O(gate144inter7));
  inv1  gate1717(.a(G471), .O(gate144inter8));
  nand2 gate1718(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1719(.a(s_167), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1720(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1721(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1722(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2227(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2228(.a(gate151inter0), .b(s_240), .O(gate151inter1));
  and2  gate2229(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2230(.a(s_240), .O(gate151inter3));
  inv1  gate2231(.a(s_241), .O(gate151inter4));
  nand2 gate2232(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2233(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2234(.a(G510), .O(gate151inter7));
  inv1  gate2235(.a(G513), .O(gate151inter8));
  nand2 gate2236(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2237(.a(s_241), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2238(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2239(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2240(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1233(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1234(.a(gate158inter0), .b(s_98), .O(gate158inter1));
  and2  gate1235(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1236(.a(s_98), .O(gate158inter3));
  inv1  gate1237(.a(s_99), .O(gate158inter4));
  nand2 gate1238(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1239(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1240(.a(G441), .O(gate158inter7));
  inv1  gate1241(.a(G528), .O(gate158inter8));
  nand2 gate1242(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1243(.a(s_99), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1244(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1245(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1246(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate673(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate674(.a(gate172inter0), .b(s_18), .O(gate172inter1));
  and2  gate675(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate676(.a(s_18), .O(gate172inter3));
  inv1  gate677(.a(s_19), .O(gate172inter4));
  nand2 gate678(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate679(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate680(.a(G483), .O(gate172inter7));
  inv1  gate681(.a(G549), .O(gate172inter8));
  nand2 gate682(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate683(.a(s_19), .b(gate172inter3), .O(gate172inter10));
  nor2  gate684(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate685(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate686(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate743(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate744(.a(gate175inter0), .b(s_28), .O(gate175inter1));
  and2  gate745(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate746(.a(s_28), .O(gate175inter3));
  inv1  gate747(.a(s_29), .O(gate175inter4));
  nand2 gate748(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate749(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate750(.a(G492), .O(gate175inter7));
  inv1  gate751(.a(G555), .O(gate175inter8));
  nand2 gate752(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate753(.a(s_29), .b(gate175inter3), .O(gate175inter10));
  nor2  gate754(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate755(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate756(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1695(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1696(.a(gate182inter0), .b(s_164), .O(gate182inter1));
  and2  gate1697(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1698(.a(s_164), .O(gate182inter3));
  inv1  gate1699(.a(s_165), .O(gate182inter4));
  nand2 gate1700(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1701(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1702(.a(G513), .O(gate182inter7));
  inv1  gate1703(.a(G564), .O(gate182inter8));
  nand2 gate1704(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1705(.a(s_165), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1706(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1707(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1708(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate967(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate968(.a(gate185inter0), .b(s_60), .O(gate185inter1));
  and2  gate969(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate970(.a(s_60), .O(gate185inter3));
  inv1  gate971(.a(s_61), .O(gate185inter4));
  nand2 gate972(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate973(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate974(.a(G570), .O(gate185inter7));
  inv1  gate975(.a(G571), .O(gate185inter8));
  nand2 gate976(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate977(.a(s_61), .b(gate185inter3), .O(gate185inter10));
  nor2  gate978(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate979(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate980(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1513(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1514(.a(gate188inter0), .b(s_138), .O(gate188inter1));
  and2  gate1515(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1516(.a(s_138), .O(gate188inter3));
  inv1  gate1517(.a(s_139), .O(gate188inter4));
  nand2 gate1518(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1519(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1520(.a(G576), .O(gate188inter7));
  inv1  gate1521(.a(G577), .O(gate188inter8));
  nand2 gate1522(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1523(.a(s_139), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1524(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1525(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1526(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2017(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2018(.a(gate190inter0), .b(s_210), .O(gate190inter1));
  and2  gate2019(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2020(.a(s_210), .O(gate190inter3));
  inv1  gate2021(.a(s_211), .O(gate190inter4));
  nand2 gate2022(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2023(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2024(.a(G580), .O(gate190inter7));
  inv1  gate2025(.a(G581), .O(gate190inter8));
  nand2 gate2026(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2027(.a(s_211), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2028(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2029(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2030(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1555(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1556(.a(gate193inter0), .b(s_144), .O(gate193inter1));
  and2  gate1557(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1558(.a(s_144), .O(gate193inter3));
  inv1  gate1559(.a(s_145), .O(gate193inter4));
  nand2 gate1560(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1561(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1562(.a(G586), .O(gate193inter7));
  inv1  gate1563(.a(G587), .O(gate193inter8));
  nand2 gate1564(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1565(.a(s_145), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1566(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1567(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1568(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1429(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1430(.a(gate197inter0), .b(s_126), .O(gate197inter1));
  and2  gate1431(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1432(.a(s_126), .O(gate197inter3));
  inv1  gate1433(.a(s_127), .O(gate197inter4));
  nand2 gate1434(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1435(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1436(.a(G594), .O(gate197inter7));
  inv1  gate1437(.a(G595), .O(gate197inter8));
  nand2 gate1438(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1439(.a(s_127), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1440(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1441(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1442(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1835(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1836(.a(gate199inter0), .b(s_184), .O(gate199inter1));
  and2  gate1837(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1838(.a(s_184), .O(gate199inter3));
  inv1  gate1839(.a(s_185), .O(gate199inter4));
  nand2 gate1840(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1841(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1842(.a(G598), .O(gate199inter7));
  inv1  gate1843(.a(G599), .O(gate199inter8));
  nand2 gate1844(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1845(.a(s_185), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1846(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1847(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1848(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2031(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2032(.a(gate201inter0), .b(s_212), .O(gate201inter1));
  and2  gate2033(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2034(.a(s_212), .O(gate201inter3));
  inv1  gate2035(.a(s_213), .O(gate201inter4));
  nand2 gate2036(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2037(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2038(.a(G602), .O(gate201inter7));
  inv1  gate2039(.a(G607), .O(gate201inter8));
  nand2 gate2040(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2041(.a(s_213), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2042(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2043(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2044(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1723(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1724(.a(gate203inter0), .b(s_168), .O(gate203inter1));
  and2  gate1725(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1726(.a(s_168), .O(gate203inter3));
  inv1  gate1727(.a(s_169), .O(gate203inter4));
  nand2 gate1728(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1729(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1730(.a(G602), .O(gate203inter7));
  inv1  gate1731(.a(G612), .O(gate203inter8));
  nand2 gate1732(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1733(.a(s_169), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1734(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1735(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1736(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1597(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1598(.a(gate206inter0), .b(s_150), .O(gate206inter1));
  and2  gate1599(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1600(.a(s_150), .O(gate206inter3));
  inv1  gate1601(.a(s_151), .O(gate206inter4));
  nand2 gate1602(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1603(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1604(.a(G632), .O(gate206inter7));
  inv1  gate1605(.a(G637), .O(gate206inter8));
  nand2 gate1606(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1607(.a(s_151), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1608(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1609(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1610(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate897(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate898(.a(gate207inter0), .b(s_50), .O(gate207inter1));
  and2  gate899(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate900(.a(s_50), .O(gate207inter3));
  inv1  gate901(.a(s_51), .O(gate207inter4));
  nand2 gate902(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate903(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate904(.a(G622), .O(gate207inter7));
  inv1  gate905(.a(G632), .O(gate207inter8));
  nand2 gate906(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate907(.a(s_51), .b(gate207inter3), .O(gate207inter10));
  nor2  gate908(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate909(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate910(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1527(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1528(.a(gate209inter0), .b(s_140), .O(gate209inter1));
  and2  gate1529(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1530(.a(s_140), .O(gate209inter3));
  inv1  gate1531(.a(s_141), .O(gate209inter4));
  nand2 gate1532(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1533(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1534(.a(G602), .O(gate209inter7));
  inv1  gate1535(.a(G666), .O(gate209inter8));
  nand2 gate1536(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1537(.a(s_141), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1538(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1539(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1540(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate953(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate954(.a(gate212inter0), .b(s_58), .O(gate212inter1));
  and2  gate955(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate956(.a(s_58), .O(gate212inter3));
  inv1  gate957(.a(s_59), .O(gate212inter4));
  nand2 gate958(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate959(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate960(.a(G617), .O(gate212inter7));
  inv1  gate961(.a(G669), .O(gate212inter8));
  nand2 gate962(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate963(.a(s_59), .b(gate212inter3), .O(gate212inter10));
  nor2  gate964(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate965(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate966(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1037(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1038(.a(gate214inter0), .b(s_70), .O(gate214inter1));
  and2  gate1039(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1040(.a(s_70), .O(gate214inter3));
  inv1  gate1041(.a(s_71), .O(gate214inter4));
  nand2 gate1042(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1043(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1044(.a(G612), .O(gate214inter7));
  inv1  gate1045(.a(G672), .O(gate214inter8));
  nand2 gate1046(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1047(.a(s_71), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1048(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1049(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1050(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2157(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2158(.a(gate216inter0), .b(s_230), .O(gate216inter1));
  and2  gate2159(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2160(.a(s_230), .O(gate216inter3));
  inv1  gate2161(.a(s_231), .O(gate216inter4));
  nand2 gate2162(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2163(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2164(.a(G617), .O(gate216inter7));
  inv1  gate2165(.a(G675), .O(gate216inter8));
  nand2 gate2166(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2167(.a(s_231), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2168(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2169(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2170(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1023(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1024(.a(gate217inter0), .b(s_68), .O(gate217inter1));
  and2  gate1025(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1026(.a(s_68), .O(gate217inter3));
  inv1  gate1027(.a(s_69), .O(gate217inter4));
  nand2 gate1028(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1029(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1030(.a(G622), .O(gate217inter7));
  inv1  gate1031(.a(G678), .O(gate217inter8));
  nand2 gate1032(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1033(.a(s_69), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1034(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1035(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1036(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1737(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1738(.a(gate219inter0), .b(s_170), .O(gate219inter1));
  and2  gate1739(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1740(.a(s_170), .O(gate219inter3));
  inv1  gate1741(.a(s_171), .O(gate219inter4));
  nand2 gate1742(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1743(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1744(.a(G632), .O(gate219inter7));
  inv1  gate1745(.a(G681), .O(gate219inter8));
  nand2 gate1746(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1747(.a(s_171), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1748(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1749(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1750(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1905(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1906(.a(gate223inter0), .b(s_194), .O(gate223inter1));
  and2  gate1907(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1908(.a(s_194), .O(gate223inter3));
  inv1  gate1909(.a(s_195), .O(gate223inter4));
  nand2 gate1910(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1911(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1912(.a(G627), .O(gate223inter7));
  inv1  gate1913(.a(G687), .O(gate223inter8));
  nand2 gate1914(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1915(.a(s_195), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1916(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1917(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1918(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate2297(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2298(.a(gate224inter0), .b(s_250), .O(gate224inter1));
  and2  gate2299(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2300(.a(s_250), .O(gate224inter3));
  inv1  gate2301(.a(s_251), .O(gate224inter4));
  nand2 gate2302(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2303(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2304(.a(G637), .O(gate224inter7));
  inv1  gate2305(.a(G687), .O(gate224inter8));
  nand2 gate2306(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2307(.a(s_251), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2308(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2309(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2310(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1989(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1990(.a(gate225inter0), .b(s_206), .O(gate225inter1));
  and2  gate1991(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1992(.a(s_206), .O(gate225inter3));
  inv1  gate1993(.a(s_207), .O(gate225inter4));
  nand2 gate1994(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1995(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1996(.a(G690), .O(gate225inter7));
  inv1  gate1997(.a(G691), .O(gate225inter8));
  nand2 gate1998(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1999(.a(s_207), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2000(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2001(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2002(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1415(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1416(.a(gate226inter0), .b(s_124), .O(gate226inter1));
  and2  gate1417(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1418(.a(s_124), .O(gate226inter3));
  inv1  gate1419(.a(s_125), .O(gate226inter4));
  nand2 gate1420(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1421(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1422(.a(G692), .O(gate226inter7));
  inv1  gate1423(.a(G693), .O(gate226inter8));
  nand2 gate1424(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1425(.a(s_125), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1426(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1427(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1428(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1079(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1080(.a(gate233inter0), .b(s_76), .O(gate233inter1));
  and2  gate1081(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1082(.a(s_76), .O(gate233inter3));
  inv1  gate1083(.a(s_77), .O(gate233inter4));
  nand2 gate1084(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1085(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1086(.a(G242), .O(gate233inter7));
  inv1  gate1087(.a(G718), .O(gate233inter8));
  nand2 gate1088(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1089(.a(s_77), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1090(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1091(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1092(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1387(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1388(.a(gate234inter0), .b(s_120), .O(gate234inter1));
  and2  gate1389(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1390(.a(s_120), .O(gate234inter3));
  inv1  gate1391(.a(s_121), .O(gate234inter4));
  nand2 gate1392(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1393(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1394(.a(G245), .O(gate234inter7));
  inv1  gate1395(.a(G721), .O(gate234inter8));
  nand2 gate1396(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1397(.a(s_121), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1398(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1399(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1400(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate603(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate604(.a(gate235inter0), .b(s_8), .O(gate235inter1));
  and2  gate605(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate606(.a(s_8), .O(gate235inter3));
  inv1  gate607(.a(s_9), .O(gate235inter4));
  nand2 gate608(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate609(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate610(.a(G248), .O(gate235inter7));
  inv1  gate611(.a(G724), .O(gate235inter8));
  nand2 gate612(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate613(.a(s_9), .b(gate235inter3), .O(gate235inter10));
  nor2  gate614(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate615(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate616(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate1163(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1164(.a(gate236inter0), .b(s_88), .O(gate236inter1));
  and2  gate1165(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1166(.a(s_88), .O(gate236inter3));
  inv1  gate1167(.a(s_89), .O(gate236inter4));
  nand2 gate1168(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1169(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1170(.a(G251), .O(gate236inter7));
  inv1  gate1171(.a(G727), .O(gate236inter8));
  nand2 gate1172(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1173(.a(s_89), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1174(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1175(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1176(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1779(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1780(.a(gate237inter0), .b(s_176), .O(gate237inter1));
  and2  gate1781(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1782(.a(s_176), .O(gate237inter3));
  inv1  gate1783(.a(s_177), .O(gate237inter4));
  nand2 gate1784(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1785(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1786(.a(G254), .O(gate237inter7));
  inv1  gate1787(.a(G706), .O(gate237inter8));
  nand2 gate1788(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1789(.a(s_177), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1790(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1791(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1792(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate883(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate884(.a(gate238inter0), .b(s_48), .O(gate238inter1));
  and2  gate885(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate886(.a(s_48), .O(gate238inter3));
  inv1  gate887(.a(s_49), .O(gate238inter4));
  nand2 gate888(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate889(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate890(.a(G257), .O(gate238inter7));
  inv1  gate891(.a(G709), .O(gate238inter8));
  nand2 gate892(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate893(.a(s_49), .b(gate238inter3), .O(gate238inter10));
  nor2  gate894(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate895(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate896(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2241(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2242(.a(gate244inter0), .b(s_242), .O(gate244inter1));
  and2  gate2243(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2244(.a(s_242), .O(gate244inter3));
  inv1  gate2245(.a(s_243), .O(gate244inter4));
  nand2 gate2246(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2247(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2248(.a(G721), .O(gate244inter7));
  inv1  gate2249(.a(G733), .O(gate244inter8));
  nand2 gate2250(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2251(.a(s_243), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2252(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2253(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2254(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2353(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2354(.a(gate249inter0), .b(s_258), .O(gate249inter1));
  and2  gate2355(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2356(.a(s_258), .O(gate249inter3));
  inv1  gate2357(.a(s_259), .O(gate249inter4));
  nand2 gate2358(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2359(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2360(.a(G254), .O(gate249inter7));
  inv1  gate2361(.a(G742), .O(gate249inter8));
  nand2 gate2362(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2363(.a(s_259), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2364(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2365(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2366(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2437(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2438(.a(gate254inter0), .b(s_270), .O(gate254inter1));
  and2  gate2439(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2440(.a(s_270), .O(gate254inter3));
  inv1  gate2441(.a(s_271), .O(gate254inter4));
  nand2 gate2442(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2443(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2444(.a(G712), .O(gate254inter7));
  inv1  gate2445(.a(G748), .O(gate254inter8));
  nand2 gate2446(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2447(.a(s_271), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2448(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2449(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2450(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate575(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate576(.a(gate256inter0), .b(s_4), .O(gate256inter1));
  and2  gate577(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate578(.a(s_4), .O(gate256inter3));
  inv1  gate579(.a(s_5), .O(gate256inter4));
  nand2 gate580(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate581(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate582(.a(G715), .O(gate256inter7));
  inv1  gate583(.a(G751), .O(gate256inter8));
  nand2 gate584(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate585(.a(s_5), .b(gate256inter3), .O(gate256inter10));
  nor2  gate586(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate587(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate588(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate869(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate870(.a(gate257inter0), .b(s_46), .O(gate257inter1));
  and2  gate871(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate872(.a(s_46), .O(gate257inter3));
  inv1  gate873(.a(s_47), .O(gate257inter4));
  nand2 gate874(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate875(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate876(.a(G754), .O(gate257inter7));
  inv1  gate877(.a(G755), .O(gate257inter8));
  nand2 gate878(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate879(.a(s_47), .b(gate257inter3), .O(gate257inter10));
  nor2  gate880(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate881(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate882(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate2185(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2186(.a(gate259inter0), .b(s_234), .O(gate259inter1));
  and2  gate2187(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2188(.a(s_234), .O(gate259inter3));
  inv1  gate2189(.a(s_235), .O(gate259inter4));
  nand2 gate2190(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2191(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2192(.a(G758), .O(gate259inter7));
  inv1  gate2193(.a(G759), .O(gate259inter8));
  nand2 gate2194(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2195(.a(s_235), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2196(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2197(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2198(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2143(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2144(.a(gate265inter0), .b(s_228), .O(gate265inter1));
  and2  gate2145(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2146(.a(s_228), .O(gate265inter3));
  inv1  gate2147(.a(s_229), .O(gate265inter4));
  nand2 gate2148(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2149(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2150(.a(G642), .O(gate265inter7));
  inv1  gate2151(.a(G770), .O(gate265inter8));
  nand2 gate2152(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2153(.a(s_229), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2154(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2155(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2156(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate631(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate632(.a(gate266inter0), .b(s_12), .O(gate266inter1));
  and2  gate633(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate634(.a(s_12), .O(gate266inter3));
  inv1  gate635(.a(s_13), .O(gate266inter4));
  nand2 gate636(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate637(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate638(.a(G645), .O(gate266inter7));
  inv1  gate639(.a(G773), .O(gate266inter8));
  nand2 gate640(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate641(.a(s_13), .b(gate266inter3), .O(gate266inter10));
  nor2  gate642(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate643(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate644(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate547(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate548(.a(gate268inter0), .b(s_0), .O(gate268inter1));
  and2  gate549(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate550(.a(s_0), .O(gate268inter3));
  inv1  gate551(.a(s_1), .O(gate268inter4));
  nand2 gate552(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate553(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate554(.a(G651), .O(gate268inter7));
  inv1  gate555(.a(G779), .O(gate268inter8));
  nand2 gate556(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate557(.a(s_1), .b(gate268inter3), .O(gate268inter10));
  nor2  gate558(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate559(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate560(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate701(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate702(.a(gate273inter0), .b(s_22), .O(gate273inter1));
  and2  gate703(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate704(.a(s_22), .O(gate273inter3));
  inv1  gate705(.a(s_23), .O(gate273inter4));
  nand2 gate706(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate707(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate708(.a(G642), .O(gate273inter7));
  inv1  gate709(.a(G794), .O(gate273inter8));
  nand2 gate710(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate711(.a(s_23), .b(gate273inter3), .O(gate273inter10));
  nor2  gate712(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate713(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate714(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1975(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1976(.a(gate277inter0), .b(s_204), .O(gate277inter1));
  and2  gate1977(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1978(.a(s_204), .O(gate277inter3));
  inv1  gate1979(.a(s_205), .O(gate277inter4));
  nand2 gate1980(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1981(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1982(.a(G648), .O(gate277inter7));
  inv1  gate1983(.a(G800), .O(gate277inter8));
  nand2 gate1984(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1985(.a(s_205), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1986(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1987(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1988(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1359(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1360(.a(gate283inter0), .b(s_116), .O(gate283inter1));
  and2  gate1361(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1362(.a(s_116), .O(gate283inter3));
  inv1  gate1363(.a(s_117), .O(gate283inter4));
  nand2 gate1364(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1365(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1366(.a(G657), .O(gate283inter7));
  inv1  gate1367(.a(G809), .O(gate283inter8));
  nand2 gate1368(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1369(.a(s_117), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1370(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1371(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1372(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1947(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1948(.a(gate284inter0), .b(s_200), .O(gate284inter1));
  and2  gate1949(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1950(.a(s_200), .O(gate284inter3));
  inv1  gate1951(.a(s_201), .O(gate284inter4));
  nand2 gate1952(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1953(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1954(.a(G785), .O(gate284inter7));
  inv1  gate1955(.a(G809), .O(gate284inter8));
  nand2 gate1956(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1957(.a(s_201), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1958(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1959(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1960(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2311(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2312(.a(gate290inter0), .b(s_252), .O(gate290inter1));
  and2  gate2313(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2314(.a(s_252), .O(gate290inter3));
  inv1  gate2315(.a(s_253), .O(gate290inter4));
  nand2 gate2316(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2317(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2318(.a(G820), .O(gate290inter7));
  inv1  gate2319(.a(G821), .O(gate290inter8));
  nand2 gate2320(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2321(.a(s_253), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2322(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2323(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2324(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1219(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1220(.a(gate292inter0), .b(s_96), .O(gate292inter1));
  and2  gate1221(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1222(.a(s_96), .O(gate292inter3));
  inv1  gate1223(.a(s_97), .O(gate292inter4));
  nand2 gate1224(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1225(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1226(.a(G824), .O(gate292inter7));
  inv1  gate1227(.a(G825), .O(gate292inter8));
  nand2 gate1228(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1229(.a(s_97), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1230(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1231(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1232(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate911(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate912(.a(gate296inter0), .b(s_52), .O(gate296inter1));
  and2  gate913(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate914(.a(s_52), .O(gate296inter3));
  inv1  gate915(.a(s_53), .O(gate296inter4));
  nand2 gate916(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate917(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate918(.a(G826), .O(gate296inter7));
  inv1  gate919(.a(G827), .O(gate296inter8));
  nand2 gate920(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate921(.a(s_53), .b(gate296inter3), .O(gate296inter10));
  nor2  gate922(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate923(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate924(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2367(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2368(.a(gate388inter0), .b(s_260), .O(gate388inter1));
  and2  gate2369(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2370(.a(s_260), .O(gate388inter3));
  inv1  gate2371(.a(s_261), .O(gate388inter4));
  nand2 gate2372(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2373(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2374(.a(G2), .O(gate388inter7));
  inv1  gate2375(.a(G1039), .O(gate388inter8));
  nand2 gate2376(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2377(.a(s_261), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2378(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2379(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2380(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1135(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1136(.a(gate392inter0), .b(s_84), .O(gate392inter1));
  and2  gate1137(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1138(.a(s_84), .O(gate392inter3));
  inv1  gate1139(.a(s_85), .O(gate392inter4));
  nand2 gate1140(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1141(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1142(.a(G6), .O(gate392inter7));
  inv1  gate1143(.a(G1051), .O(gate392inter8));
  nand2 gate1144(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1145(.a(s_85), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1146(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1147(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1148(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1247(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1248(.a(gate393inter0), .b(s_100), .O(gate393inter1));
  and2  gate1249(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1250(.a(s_100), .O(gate393inter3));
  inv1  gate1251(.a(s_101), .O(gate393inter4));
  nand2 gate1252(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1253(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1254(.a(G7), .O(gate393inter7));
  inv1  gate1255(.a(G1054), .O(gate393inter8));
  nand2 gate1256(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1257(.a(s_101), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1258(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1259(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1260(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1611(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1612(.a(gate396inter0), .b(s_152), .O(gate396inter1));
  and2  gate1613(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1614(.a(s_152), .O(gate396inter3));
  inv1  gate1615(.a(s_153), .O(gate396inter4));
  nand2 gate1616(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1617(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1618(.a(G10), .O(gate396inter7));
  inv1  gate1619(.a(G1063), .O(gate396inter8));
  nand2 gate1620(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1621(.a(s_153), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1622(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1623(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1624(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1009(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1010(.a(gate401inter0), .b(s_66), .O(gate401inter1));
  and2  gate1011(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1012(.a(s_66), .O(gate401inter3));
  inv1  gate1013(.a(s_67), .O(gate401inter4));
  nand2 gate1014(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1015(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1016(.a(G15), .O(gate401inter7));
  inv1  gate1017(.a(G1078), .O(gate401inter8));
  nand2 gate1018(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1019(.a(s_67), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1020(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1021(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1022(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate2577(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2578(.a(gate402inter0), .b(s_290), .O(gate402inter1));
  and2  gate2579(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2580(.a(s_290), .O(gate402inter3));
  inv1  gate2581(.a(s_291), .O(gate402inter4));
  nand2 gate2582(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2583(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2584(.a(G16), .O(gate402inter7));
  inv1  gate2585(.a(G1081), .O(gate402inter8));
  nand2 gate2586(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2587(.a(s_291), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2588(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2589(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2590(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1289(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1290(.a(gate407inter0), .b(s_106), .O(gate407inter1));
  and2  gate1291(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1292(.a(s_106), .O(gate407inter3));
  inv1  gate1293(.a(s_107), .O(gate407inter4));
  nand2 gate1294(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1295(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1296(.a(G21), .O(gate407inter7));
  inv1  gate1297(.a(G1096), .O(gate407inter8));
  nand2 gate1298(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1299(.a(s_107), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1300(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1301(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1302(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2269(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2270(.a(gate412inter0), .b(s_246), .O(gate412inter1));
  and2  gate2271(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2272(.a(s_246), .O(gate412inter3));
  inv1  gate2273(.a(s_247), .O(gate412inter4));
  nand2 gate2274(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2275(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2276(.a(G26), .O(gate412inter7));
  inv1  gate2277(.a(G1111), .O(gate412inter8));
  nand2 gate2278(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2279(.a(s_247), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2280(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2281(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2282(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate617(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate618(.a(gate418inter0), .b(s_10), .O(gate418inter1));
  and2  gate619(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate620(.a(s_10), .O(gate418inter3));
  inv1  gate621(.a(s_11), .O(gate418inter4));
  nand2 gate622(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate623(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate624(.a(G32), .O(gate418inter7));
  inv1  gate625(.a(G1129), .O(gate418inter8));
  nand2 gate626(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate627(.a(s_11), .b(gate418inter3), .O(gate418inter10));
  nor2  gate628(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate629(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate630(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1499(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1500(.a(gate421inter0), .b(s_136), .O(gate421inter1));
  and2  gate1501(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1502(.a(s_136), .O(gate421inter3));
  inv1  gate1503(.a(s_137), .O(gate421inter4));
  nand2 gate1504(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1505(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1506(.a(G2), .O(gate421inter7));
  inv1  gate1507(.a(G1135), .O(gate421inter8));
  nand2 gate1508(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1509(.a(s_137), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1510(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1511(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1512(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2059(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2060(.a(gate424inter0), .b(s_216), .O(gate424inter1));
  and2  gate2061(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2062(.a(s_216), .O(gate424inter3));
  inv1  gate2063(.a(s_217), .O(gate424inter4));
  nand2 gate2064(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2065(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2066(.a(G1042), .O(gate424inter7));
  inv1  gate2067(.a(G1138), .O(gate424inter8));
  nand2 gate2068(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2069(.a(s_217), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2070(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2071(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2072(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate813(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate814(.a(gate425inter0), .b(s_38), .O(gate425inter1));
  and2  gate815(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate816(.a(s_38), .O(gate425inter3));
  inv1  gate817(.a(s_39), .O(gate425inter4));
  nand2 gate818(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate819(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate820(.a(G4), .O(gate425inter7));
  inv1  gate821(.a(G1141), .O(gate425inter8));
  nand2 gate822(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate823(.a(s_39), .b(gate425inter3), .O(gate425inter10));
  nor2  gate824(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate825(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate826(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1667(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1668(.a(gate426inter0), .b(s_160), .O(gate426inter1));
  and2  gate1669(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1670(.a(s_160), .O(gate426inter3));
  inv1  gate1671(.a(s_161), .O(gate426inter4));
  nand2 gate1672(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1673(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1674(.a(G1045), .O(gate426inter7));
  inv1  gate1675(.a(G1141), .O(gate426inter8));
  nand2 gate1676(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1677(.a(s_161), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1678(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1679(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1680(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2087(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2088(.a(gate430inter0), .b(s_220), .O(gate430inter1));
  and2  gate2089(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2090(.a(s_220), .O(gate430inter3));
  inv1  gate2091(.a(s_221), .O(gate430inter4));
  nand2 gate2092(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2093(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2094(.a(G1051), .O(gate430inter7));
  inv1  gate2095(.a(G1147), .O(gate430inter8));
  nand2 gate2096(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2097(.a(s_221), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2098(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2099(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2100(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1205(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1206(.a(gate434inter0), .b(s_94), .O(gate434inter1));
  and2  gate1207(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1208(.a(s_94), .O(gate434inter3));
  inv1  gate1209(.a(s_95), .O(gate434inter4));
  nand2 gate1210(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1211(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1212(.a(G1057), .O(gate434inter7));
  inv1  gate1213(.a(G1153), .O(gate434inter8));
  nand2 gate1214(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1215(.a(s_95), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1216(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1217(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1218(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1345(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1346(.a(gate438inter0), .b(s_114), .O(gate438inter1));
  and2  gate1347(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1348(.a(s_114), .O(gate438inter3));
  inv1  gate1349(.a(s_115), .O(gate438inter4));
  nand2 gate1350(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1351(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1352(.a(G1063), .O(gate438inter7));
  inv1  gate1353(.a(G1159), .O(gate438inter8));
  nand2 gate1354(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1355(.a(s_115), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1356(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1357(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1358(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2045(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2046(.a(gate443inter0), .b(s_214), .O(gate443inter1));
  and2  gate2047(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2048(.a(s_214), .O(gate443inter3));
  inv1  gate2049(.a(s_215), .O(gate443inter4));
  nand2 gate2050(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2051(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2052(.a(G13), .O(gate443inter7));
  inv1  gate2053(.a(G1168), .O(gate443inter8));
  nand2 gate2054(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2055(.a(s_215), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2056(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2057(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2058(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1443(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1444(.a(gate446inter0), .b(s_128), .O(gate446inter1));
  and2  gate1445(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1446(.a(s_128), .O(gate446inter3));
  inv1  gate1447(.a(s_129), .O(gate446inter4));
  nand2 gate1448(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1449(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1450(.a(G1075), .O(gate446inter7));
  inv1  gate1451(.a(G1171), .O(gate446inter8));
  nand2 gate1452(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1453(.a(s_129), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1454(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1455(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1456(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1919(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1920(.a(gate447inter0), .b(s_196), .O(gate447inter1));
  and2  gate1921(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1922(.a(s_196), .O(gate447inter3));
  inv1  gate1923(.a(s_197), .O(gate447inter4));
  nand2 gate1924(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1925(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1926(.a(G15), .O(gate447inter7));
  inv1  gate1927(.a(G1174), .O(gate447inter8));
  nand2 gate1928(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1929(.a(s_197), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1930(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1931(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1932(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2563(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2564(.a(gate453inter0), .b(s_288), .O(gate453inter1));
  and2  gate2565(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2566(.a(s_288), .O(gate453inter3));
  inv1  gate2567(.a(s_289), .O(gate453inter4));
  nand2 gate2568(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2569(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2570(.a(G18), .O(gate453inter7));
  inv1  gate2571(.a(G1183), .O(gate453inter8));
  nand2 gate2572(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2573(.a(s_289), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2574(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2575(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2576(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2073(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2074(.a(gate456inter0), .b(s_218), .O(gate456inter1));
  and2  gate2075(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2076(.a(s_218), .O(gate456inter3));
  inv1  gate2077(.a(s_219), .O(gate456inter4));
  nand2 gate2078(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2079(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2080(.a(G1090), .O(gate456inter7));
  inv1  gate2081(.a(G1186), .O(gate456inter8));
  nand2 gate2082(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2083(.a(s_219), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2084(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2085(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2086(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate771(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate772(.a(gate461inter0), .b(s_32), .O(gate461inter1));
  and2  gate773(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate774(.a(s_32), .O(gate461inter3));
  inv1  gate775(.a(s_33), .O(gate461inter4));
  nand2 gate776(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate777(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate778(.a(G22), .O(gate461inter7));
  inv1  gate779(.a(G1195), .O(gate461inter8));
  nand2 gate780(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate781(.a(s_33), .b(gate461inter3), .O(gate461inter10));
  nor2  gate782(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate783(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate784(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2479(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2480(.a(gate467inter0), .b(s_276), .O(gate467inter1));
  and2  gate2481(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2482(.a(s_276), .O(gate467inter3));
  inv1  gate2483(.a(s_277), .O(gate467inter4));
  nand2 gate2484(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2485(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2486(.a(G25), .O(gate467inter7));
  inv1  gate2487(.a(G1204), .O(gate467inter8));
  nand2 gate2488(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2489(.a(s_277), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2490(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2491(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2492(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1653(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1654(.a(gate469inter0), .b(s_158), .O(gate469inter1));
  and2  gate1655(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1656(.a(s_158), .O(gate469inter3));
  inv1  gate1657(.a(s_159), .O(gate469inter4));
  nand2 gate1658(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1659(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1660(.a(G26), .O(gate469inter7));
  inv1  gate1661(.a(G1207), .O(gate469inter8));
  nand2 gate1662(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1663(.a(s_159), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1664(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1665(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1666(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2381(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2382(.a(gate470inter0), .b(s_262), .O(gate470inter1));
  and2  gate2383(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2384(.a(s_262), .O(gate470inter3));
  inv1  gate2385(.a(s_263), .O(gate470inter4));
  nand2 gate2386(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2387(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2388(.a(G1111), .O(gate470inter7));
  inv1  gate2389(.a(G1207), .O(gate470inter8));
  nand2 gate2390(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2391(.a(s_263), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2392(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2393(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2394(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1373(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1374(.a(gate472inter0), .b(s_118), .O(gate472inter1));
  and2  gate1375(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1376(.a(s_118), .O(gate472inter3));
  inv1  gate1377(.a(s_119), .O(gate472inter4));
  nand2 gate1378(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1379(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1380(.a(G1114), .O(gate472inter7));
  inv1  gate1381(.a(G1210), .O(gate472inter8));
  nand2 gate1382(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1383(.a(s_119), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1384(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1385(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1386(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1093(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1094(.a(gate477inter0), .b(s_78), .O(gate477inter1));
  and2  gate1095(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1096(.a(s_78), .O(gate477inter3));
  inv1  gate1097(.a(s_79), .O(gate477inter4));
  nand2 gate1098(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1099(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1100(.a(G30), .O(gate477inter7));
  inv1  gate1101(.a(G1219), .O(gate477inter8));
  nand2 gate1102(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1103(.a(s_79), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1104(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1105(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1106(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1681(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1682(.a(gate479inter0), .b(s_162), .O(gate479inter1));
  and2  gate1683(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1684(.a(s_162), .O(gate479inter3));
  inv1  gate1685(.a(s_163), .O(gate479inter4));
  nand2 gate1686(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1687(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1688(.a(G31), .O(gate479inter7));
  inv1  gate1689(.a(G1222), .O(gate479inter8));
  nand2 gate1690(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1691(.a(s_163), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1692(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1693(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1694(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1177(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1178(.a(gate485inter0), .b(s_90), .O(gate485inter1));
  and2  gate1179(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1180(.a(s_90), .O(gate485inter3));
  inv1  gate1181(.a(s_91), .O(gate485inter4));
  nand2 gate1182(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1183(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1184(.a(G1232), .O(gate485inter7));
  inv1  gate1185(.a(G1233), .O(gate485inter8));
  nand2 gate1186(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1187(.a(s_91), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1188(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1189(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1190(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate925(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate926(.a(gate487inter0), .b(s_54), .O(gate487inter1));
  and2  gate927(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate928(.a(s_54), .O(gate487inter3));
  inv1  gate929(.a(s_55), .O(gate487inter4));
  nand2 gate930(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate931(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate932(.a(G1236), .O(gate487inter7));
  inv1  gate933(.a(G1237), .O(gate487inter8));
  nand2 gate934(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate935(.a(s_55), .b(gate487inter3), .O(gate487inter10));
  nor2  gate936(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate937(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate938(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1471(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1472(.a(gate488inter0), .b(s_132), .O(gate488inter1));
  and2  gate1473(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1474(.a(s_132), .O(gate488inter3));
  inv1  gate1475(.a(s_133), .O(gate488inter4));
  nand2 gate1476(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1477(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1478(.a(G1238), .O(gate488inter7));
  inv1  gate1479(.a(G1239), .O(gate488inter8));
  nand2 gate1480(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1481(.a(s_133), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1482(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1483(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1484(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2521(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2522(.a(gate490inter0), .b(s_282), .O(gate490inter1));
  and2  gate2523(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2524(.a(s_282), .O(gate490inter3));
  inv1  gate2525(.a(s_283), .O(gate490inter4));
  nand2 gate2526(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2527(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2528(.a(G1242), .O(gate490inter7));
  inv1  gate2529(.a(G1243), .O(gate490inter8));
  nand2 gate2530(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2531(.a(s_283), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2532(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2533(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2534(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1107(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1108(.a(gate491inter0), .b(s_80), .O(gate491inter1));
  and2  gate1109(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1110(.a(s_80), .O(gate491inter3));
  inv1  gate1111(.a(s_81), .O(gate491inter4));
  nand2 gate1112(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1113(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1114(.a(G1244), .O(gate491inter7));
  inv1  gate1115(.a(G1245), .O(gate491inter8));
  nand2 gate1116(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1117(.a(s_81), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1118(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1119(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1120(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2283(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2284(.a(gate496inter0), .b(s_248), .O(gate496inter1));
  and2  gate2285(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2286(.a(s_248), .O(gate496inter3));
  inv1  gate2287(.a(s_249), .O(gate496inter4));
  nand2 gate2288(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2289(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2290(.a(G1254), .O(gate496inter7));
  inv1  gate2291(.a(G1255), .O(gate496inter8));
  nand2 gate2292(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2293(.a(s_249), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2294(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2295(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2296(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1541(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1542(.a(gate503inter0), .b(s_142), .O(gate503inter1));
  and2  gate1543(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1544(.a(s_142), .O(gate503inter3));
  inv1  gate1545(.a(s_143), .O(gate503inter4));
  nand2 gate1546(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1547(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1548(.a(G1268), .O(gate503inter7));
  inv1  gate1549(.a(G1269), .O(gate503inter8));
  nand2 gate1550(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1551(.a(s_143), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1552(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1553(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1554(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2465(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2466(.a(gate504inter0), .b(s_274), .O(gate504inter1));
  and2  gate2467(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2468(.a(s_274), .O(gate504inter3));
  inv1  gate2469(.a(s_275), .O(gate504inter4));
  nand2 gate2470(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2471(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2472(.a(G1270), .O(gate504inter7));
  inv1  gate2473(.a(G1271), .O(gate504inter8));
  nand2 gate2474(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2475(.a(s_275), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2476(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2477(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2478(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1849(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1850(.a(gate506inter0), .b(s_186), .O(gate506inter1));
  and2  gate1851(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1852(.a(s_186), .O(gate506inter3));
  inv1  gate1853(.a(s_187), .O(gate506inter4));
  nand2 gate1854(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1855(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1856(.a(G1274), .O(gate506inter7));
  inv1  gate1857(.a(G1275), .O(gate506inter8));
  nand2 gate1858(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1859(.a(s_187), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1860(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1861(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1862(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1793(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1794(.a(gate507inter0), .b(s_178), .O(gate507inter1));
  and2  gate1795(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1796(.a(s_178), .O(gate507inter3));
  inv1  gate1797(.a(s_179), .O(gate507inter4));
  nand2 gate1798(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1799(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1800(.a(G1276), .O(gate507inter7));
  inv1  gate1801(.a(G1277), .O(gate507inter8));
  nand2 gate1802(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1803(.a(s_179), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1804(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1805(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1806(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2395(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2396(.a(gate511inter0), .b(s_264), .O(gate511inter1));
  and2  gate2397(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2398(.a(s_264), .O(gate511inter3));
  inv1  gate2399(.a(s_265), .O(gate511inter4));
  nand2 gate2400(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2401(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2402(.a(G1284), .O(gate511inter7));
  inv1  gate2403(.a(G1285), .O(gate511inter8));
  nand2 gate2404(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2405(.a(s_265), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2406(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2407(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2408(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1331(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1332(.a(gate512inter0), .b(s_112), .O(gate512inter1));
  and2  gate1333(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1334(.a(s_112), .O(gate512inter3));
  inv1  gate1335(.a(s_113), .O(gate512inter4));
  nand2 gate1336(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1337(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1338(.a(G1286), .O(gate512inter7));
  inv1  gate1339(.a(G1287), .O(gate512inter8));
  nand2 gate1340(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1341(.a(s_113), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1342(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1343(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1344(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule