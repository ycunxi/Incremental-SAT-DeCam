module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate805(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate806(.a(gate19inter0), .b(s_92), .O(gate19inter1));
  and2  gate807(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate808(.a(s_92), .O(gate19inter3));
  inv1  gate809(.a(s_93), .O(gate19inter4));
  nand2 gate810(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate811(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate812(.a(N118), .O(gate19inter7));
  inv1  gate813(.a(N4), .O(gate19inter8));
  nand2 gate814(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate815(.a(s_93), .b(gate19inter3), .O(gate19inter10));
  nor2  gate816(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate817(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate818(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate917(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate918(.a(gate20inter0), .b(s_108), .O(gate20inter1));
  and2  gate919(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate920(.a(s_108), .O(gate20inter3));
  inv1  gate921(.a(s_109), .O(gate20inter4));
  nand2 gate922(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate923(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate924(.a(N8), .O(gate20inter7));
  inv1  gate925(.a(N119), .O(gate20inter8));
  nand2 gate926(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate927(.a(s_109), .b(gate20inter3), .O(gate20inter10));
  nor2  gate928(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate929(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate930(.a(gate20inter12), .b(gate20inter1), .O(N157));

  xor2  gate679(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate680(.a(gate21inter0), .b(s_74), .O(gate21inter1));
  and2  gate681(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate682(.a(s_74), .O(gate21inter3));
  inv1  gate683(.a(s_75), .O(gate21inter4));
  nand2 gate684(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate685(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate686(.a(N14), .O(gate21inter7));
  inv1  gate687(.a(N119), .O(gate21inter8));
  nand2 gate688(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate689(.a(s_75), .b(gate21inter3), .O(gate21inter10));
  nor2  gate690(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate691(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate692(.a(gate21inter12), .b(gate21inter1), .O(N158));
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate427(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate428(.a(gate23inter0), .b(s_38), .O(gate23inter1));
  and2  gate429(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate430(.a(s_38), .O(gate23inter3));
  inv1  gate431(.a(s_39), .O(gate23inter4));
  nand2 gate432(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate433(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate434(.a(N126), .O(gate23inter7));
  inv1  gate435(.a(N30), .O(gate23inter8));
  nand2 gate436(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate437(.a(s_39), .b(gate23inter3), .O(gate23inter10));
  nor2  gate438(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate439(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate440(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );

  xor2  gate455(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate456(.a(gate25inter0), .b(s_42), .O(gate25inter1));
  and2  gate457(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate458(.a(s_42), .O(gate25inter3));
  inv1  gate459(.a(s_43), .O(gate25inter4));
  nand2 gate460(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate461(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate462(.a(N134), .O(gate25inter7));
  inv1  gate463(.a(N56), .O(gate25inter8));
  nand2 gate464(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate465(.a(s_43), .b(gate25inter3), .O(gate25inter10));
  nor2  gate466(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate467(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate468(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate273(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate274(.a(gate29inter0), .b(s_16), .O(gate29inter1));
  and2  gate275(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate276(.a(s_16), .O(gate29inter3));
  inv1  gate277(.a(s_17), .O(gate29inter4));
  nand2 gate278(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate279(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate280(.a(N150), .O(gate29inter7));
  inv1  gate281(.a(N108), .O(gate29inter8));
  nand2 gate282(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate283(.a(s_17), .b(gate29inter3), .O(gate29inter10));
  nor2  gate284(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate285(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate286(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );

  xor2  gate707(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate708(.a(gate31inter0), .b(s_78), .O(gate31inter1));
  and2  gate709(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate710(.a(s_78), .O(gate31inter3));
  inv1  gate711(.a(s_79), .O(gate31inter4));
  nand2 gate712(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate713(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate714(.a(N27), .O(gate31inter7));
  inv1  gate715(.a(N123), .O(gate31inter8));
  nand2 gate716(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate717(.a(s_79), .b(gate31inter3), .O(gate31inter10));
  nor2  gate718(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate719(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate720(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate595(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate596(.a(gate34inter0), .b(s_62), .O(gate34inter1));
  and2  gate597(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate598(.a(s_62), .O(gate34inter3));
  inv1  gate599(.a(s_63), .O(gate34inter4));
  nand2 gate600(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate601(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate602(.a(N47), .O(gate34inter7));
  inv1  gate603(.a(N131), .O(gate34inter8));
  nand2 gate604(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate605(.a(s_63), .b(gate34inter3), .O(gate34inter10));
  nor2  gate606(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate607(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate608(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate567(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate568(.a(gate35inter0), .b(s_58), .O(gate35inter1));
  and2  gate569(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate570(.a(s_58), .O(gate35inter3));
  inv1  gate571(.a(s_59), .O(gate35inter4));
  nand2 gate572(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate573(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate574(.a(N53), .O(gate35inter7));
  inv1  gate575(.a(N131), .O(gate35inter8));
  nand2 gate576(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate577(.a(s_59), .b(gate35inter3), .O(gate35inter10));
  nor2  gate578(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate579(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate580(.a(gate35inter12), .b(gate35inter1), .O(N188));

  xor2  gate525(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate526(.a(gate36inter0), .b(s_52), .O(gate36inter1));
  and2  gate527(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate528(.a(s_52), .O(gate36inter3));
  inv1  gate529(.a(s_53), .O(gate36inter4));
  nand2 gate530(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate531(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate532(.a(N60), .O(gate36inter7));
  inv1  gate533(.a(N135), .O(gate36inter8));
  nand2 gate534(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate535(.a(s_53), .b(gate36inter3), .O(gate36inter10));
  nor2  gate536(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate537(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate538(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate161(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate162(.a(gate38inter0), .b(s_0), .O(gate38inter1));
  and2  gate163(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate164(.a(s_0), .O(gate38inter3));
  inv1  gate165(.a(s_1), .O(gate38inter4));
  nand2 gate166(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate167(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate168(.a(N73), .O(gate38inter7));
  inv1  gate169(.a(N139), .O(gate38inter8));
  nand2 gate170(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate171(.a(s_1), .b(gate38inter3), .O(gate38inter10));
  nor2  gate172(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate173(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate174(.a(gate38inter12), .b(gate38inter1), .O(N191));
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate441(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate442(.a(gate40inter0), .b(s_40), .O(gate40inter1));
  and2  gate443(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate444(.a(s_40), .O(gate40inter3));
  inv1  gate445(.a(s_41), .O(gate40inter4));
  nand2 gate446(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate447(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate448(.a(N86), .O(gate40inter7));
  inv1  gate449(.a(N143), .O(gate40inter8));
  nand2 gate450(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate451(.a(s_41), .b(gate40inter3), .O(gate40inter10));
  nor2  gate452(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate453(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate454(.a(gate40inter12), .b(gate40inter1), .O(N193));

  xor2  gate189(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate190(.a(gate41inter0), .b(s_4), .O(gate41inter1));
  and2  gate191(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate192(.a(s_4), .O(gate41inter3));
  inv1  gate193(.a(s_5), .O(gate41inter4));
  nand2 gate194(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate195(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate196(.a(N92), .O(gate41inter7));
  inv1  gate197(.a(N143), .O(gate41inter8));
  nand2 gate198(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate199(.a(s_5), .b(gate41inter3), .O(gate41inter10));
  nor2  gate200(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate201(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate202(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate469(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate470(.a(gate43inter0), .b(s_44), .O(gate43inter1));
  and2  gate471(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate472(.a(s_44), .O(gate43inter3));
  inv1  gate473(.a(s_45), .O(gate43inter4));
  nand2 gate474(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate475(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate476(.a(N105), .O(gate43inter7));
  inv1  gate477(.a(N147), .O(gate43inter8));
  nand2 gate478(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate479(.a(s_45), .b(gate43inter3), .O(gate43inter10));
  nor2  gate480(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate481(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate482(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );

  xor2  gate791(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate792(.a(gate45inter0), .b(s_90), .O(gate45inter1));
  and2  gate793(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate794(.a(s_90), .O(gate45inter3));
  inv1  gate795(.a(s_91), .O(gate45inter4));
  nand2 gate796(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate797(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate798(.a(N115), .O(gate45inter7));
  inv1  gate799(.a(N151), .O(gate45inter8));
  nand2 gate800(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate801(.a(s_91), .b(gate45inter3), .O(gate45inter10));
  nor2  gate802(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate803(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate804(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate301(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate302(.a(gate50inter0), .b(s_20), .O(gate50inter1));
  and2  gate303(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate304(.a(s_20), .O(gate50inter3));
  inv1  gate305(.a(s_21), .O(gate50inter4));
  nand2 gate306(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate307(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate308(.a(N203), .O(gate50inter7));
  inv1  gate309(.a(N154), .O(gate50inter8));
  nand2 gate310(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate311(.a(s_21), .b(gate50inter3), .O(gate50inter10));
  nor2  gate312(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate313(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate314(.a(gate50inter12), .b(gate50inter1), .O(N224));
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate903(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate904(.a(gate52inter0), .b(s_106), .O(gate52inter1));
  and2  gate905(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate906(.a(s_106), .O(gate52inter3));
  inv1  gate907(.a(s_107), .O(gate52inter4));
  nand2 gate908(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate909(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate910(.a(N203), .O(gate52inter7));
  inv1  gate911(.a(N162), .O(gate52inter8));
  nand2 gate912(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate913(.a(s_107), .b(gate52inter3), .O(gate52inter10));
  nor2  gate914(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate915(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate916(.a(gate52inter12), .b(gate52inter1), .O(N230));

  xor2  gate329(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate330(.a(gate53inter0), .b(s_24), .O(gate53inter1));
  and2  gate331(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate332(.a(s_24), .O(gate53inter3));
  inv1  gate333(.a(s_25), .O(gate53inter4));
  nand2 gate334(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate335(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate336(.a(N203), .O(gate53inter7));
  inv1  gate337(.a(N165), .O(gate53inter8));
  nand2 gate338(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate339(.a(s_25), .b(gate53inter3), .O(gate53inter10));
  nor2  gate340(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate341(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate342(.a(gate53inter12), .b(gate53inter1), .O(N233));
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate665(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate666(.a(gate60inter0), .b(s_72), .O(gate60inter1));
  and2  gate667(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate668(.a(s_72), .O(gate60inter3));
  inv1  gate669(.a(s_73), .O(gate60inter4));
  nand2 gate670(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate671(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate672(.a(N213), .O(gate60inter7));
  inv1  gate673(.a(N24), .O(gate60inter8));
  nand2 gate674(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate675(.a(s_73), .b(gate60inter3), .O(gate60inter10));
  nor2  gate676(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate677(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate678(.a(gate60inter12), .b(gate60inter1), .O(N250));

  xor2  gate217(.a(N180), .b(N203), .O(gate61inter0));
  nand2 gate218(.a(gate61inter0), .b(s_8), .O(gate61inter1));
  and2  gate219(.a(N180), .b(N203), .O(gate61inter2));
  inv1  gate220(.a(s_8), .O(gate61inter3));
  inv1  gate221(.a(s_9), .O(gate61inter4));
  nand2 gate222(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate223(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate224(.a(N203), .O(gate61inter7));
  inv1  gate225(.a(N180), .O(gate61inter8));
  nand2 gate226(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate227(.a(s_9), .b(gate61inter3), .O(gate61inter10));
  nor2  gate228(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate229(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate230(.a(gate61inter12), .b(gate61inter1), .O(N251));
nand2 gate62( .a(N213), .b(N37), .O(N254) );

  xor2  gate847(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate848(.a(gate63inter0), .b(s_98), .O(gate63inter1));
  and2  gate849(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate850(.a(s_98), .O(gate63inter3));
  inv1  gate851(.a(s_99), .O(gate63inter4));
  nand2 gate852(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate853(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate854(.a(N213), .O(gate63inter7));
  inv1  gate855(.a(N50), .O(gate63inter8));
  nand2 gate856(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate857(.a(s_99), .b(gate63inter3), .O(gate63inter10));
  nor2  gate858(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate859(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate860(.a(gate63inter12), .b(gate63inter1), .O(N255));

  xor2  gate833(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate834(.a(gate64inter0), .b(s_96), .O(gate64inter1));
  and2  gate835(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate836(.a(s_96), .O(gate64inter3));
  inv1  gate837(.a(s_97), .O(gate64inter4));
  nand2 gate838(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate839(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate840(.a(N213), .O(gate64inter7));
  inv1  gate841(.a(N63), .O(gate64inter8));
  nand2 gate842(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate843(.a(s_97), .b(gate64inter3), .O(gate64inter10));
  nor2  gate844(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate845(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate846(.a(gate64inter12), .b(gate64inter1), .O(N256));

  xor2  gate511(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate512(.a(gate65inter0), .b(s_50), .O(gate65inter1));
  and2  gate513(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate514(.a(s_50), .O(gate65inter3));
  inv1  gate515(.a(s_51), .O(gate65inter4));
  nand2 gate516(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate517(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate518(.a(N213), .O(gate65inter7));
  inv1  gate519(.a(N76), .O(gate65inter8));
  nand2 gate520(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate521(.a(s_51), .b(gate65inter3), .O(gate65inter10));
  nor2  gate522(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate523(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate524(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate315(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate316(.a(gate68inter0), .b(s_22), .O(gate68inter1));
  and2  gate317(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate318(.a(s_22), .O(gate68inter3));
  inv1  gate319(.a(s_23), .O(gate68inter4));
  nand2 gate320(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate321(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate322(.a(N224), .O(gate68inter7));
  inv1  gate323(.a(N157), .O(gate68inter8));
  nand2 gate324(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate325(.a(s_23), .b(gate68inter3), .O(gate68inter10));
  nor2  gate326(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate327(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate328(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate399(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate400(.a(gate71inter0), .b(s_34), .O(gate71inter1));
  and2  gate401(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate402(.a(s_34), .O(gate71inter3));
  inv1  gate403(.a(s_35), .O(gate71inter4));
  nand2 gate404(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate405(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate406(.a(N230), .O(gate71inter7));
  inv1  gate407(.a(N185), .O(gate71inter8));
  nand2 gate408(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate409(.a(s_35), .b(gate71inter3), .O(gate71inter10));
  nor2  gate410(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate411(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate412(.a(gate71inter12), .b(gate71inter1), .O(N267));

  xor2  gate483(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate484(.a(gate72inter0), .b(s_46), .O(gate72inter1));
  and2  gate485(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate486(.a(s_46), .O(gate72inter3));
  inv1  gate487(.a(s_47), .O(gate72inter4));
  nand2 gate488(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate489(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate490(.a(N233), .O(gate72inter7));
  inv1  gate491(.a(N187), .O(gate72inter8));
  nand2 gate492(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate493(.a(s_47), .b(gate72inter3), .O(gate72inter10));
  nor2  gate494(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate495(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate496(.a(gate72inter12), .b(gate72inter1), .O(N270));

  xor2  gate693(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate694(.a(gate73inter0), .b(s_76), .O(gate73inter1));
  and2  gate695(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate696(.a(s_76), .O(gate73inter3));
  inv1  gate697(.a(s_77), .O(gate73inter4));
  nand2 gate698(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate699(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate700(.a(N236), .O(gate73inter7));
  inv1  gate701(.a(N189), .O(gate73inter8));
  nand2 gate702(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate703(.a(s_77), .b(gate73inter3), .O(gate73inter10));
  nor2  gate704(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate705(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate706(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate581(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate582(.a(gate75inter0), .b(s_60), .O(gate75inter1));
  and2  gate583(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate584(.a(s_60), .O(gate75inter3));
  inv1  gate585(.a(s_61), .O(gate75inter4));
  nand2 gate586(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate587(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate588(.a(N243), .O(gate75inter7));
  inv1  gate589(.a(N193), .O(gate75inter8));
  nand2 gate590(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate591(.a(s_61), .b(gate75inter3), .O(gate75inter10));
  nor2  gate592(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate593(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate594(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate539(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate540(.a(gate83inter0), .b(s_54), .O(gate83inter1));
  and2  gate541(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate542(.a(s_54), .O(gate83inter3));
  inv1  gate543(.a(s_55), .O(gate83inter4));
  nand2 gate544(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate545(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate546(.a(N243), .O(gate83inter7));
  inv1  gate547(.a(N194), .O(gate83inter8));
  nand2 gate548(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate549(.a(s_55), .b(gate83inter3), .O(gate83inter10));
  nor2  gate550(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate551(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate552(.a(gate83inter12), .b(gate83inter1), .O(N293));

  xor2  gate413(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate414(.a(gate84inter0), .b(s_36), .O(gate84inter1));
  and2  gate415(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate416(.a(s_36), .O(gate84inter3));
  inv1  gate417(.a(s_37), .O(gate84inter4));
  nand2 gate418(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate419(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate420(.a(N247), .O(gate84inter7));
  inv1  gate421(.a(N196), .O(gate84inter8));
  nand2 gate422(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate423(.a(s_37), .b(gate84inter3), .O(gate84inter10));
  nor2  gate424(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate425(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate426(.a(gate84inter12), .b(gate84inter1), .O(N294));

  xor2  gate357(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate358(.a(gate85inter0), .b(s_28), .O(gate85inter1));
  and2  gate359(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate360(.a(s_28), .O(gate85inter3));
  inv1  gate361(.a(s_29), .O(gate85inter4));
  nand2 gate362(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate363(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate364(.a(N251), .O(gate85inter7));
  inv1  gate365(.a(N198), .O(gate85inter8));
  nand2 gate366(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate367(.a(s_29), .b(gate85inter3), .O(gate85inter10));
  nor2  gate368(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate369(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate370(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate385(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate386(.a(gate99inter0), .b(s_32), .O(gate99inter1));
  and2  gate387(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate388(.a(s_32), .O(gate99inter3));
  inv1  gate389(.a(s_33), .O(gate99inter4));
  nand2 gate390(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate391(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate392(.a(N309), .O(gate99inter7));
  inv1  gate393(.a(N260), .O(gate99inter8));
  nand2 gate394(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate395(.a(s_33), .b(gate99inter3), .O(gate99inter10));
  nor2  gate396(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate397(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate398(.a(gate99inter12), .b(gate99inter1), .O(N330));

  xor2  gate861(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate862(.a(gate100inter0), .b(s_100), .O(gate100inter1));
  and2  gate863(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate864(.a(s_100), .O(gate100inter3));
  inv1  gate865(.a(s_101), .O(gate100inter4));
  nand2 gate866(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate867(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate868(.a(N309), .O(gate100inter7));
  inv1  gate869(.a(N264), .O(gate100inter8));
  nand2 gate870(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate871(.a(s_101), .b(gate100inter3), .O(gate100inter10));
  nor2  gate872(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate873(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate874(.a(gate100inter12), .b(gate100inter1), .O(N331));

  xor2  gate875(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate876(.a(gate101inter0), .b(s_102), .O(gate101inter1));
  and2  gate877(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate878(.a(s_102), .O(gate101inter3));
  inv1  gate879(.a(s_103), .O(gate101inter4));
  nand2 gate880(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate881(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate882(.a(N309), .O(gate101inter7));
  inv1  gate883(.a(N267), .O(gate101inter8));
  nand2 gate884(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate885(.a(s_103), .b(gate101inter3), .O(gate101inter10));
  nor2  gate886(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate887(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate888(.a(gate101inter12), .b(gate101inter1), .O(N332));

  xor2  gate637(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate638(.a(gate102inter0), .b(s_68), .O(gate102inter1));
  and2  gate639(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate640(.a(s_68), .O(gate102inter3));
  inv1  gate641(.a(s_69), .O(gate102inter4));
  nand2 gate642(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate643(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate644(.a(N309), .O(gate102inter7));
  inv1  gate645(.a(N270), .O(gate102inter8));
  nand2 gate646(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate647(.a(s_69), .b(gate102inter3), .O(gate102inter10));
  nor2  gate648(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate649(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate650(.a(gate102inter12), .b(gate102inter1), .O(N333));

  xor2  gate763(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate764(.a(gate103inter0), .b(s_86), .O(gate103inter1));
  and2  gate765(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate766(.a(s_86), .O(gate103inter3));
  inv1  gate767(.a(s_87), .O(gate103inter4));
  nand2 gate768(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate769(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate770(.a(N8), .O(gate103inter7));
  inv1  gate771(.a(N319), .O(gate103inter8));
  nand2 gate772(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate773(.a(s_87), .b(gate103inter3), .O(gate103inter10));
  nor2  gate774(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate775(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate776(.a(gate103inter12), .b(gate103inter1), .O(N334));

  xor2  gate889(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate890(.a(gate104inter0), .b(s_104), .O(gate104inter1));
  and2  gate891(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate892(.a(s_104), .O(gate104inter3));
  inv1  gate893(.a(s_105), .O(gate104inter4));
  nand2 gate894(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate895(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate896(.a(N309), .O(gate104inter7));
  inv1  gate897(.a(N273), .O(gate104inter8));
  nand2 gate898(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate899(.a(s_105), .b(gate104inter3), .O(gate104inter10));
  nor2  gate900(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate901(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate902(.a(gate104inter12), .b(gate104inter1), .O(N335));

  xor2  gate735(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate736(.a(gate105inter0), .b(s_82), .O(gate105inter1));
  and2  gate737(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate738(.a(s_82), .O(gate105inter3));
  inv1  gate739(.a(s_83), .O(gate105inter4));
  nand2 gate740(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate741(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate742(.a(N319), .O(gate105inter7));
  inv1  gate743(.a(N21), .O(gate105inter8));
  nand2 gate744(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate745(.a(s_83), .b(gate105inter3), .O(gate105inter10));
  nor2  gate746(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate747(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate748(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );

  xor2  gate343(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate344(.a(gate107inter0), .b(s_26), .O(gate107inter1));
  and2  gate345(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate346(.a(s_26), .O(gate107inter3));
  inv1  gate347(.a(s_27), .O(gate107inter4));
  nand2 gate348(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate349(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate350(.a(N319), .O(gate107inter7));
  inv1  gate351(.a(N34), .O(gate107inter8));
  nand2 gate352(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate353(.a(s_27), .b(gate107inter3), .O(gate107inter10));
  nor2  gate354(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate355(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate356(.a(gate107inter12), .b(gate107inter1), .O(N338));

  xor2  gate497(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate498(.a(gate108inter0), .b(s_48), .O(gate108inter1));
  and2  gate499(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate500(.a(s_48), .O(gate108inter3));
  inv1  gate501(.a(s_49), .O(gate108inter4));
  nand2 gate502(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate503(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate504(.a(N309), .O(gate108inter7));
  inv1  gate505(.a(N279), .O(gate108inter8));
  nand2 gate506(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate507(.a(s_49), .b(gate108inter3), .O(gate108inter10));
  nor2  gate508(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate509(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate510(.a(gate108inter12), .b(gate108inter1), .O(N339));

  xor2  gate819(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate820(.a(gate109inter0), .b(s_94), .O(gate109inter1));
  and2  gate821(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate822(.a(s_94), .O(gate109inter3));
  inv1  gate823(.a(s_95), .O(gate109inter4));
  nand2 gate824(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate825(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate826(.a(N319), .O(gate109inter7));
  inv1  gate827(.a(N47), .O(gate109inter8));
  nand2 gate828(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate829(.a(s_95), .b(gate109inter3), .O(gate109inter10));
  nor2  gate830(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate831(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate832(.a(gate109inter12), .b(gate109inter1), .O(N340));
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate553(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate554(.a(gate111inter0), .b(s_56), .O(gate111inter1));
  and2  gate555(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate556(.a(s_56), .O(gate111inter3));
  inv1  gate557(.a(s_57), .O(gate111inter4));
  nand2 gate558(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate559(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate560(.a(N319), .O(gate111inter7));
  inv1  gate561(.a(N60), .O(gate111inter8));
  nand2 gate562(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate563(.a(s_57), .b(gate111inter3), .O(gate111inter10));
  nor2  gate564(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate565(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate566(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate721(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate722(.a(gate113inter0), .b(s_80), .O(gate113inter1));
  and2  gate723(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate724(.a(s_80), .O(gate113inter3));
  inv1  gate725(.a(s_81), .O(gate113inter4));
  nand2 gate726(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate727(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate728(.a(N319), .O(gate113inter7));
  inv1  gate729(.a(N73), .O(gate113inter8));
  nand2 gate730(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate731(.a(s_81), .b(gate113inter3), .O(gate113inter10));
  nor2  gate732(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate733(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate734(.a(gate113inter12), .b(gate113inter1), .O(N344));

  xor2  gate203(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate204(.a(gate114inter0), .b(s_6), .O(gate114inter1));
  and2  gate205(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate206(.a(s_6), .O(gate114inter3));
  inv1  gate207(.a(s_7), .O(gate114inter4));
  nand2 gate208(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate209(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate210(.a(N319), .O(gate114inter7));
  inv1  gate211(.a(N86), .O(gate114inter8));
  nand2 gate212(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate213(.a(s_7), .b(gate114inter3), .O(gate114inter10));
  nor2  gate214(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate215(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate216(.a(gate114inter12), .b(gate114inter1), .O(N345));

  xor2  gate259(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate260(.a(gate115inter0), .b(s_14), .O(gate115inter1));
  and2  gate261(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate262(.a(s_14), .O(gate115inter3));
  inv1  gate263(.a(s_15), .O(gate115inter4));
  nand2 gate264(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate265(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate266(.a(N319), .O(gate115inter7));
  inv1  gate267(.a(N99), .O(gate115inter8));
  nand2 gate268(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate269(.a(s_15), .b(gate115inter3), .O(gate115inter10));
  nor2  gate270(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate271(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate272(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );

  xor2  gate623(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate624(.a(gate117inter0), .b(s_66), .O(gate117inter1));
  and2  gate625(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate626(.a(s_66), .O(gate117inter3));
  inv1  gate627(.a(s_67), .O(gate117inter4));
  nand2 gate628(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate629(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate630(.a(N330), .O(gate117inter7));
  inv1  gate631(.a(N300), .O(gate117inter8));
  nand2 gate632(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate633(.a(s_67), .b(gate117inter3), .O(gate117inter10));
  nor2  gate634(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate635(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate636(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate651(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate652(.a(gate119inter0), .b(s_70), .O(gate119inter1));
  and2  gate653(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate654(.a(s_70), .O(gate119inter3));
  inv1  gate655(.a(s_71), .O(gate119inter4));
  nand2 gate656(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate657(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate658(.a(N332), .O(gate119inter7));
  inv1  gate659(.a(N302), .O(gate119inter8));
  nand2 gate660(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate661(.a(s_71), .b(gate119inter3), .O(gate119inter10));
  nor2  gate662(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate663(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate664(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate371(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate372(.a(gate121inter0), .b(s_30), .O(gate121inter1));
  and2  gate373(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate374(.a(s_30), .O(gate121inter3));
  inv1  gate375(.a(s_31), .O(gate121inter4));
  nand2 gate376(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate377(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate378(.a(N335), .O(gate121inter7));
  inv1  gate379(.a(N304), .O(gate121inter8));
  nand2 gate380(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate381(.a(s_31), .b(gate121inter3), .O(gate121inter10));
  nor2  gate382(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate383(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate384(.a(gate121inter12), .b(gate121inter1), .O(N352));

  xor2  gate931(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate932(.a(gate122inter0), .b(s_110), .O(gate122inter1));
  and2  gate933(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate934(.a(s_110), .O(gate122inter3));
  inv1  gate935(.a(s_111), .O(gate122inter4));
  nand2 gate936(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate937(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate938(.a(N337), .O(gate122inter7));
  inv1  gate939(.a(N305), .O(gate122inter8));
  nand2 gate940(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate941(.a(s_111), .b(gate122inter3), .O(gate122inter10));
  nor2  gate942(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate943(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate944(.a(gate122inter12), .b(gate122inter1), .O(N353));
nand2 gate123( .a(N339), .b(N306), .O(N354) );

  xor2  gate749(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate750(.a(gate124inter0), .b(s_84), .O(gate124inter1));
  and2  gate751(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate752(.a(s_84), .O(gate124inter3));
  inv1  gate753(.a(s_85), .O(gate124inter4));
  nand2 gate754(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate755(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate756(.a(N341), .O(gate124inter7));
  inv1  gate757(.a(N307), .O(gate124inter8));
  nand2 gate758(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate759(.a(s_85), .b(gate124inter3), .O(gate124inter10));
  nor2  gate760(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate761(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate762(.a(gate124inter12), .b(gate124inter1), .O(N355));

  xor2  gate609(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate610(.a(gate125inter0), .b(s_64), .O(gate125inter1));
  and2  gate611(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate612(.a(s_64), .O(gate125inter3));
  inv1  gate613(.a(s_65), .O(gate125inter4));
  nand2 gate614(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate615(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate616(.a(N343), .O(gate125inter7));
  inv1  gate617(.a(N308), .O(gate125inter8));
  nand2 gate618(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate619(.a(s_65), .b(gate125inter3), .O(gate125inter10));
  nor2  gate620(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate621(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate622(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate245(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate246(.a(gate129inter0), .b(s_12), .O(gate129inter1));
  and2  gate247(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate248(.a(s_12), .O(gate129inter3));
  inv1  gate249(.a(s_13), .O(gate129inter4));
  nand2 gate250(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate251(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate252(.a(N14), .O(gate129inter7));
  inv1  gate253(.a(N360), .O(gate129inter8));
  nand2 gate254(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate255(.a(s_13), .b(gate129inter3), .O(gate129inter10));
  nor2  gate256(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate257(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate258(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate287(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate288(.a(gate132inter0), .b(s_18), .O(gate132inter1));
  and2  gate289(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate290(.a(s_18), .O(gate132inter3));
  inv1  gate291(.a(s_19), .O(gate132inter4));
  nand2 gate292(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate293(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate294(.a(N360), .O(gate132inter7));
  inv1  gate295(.a(N53), .O(gate132inter8));
  nand2 gate296(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate297(.a(s_19), .b(gate132inter3), .O(gate132inter10));
  nor2  gate298(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate299(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate300(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );

  xor2  gate175(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate176(.a(gate134inter0), .b(s_2), .O(gate134inter1));
  and2  gate177(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate178(.a(s_2), .O(gate134inter3));
  inv1  gate179(.a(s_3), .O(gate134inter4));
  nand2 gate180(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate181(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate182(.a(N360), .O(gate134inter7));
  inv1  gate183(.a(N79), .O(gate134inter8));
  nand2 gate184(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate185(.a(s_3), .b(gate134inter3), .O(gate134inter10));
  nor2  gate186(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate187(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate188(.a(gate134inter12), .b(gate134inter1), .O(N376));
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );

  xor2  gate777(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate778(.a(gate137inter0), .b(s_88), .O(gate137inter1));
  and2  gate779(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate780(.a(s_88), .O(gate137inter3));
  inv1  gate781(.a(s_89), .O(gate137inter4));
  nand2 gate782(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate783(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate784(.a(N360), .O(gate137inter7));
  inv1  gate785(.a(N115), .O(gate137inter8));
  nand2 gate786(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate787(.a(s_89), .b(gate137inter3), .O(gate137inter10));
  nor2  gate788(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate789(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate790(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate231(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate232(.a(gate153inter0), .b(s_10), .O(gate153inter1));
  and2  gate233(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate234(.a(s_10), .O(gate153inter3));
  inv1  gate235(.a(s_11), .O(gate153inter4));
  nand2 gate236(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate237(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate238(.a(N415), .O(gate153inter7));
  inv1  gate239(.a(N416), .O(gate153inter8));
  nand2 gate240(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate241(.a(s_11), .b(gate153inter3), .O(gate153inter10));
  nor2  gate242(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate243(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate244(.a(gate153inter12), .b(gate153inter1), .O(N421));
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule