module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate853inter0, gate853inter1, gate853inter2, gate853inter3, gate853inter4, gate853inter5, gate853inter6, gate853inter7, gate853inter8, gate853inter9, gate853inter10, gate853inter11, gate853inter12, gate349inter0, gate349inter1, gate349inter2, gate349inter3, gate349inter4, gate349inter5, gate349inter6, gate349inter7, gate349inter8, gate349inter9, gate349inter10, gate349inter11, gate349inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate552inter0, gate552inter1, gate552inter2, gate552inter3, gate552inter4, gate552inter5, gate552inter6, gate552inter7, gate552inter8, gate552inter9, gate552inter10, gate552inter11, gate552inter12, gate368inter0, gate368inter1, gate368inter2, gate368inter3, gate368inter4, gate368inter5, gate368inter6, gate368inter7, gate368inter8, gate368inter9, gate368inter10, gate368inter11, gate368inter12, gate556inter0, gate556inter1, gate556inter2, gate556inter3, gate556inter4, gate556inter5, gate556inter6, gate556inter7, gate556inter8, gate556inter9, gate556inter10, gate556inter11, gate556inter12, gate340inter0, gate340inter1, gate340inter2, gate340inter3, gate340inter4, gate340inter5, gate340inter6, gate340inter7, gate340inter8, gate340inter9, gate340inter10, gate340inter11, gate340inter12, gate866inter0, gate866inter1, gate866inter2, gate866inter3, gate866inter4, gate866inter5, gate866inter6, gate866inter7, gate866inter8, gate866inter9, gate866inter10, gate866inter11, gate866inter12, gate816inter0, gate816inter1, gate816inter2, gate816inter3, gate816inter4, gate816inter5, gate816inter6, gate816inter7, gate816inter8, gate816inter9, gate816inter10, gate816inter11, gate816inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate519inter0, gate519inter1, gate519inter2, gate519inter3, gate519inter4, gate519inter5, gate519inter6, gate519inter7, gate519inter8, gate519inter9, gate519inter10, gate519inter11, gate519inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate801inter0, gate801inter1, gate801inter2, gate801inter3, gate801inter4, gate801inter5, gate801inter6, gate801inter7, gate801inter8, gate801inter9, gate801inter10, gate801inter11, gate801inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate526inter0, gate526inter1, gate526inter2, gate526inter3, gate526inter4, gate526inter5, gate526inter6, gate526inter7, gate526inter8, gate526inter9, gate526inter10, gate526inter11, gate526inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate618inter0, gate618inter1, gate618inter2, gate618inter3, gate618inter4, gate618inter5, gate618inter6, gate618inter7, gate618inter8, gate618inter9, gate618inter10, gate618inter11, gate618inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate767inter0, gate767inter1, gate767inter2, gate767inter3, gate767inter4, gate767inter5, gate767inter6, gate767inter7, gate767inter8, gate767inter9, gate767inter10, gate767inter11, gate767inter12, gate805inter0, gate805inter1, gate805inter2, gate805inter3, gate805inter4, gate805inter5, gate805inter6, gate805inter7, gate805inter8, gate805inter9, gate805inter10, gate805inter11, gate805inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate766inter0, gate766inter1, gate766inter2, gate766inter3, gate766inter4, gate766inter5, gate766inter6, gate766inter7, gate766inter8, gate766inter9, gate766inter10, gate766inter11, gate766inter12, gate775inter0, gate775inter1, gate775inter2, gate775inter3, gate775inter4, gate775inter5, gate775inter6, gate775inter7, gate775inter8, gate775inter9, gate775inter10, gate775inter11, gate775inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate541inter0, gate541inter1, gate541inter2, gate541inter3, gate541inter4, gate541inter5, gate541inter6, gate541inter7, gate541inter8, gate541inter9, gate541inter10, gate541inter11, gate541inter12, gate826inter0, gate826inter1, gate826inter2, gate826inter3, gate826inter4, gate826inter5, gate826inter6, gate826inter7, gate826inter8, gate826inter9, gate826inter10, gate826inter11, gate826inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate639inter0, gate639inter1, gate639inter2, gate639inter3, gate639inter4, gate639inter5, gate639inter6, gate639inter7, gate639inter8, gate639inter9, gate639inter10, gate639inter11, gate639inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate372inter0, gate372inter1, gate372inter2, gate372inter3, gate372inter4, gate372inter5, gate372inter6, gate372inter7, gate372inter8, gate372inter9, gate372inter10, gate372inter11, gate372inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate769inter0, gate769inter1, gate769inter2, gate769inter3, gate769inter4, gate769inter5, gate769inter6, gate769inter7, gate769inter8, gate769inter9, gate769inter10, gate769inter11, gate769inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate681inter0, gate681inter1, gate681inter2, gate681inter3, gate681inter4, gate681inter5, gate681inter6, gate681inter7, gate681inter8, gate681inter9, gate681inter10, gate681inter11, gate681inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate528inter0, gate528inter1, gate528inter2, gate528inter3, gate528inter4, gate528inter5, gate528inter6, gate528inter7, gate528inter8, gate528inter9, gate528inter10, gate528inter11, gate528inter12, gate679inter0, gate679inter1, gate679inter2, gate679inter3, gate679inter4, gate679inter5, gate679inter6, gate679inter7, gate679inter8, gate679inter9, gate679inter10, gate679inter11, gate679inter12, gate572inter0, gate572inter1, gate572inter2, gate572inter3, gate572inter4, gate572inter5, gate572inter6, gate572inter7, gate572inter8, gate572inter9, gate572inter10, gate572inter11, gate572inter12, gate879inter0, gate879inter1, gate879inter2, gate879inter3, gate879inter4, gate879inter5, gate879inter6, gate879inter7, gate879inter8, gate879inter9, gate879inter10, gate879inter11, gate879inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate682inter0, gate682inter1, gate682inter2, gate682inter3, gate682inter4, gate682inter5, gate682inter6, gate682inter7, gate682inter8, gate682inter9, gate682inter10, gate682inter11, gate682inter12, gate325inter0, gate325inter1, gate325inter2, gate325inter3, gate325inter4, gate325inter5, gate325inter6, gate325inter7, gate325inter8, gate325inter9, gate325inter10, gate325inter11, gate325inter12, gate319inter0, gate319inter1, gate319inter2, gate319inter3, gate319inter4, gate319inter5, gate319inter6, gate319inter7, gate319inter8, gate319inter9, gate319inter10, gate319inter11, gate319inter12, gate545inter0, gate545inter1, gate545inter2, gate545inter3, gate545inter4, gate545inter5, gate545inter6, gate545inter7, gate545inter8, gate545inter9, gate545inter10, gate545inter11, gate545inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate329inter0, gate329inter1, gate329inter2, gate329inter3, gate329inter4, gate329inter5, gate329inter6, gate329inter7, gate329inter8, gate329inter9, gate329inter10, gate329inter11, gate329inter12, gate608inter0, gate608inter1, gate608inter2, gate608inter3, gate608inter4, gate608inter5, gate608inter6, gate608inter7, gate608inter8, gate608inter9, gate608inter10, gate608inter11, gate608inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate536inter0, gate536inter1, gate536inter2, gate536inter3, gate536inter4, gate536inter5, gate536inter6, gate536inter7, gate536inter8, gate536inter9, gate536inter10, gate536inter11, gate536inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate637inter0, gate637inter1, gate637inter2, gate637inter3, gate637inter4, gate637inter5, gate637inter6, gate637inter7, gate637inter8, gate637inter9, gate637inter10, gate637inter11, gate637inter12, gate780inter0, gate780inter1, gate780inter2, gate780inter3, gate780inter4, gate780inter5, gate780inter6, gate780inter7, gate780inter8, gate780inter9, gate780inter10, gate780inter11, gate780inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate378inter0, gate378inter1, gate378inter2, gate378inter3, gate378inter4, gate378inter5, gate378inter6, gate378inter7, gate378inter8, gate378inter9, gate378inter10, gate378inter11, gate378inter12, gate758inter0, gate758inter1, gate758inter2, gate758inter3, gate758inter4, gate758inter5, gate758inter6, gate758inter7, gate758inter8, gate758inter9, gate758inter10, gate758inter11, gate758inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate863inter0, gate863inter1, gate863inter2, gate863inter3, gate863inter4, gate863inter5, gate863inter6, gate863inter7, gate863inter8, gate863inter9, gate863inter10, gate863inter11, gate863inter12, gate818inter0, gate818inter1, gate818inter2, gate818inter3, gate818inter4, gate818inter5, gate818inter6, gate818inter7, gate818inter8, gate818inter9, gate818inter10, gate818inter11, gate818inter12, gate796inter0, gate796inter1, gate796inter2, gate796inter3, gate796inter4, gate796inter5, gate796inter6, gate796inter7, gate796inter8, gate796inter9, gate796inter10, gate796inter11, gate796inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate324inter0, gate324inter1, gate324inter2, gate324inter3, gate324inter4, gate324inter5, gate324inter6, gate324inter7, gate324inter8, gate324inter9, gate324inter10, gate324inter11, gate324inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate338inter0, gate338inter1, gate338inter2, gate338inter3, gate338inter4, gate338inter5, gate338inter6, gate338inter7, gate338inter8, gate338inter9, gate338inter10, gate338inter11, gate338inter12, gate762inter0, gate762inter1, gate762inter2, gate762inter3, gate762inter4, gate762inter5, gate762inter6, gate762inter7, gate762inter8, gate762inter9, gate762inter10, gate762inter11, gate762inter12, gate851inter0, gate851inter1, gate851inter2, gate851inter3, gate851inter4, gate851inter5, gate851inter6, gate851inter7, gate851inter8, gate851inter9, gate851inter10, gate851inter11, gate851inter12, gate303inter0, gate303inter1, gate303inter2, gate303inter3, gate303inter4, gate303inter5, gate303inter6, gate303inter7, gate303inter8, gate303inter9, gate303inter10, gate303inter11, gate303inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate517inter0, gate517inter1, gate517inter2, gate517inter3, gate517inter4, gate517inter5, gate517inter6, gate517inter7, gate517inter8, gate517inter9, gate517inter10, gate517inter11, gate517inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate837inter0, gate837inter1, gate837inter2, gate837inter3, gate837inter4, gate837inter5, gate837inter6, gate837inter7, gate837inter8, gate837inter9, gate837inter10, gate837inter11, gate837inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate357inter0, gate357inter1, gate357inter2, gate357inter3, gate357inter4, gate357inter5, gate357inter6, gate357inter7, gate357inter8, gate357inter9, gate357inter10, gate357inter11, gate357inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate864inter0, gate864inter1, gate864inter2, gate864inter3, gate864inter4, gate864inter5, gate864inter6, gate864inter7, gate864inter8, gate864inter9, gate864inter10, gate864inter11, gate864inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate607inter0, gate607inter1, gate607inter2, gate607inter3, gate607inter4, gate607inter5, gate607inter6, gate607inter7, gate607inter8, gate607inter9, gate607inter10, gate607inter11, gate607inter12, gate852inter0, gate852inter1, gate852inter2, gate852inter3, gate852inter4, gate852inter5, gate852inter6, gate852inter7, gate852inter8, gate852inter9, gate852inter10, gate852inter11, gate852inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate643inter0, gate643inter1, gate643inter2, gate643inter3, gate643inter4, gate643inter5, gate643inter6, gate643inter7, gate643inter8, gate643inter9, gate643inter10, gate643inter11, gate643inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate642inter0, gate642inter1, gate642inter2, gate642inter3, gate642inter4, gate642inter5, gate642inter6, gate642inter7, gate642inter8, gate642inter9, gate642inter10, gate642inter11, gate642inter12, gate855inter0, gate855inter1, gate855inter2, gate855inter3, gate855inter4, gate855inter5, gate855inter6, gate855inter7, gate855inter8, gate855inter9, gate855inter10, gate855inter11, gate855inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate318inter0, gate318inter1, gate318inter2, gate318inter3, gate318inter4, gate318inter5, gate318inter6, gate318inter7, gate318inter8, gate318inter9, gate318inter10, gate318inter11, gate318inter12, gate621inter0, gate621inter1, gate621inter2, gate621inter3, gate621inter4, gate621inter5, gate621inter6, gate621inter7, gate621inter8, gate621inter9, gate621inter10, gate621inter11, gate621inter12, gate321inter0, gate321inter1, gate321inter2, gate321inter3, gate321inter4, gate321inter5, gate321inter6, gate321inter7, gate321inter8, gate321inter9, gate321inter10, gate321inter11, gate321inter12, gate353inter0, gate353inter1, gate353inter2, gate353inter3, gate353inter4, gate353inter5, gate353inter6, gate353inter7, gate353inter8, gate353inter9, gate353inter10, gate353inter11, gate353inter12, gate814inter0, gate814inter1, gate814inter2, gate814inter3, gate814inter4, gate814inter5, gate814inter6, gate814inter7, gate814inter8, gate814inter9, gate814inter10, gate814inter11, gate814inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate640inter0, gate640inter1, gate640inter2, gate640inter3, gate640inter4, gate640inter5, gate640inter6, gate640inter7, gate640inter8, gate640inter9, gate640inter10, gate640inter11, gate640inter12, gate561inter0, gate561inter1, gate561inter2, gate561inter3, gate561inter4, gate561inter5, gate561inter6, gate561inter7, gate561inter8, gate561inter9, gate561inter10, gate561inter11, gate561inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate798inter0, gate798inter1, gate798inter2, gate798inter3, gate798inter4, gate798inter5, gate798inter6, gate798inter7, gate798inter8, gate798inter9, gate798inter10, gate798inter11, gate798inter12, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate854inter0, gate854inter1, gate854inter2, gate854inter3, gate854inter4, gate854inter5, gate854inter6, gate854inter7, gate854inter8, gate854inter9, gate854inter10, gate854inter11, gate854inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate624inter0, gate624inter1, gate624inter2, gate624inter3, gate624inter4, gate624inter5, gate624inter6, gate624inter7, gate624inter8, gate624inter9, gate624inter10, gate624inter11, gate624inter12;



inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );

  xor2  gate2379(.a(N331), .b(N306), .O(gate75inter0));
  nand2 gate2380(.a(gate75inter0), .b(s_214), .O(gate75inter1));
  and2  gate2381(.a(N331), .b(N306), .O(gate75inter2));
  inv1  gate2382(.a(s_214), .O(gate75inter3));
  inv1  gate2383(.a(s_215), .O(gate75inter4));
  nand2 gate2384(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2385(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2386(.a(N306), .O(gate75inter7));
  inv1  gate2387(.a(N331), .O(gate75inter8));
  nand2 gate2388(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2389(.a(s_215), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2390(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2391(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2392(.a(gate75inter12), .b(gate75inter1), .O(N550));
nand2 gate76( .a(N306), .b(N331), .O(N551) );

  xor2  gate1147(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate1148(.a(gate77inter0), .b(s_38), .O(gate77inter1));
  and2  gate1149(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate1150(.a(s_38), .O(gate77inter3));
  inv1  gate1151(.a(s_39), .O(gate77inter4));
  nand2 gate1152(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1153(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1154(.a(N306), .O(gate77inter7));
  inv1  gate1155(.a(N331), .O(gate77inter8));
  nand2 gate1156(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1157(.a(s_39), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1158(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1159(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1160(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );

  xor2  gate1077(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate1078(.a(gate79inter0), .b(s_28), .O(gate79inter1));
  and2  gate1079(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate1080(.a(s_28), .O(gate79inter3));
  inv1  gate1081(.a(s_29), .O(gate79inter4));
  nand2 gate1082(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1083(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1084(.a(N306), .O(gate79inter7));
  inv1  gate1085(.a(N331), .O(gate79inter8));
  nand2 gate1086(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1087(.a(s_29), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1088(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1089(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1090(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate2631(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate2632(.a(gate96inter0), .b(s_250), .O(gate96inter1));
  and2  gate2633(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate2634(.a(s_250), .O(gate96inter3));
  inv1  gate2635(.a(s_251), .O(gate96inter4));
  nand2 gate2636(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2637(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2638(.a(N326), .O(gate96inter7));
  inv1  gate2639(.a(N277), .O(gate96inter8));
  nand2 gate2640(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2641(.a(s_251), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2642(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2643(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2644(.a(gate96inter12), .b(gate96inter1), .O(N601));
nand2 gate97( .a(N326), .b(N280), .O(N602) );

  xor2  gate2001(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate2002(.a(gate98inter0), .b(s_160), .O(gate98inter1));
  and2  gate2003(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate2004(.a(s_160), .O(gate98inter3));
  inv1  gate2005(.a(s_161), .O(gate98inter4));
  nand2 gate2006(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2007(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2008(.a(N260), .O(gate98inter7));
  inv1  gate2009(.a(N72), .O(gate98inter8));
  nand2 gate2010(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2011(.a(s_161), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2012(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2013(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2014(.a(gate98inter12), .b(gate98inter1), .O(N603));
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );

  xor2  gate1875(.a(N608), .b(N60), .O(gate161inter0));
  nand2 gate1876(.a(gate161inter0), .b(s_142), .O(gate161inter1));
  and2  gate1877(.a(N608), .b(N60), .O(gate161inter2));
  inv1  gate1878(.a(s_142), .O(gate161inter3));
  inv1  gate1879(.a(s_143), .O(gate161inter4));
  nand2 gate1880(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1881(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1882(.a(N60), .O(gate161inter7));
  inv1  gate1883(.a(N608), .O(gate161inter8));
  nand2 gate1884(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1885(.a(s_143), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1886(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1887(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1888(.a(gate161inter12), .b(gate161inter1), .O(N903));
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );

  xor2  gate1483(.a(N889), .b(N616), .O(gate234inter0));
  nand2 gate1484(.a(gate234inter0), .b(s_86), .O(gate234inter1));
  and2  gate1485(.a(N889), .b(N616), .O(gate234inter2));
  inv1  gate1486(.a(s_86), .O(gate234inter3));
  inv1  gate1487(.a(s_87), .O(gate234inter4));
  nand2 gate1488(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1489(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1490(.a(N616), .O(gate234inter7));
  inv1  gate1491(.a(N889), .O(gate234inter8));
  nand2 gate1492(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1493(.a(s_87), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1494(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1495(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1496(.a(gate234inter12), .b(gate234inter1), .O(N1055));
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );

  xor2  gate2267(.a(N895), .b(N655), .O(gate237inter0));
  nand2 gate2268(.a(gate237inter0), .b(s_198), .O(gate237inter1));
  and2  gate2269(.a(N895), .b(N655), .O(gate237inter2));
  inv1  gate2270(.a(s_198), .O(gate237inter3));
  inv1  gate2271(.a(s_199), .O(gate237inter4));
  nand2 gate2272(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2273(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2274(.a(N655), .O(gate237inter7));
  inv1  gate2275(.a(N895), .O(gate237inter8));
  nand2 gate2276(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2277(.a(s_199), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2278(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2279(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2280(.a(gate237inter12), .b(gate237inter1), .O(N1067));

  xor2  gate1665(.a(N896), .b(N652), .O(gate238inter0));
  nand2 gate1666(.a(gate238inter0), .b(s_112), .O(gate238inter1));
  and2  gate1667(.a(N896), .b(N652), .O(gate238inter2));
  inv1  gate1668(.a(s_112), .O(gate238inter3));
  inv1  gate1669(.a(s_113), .O(gate238inter4));
  nand2 gate1670(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1671(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1672(.a(N652), .O(gate238inter7));
  inv1  gate1673(.a(N896), .O(gate238inter8));
  nand2 gate1674(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1675(.a(s_113), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1676(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1677(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1678(.a(gate238inter12), .b(gate238inter1), .O(N1068));
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );

  xor2  gate2435(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate2436(.a(gate245inter0), .b(s_222), .O(gate245inter1));
  and2  gate2437(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate2438(.a(s_222), .O(gate245inter3));
  inv1  gate2439(.a(s_223), .O(gate245inter4));
  nand2 gate2440(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2441(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2442(.a(N745), .O(gate245inter7));
  inv1  gate2443(.a(N1005), .O(gate245inter8));
  nand2 gate2444(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2445(.a(s_223), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2446(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2447(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2448(.a(gate245inter12), .b(gate245inter1), .O(N1130));
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );

  xor2  gate2183(.a(N1008), .b(N751), .O(gate247inter0));
  nand2 gate2184(.a(gate247inter0), .b(s_186), .O(gate247inter1));
  and2  gate2185(.a(N1008), .b(N751), .O(gate247inter2));
  inv1  gate2186(.a(s_186), .O(gate247inter3));
  inv1  gate2187(.a(s_187), .O(gate247inter4));
  nand2 gate2188(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2189(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2190(.a(N751), .O(gate247inter7));
  inv1  gate2191(.a(N1008), .O(gate247inter8));
  nand2 gate2192(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2193(.a(s_187), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2194(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2195(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2196(.a(gate247inter12), .b(gate247inter1), .O(N1132));

  xor2  gate2561(.a(N1009), .b(N748), .O(gate248inter0));
  nand2 gate2562(.a(gate248inter0), .b(s_240), .O(gate248inter1));
  and2  gate2563(.a(N1009), .b(N748), .O(gate248inter2));
  inv1  gate2564(.a(s_240), .O(gate248inter3));
  inv1  gate2565(.a(s_241), .O(gate248inter4));
  nand2 gate2566(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2567(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2568(.a(N748), .O(gate248inter7));
  inv1  gate2569(.a(N1009), .O(gate248inter8));
  nand2 gate2570(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2571(.a(s_241), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2572(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2573(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2574(.a(gate248inter12), .b(gate248inter1), .O(N1133));
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );

  xor2  gate2015(.a(N1064), .b(N1063), .O(gate259inter0));
  nand2 gate2016(.a(gate259inter0), .b(s_162), .O(gate259inter1));
  and2  gate2017(.a(N1064), .b(N1063), .O(gate259inter2));
  inv1  gate2018(.a(s_162), .O(gate259inter3));
  inv1  gate2019(.a(s_163), .O(gate259inter4));
  nand2 gate2020(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2021(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2022(.a(N1063), .O(gate259inter7));
  inv1  gate2023(.a(N1064), .O(gate259inter8));
  nand2 gate2024(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2025(.a(s_163), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2026(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2027(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2028(.a(gate259inter12), .b(gate259inter1), .O(N1158));
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate1007(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate1008(.a(gate268inter0), .b(s_18), .O(gate268inter1));
  and2  gate1009(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate1010(.a(s_18), .O(gate268inter3));
  inv1  gate1011(.a(s_19), .O(gate268inter4));
  nand2 gate1012(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1013(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1014(.a(N921), .O(gate268inter7));
  inv1  gate1015(.a(N923), .O(gate268inter8));
  nand2 gate1016(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1017(.a(s_19), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1018(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1019(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1020(.a(gate268inter12), .b(gate268inter1), .O(N1171));

  xor2  gate2477(.a(N923), .b(N922), .O(gate269inter0));
  nand2 gate2478(.a(gate269inter0), .b(s_228), .O(gate269inter1));
  and2  gate2479(.a(N923), .b(N922), .O(gate269inter2));
  inv1  gate2480(.a(s_228), .O(gate269inter3));
  inv1  gate2481(.a(s_229), .O(gate269inter4));
  nand2 gate2482(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2483(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2484(.a(N922), .O(gate269inter7));
  inv1  gate2485(.a(N923), .O(gate269inter8));
  nand2 gate2486(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2487(.a(s_229), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2488(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2489(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2490(.a(gate269inter12), .b(gate269inter1), .O(N1188));
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate2225(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate2226(.a(gate273inter0), .b(s_192), .O(gate273inter1));
  and2  gate2227(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate2228(.a(s_192), .O(gate273inter3));
  inv1  gate2229(.a(s_193), .O(gate273inter4));
  nand2 gate2230(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2231(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2232(.a(N1013), .O(gate273inter7));
  inv1  gate2233(.a(N942), .O(gate273inter8));
  nand2 gate2234(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2235(.a(s_193), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2236(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2237(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2238(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );

  xor2  gate1917(.a(N958), .b(N1025), .O(gate281inter0));
  nand2 gate1918(.a(gate281inter0), .b(s_148), .O(gate281inter1));
  and2  gate1919(.a(N958), .b(N1025), .O(gate281inter2));
  inv1  gate1920(.a(s_148), .O(gate281inter3));
  inv1  gate1921(.a(s_149), .O(gate281inter4));
  nand2 gate1922(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1923(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1924(.a(N1025), .O(gate281inter7));
  inv1  gate1925(.a(N958), .O(gate281inter8));
  nand2 gate1926(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1927(.a(s_149), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1928(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1929(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1930(.a(gate281inter12), .b(gate281inter1), .O(N1216));
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );

  xor2  gate2645(.a(N968), .b(N1034), .O(gate286inter0));
  nand2 gate2646(.a(gate286inter0), .b(s_252), .O(gate286inter1));
  and2  gate2647(.a(N968), .b(N1034), .O(gate286inter2));
  inv1  gate2648(.a(s_252), .O(gate286inter3));
  inv1  gate2649(.a(s_253), .O(gate286inter4));
  nand2 gate2650(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2651(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2652(.a(N1034), .O(gate286inter7));
  inv1  gate2653(.a(N968), .O(gate286inter8));
  nand2 gate2654(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2655(.a(s_253), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2656(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2657(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2658(.a(gate286inter12), .b(gate286inter1), .O(N1221));
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );

  xor2  gate1161(.a(N972), .b(N1037), .O(gate289inter0));
  nand2 gate1162(.a(gate289inter0), .b(s_40), .O(gate289inter1));
  and2  gate1163(.a(N972), .b(N1037), .O(gate289inter2));
  inv1  gate1164(.a(s_40), .O(gate289inter3));
  inv1  gate1165(.a(s_41), .O(gate289inter4));
  nand2 gate1166(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1167(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1168(.a(N1037), .O(gate289inter7));
  inv1  gate1169(.a(N972), .O(gate289inter8));
  nand2 gate1170(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1171(.a(s_41), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1172(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1173(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1174(.a(gate289inter12), .b(gate289inter1), .O(N1224));
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );

  xor2  gate1189(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate1190(.a(gate298inter0), .b(s_44), .O(gate298inter1));
  and2  gate1191(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate1192(.a(s_44), .O(gate298inter3));
  inv1  gate1193(.a(s_45), .O(gate298inter4));
  nand2 gate1194(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate1195(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate1196(.a(N1121), .O(gate298inter7));
  inv1  gate1197(.a(N1122), .O(gate298inter8));
  nand2 gate1198(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate1199(.a(s_45), .b(gate298inter3), .O(gate298inter10));
  nor2  gate1200(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate1201(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate1202(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );

  xor2  gate2113(.a(N1001), .b(N1049), .O(gate303inter0));
  nand2 gate2114(.a(gate303inter0), .b(s_176), .O(gate303inter1));
  and2  gate2115(.a(N1001), .b(N1049), .O(gate303inter2));
  inv1  gate2116(.a(s_176), .O(gate303inter3));
  inv1  gate2117(.a(s_177), .O(gate303inter4));
  nand2 gate2118(.a(gate303inter4), .b(gate303inter3), .O(gate303inter5));
  nor2  gate2119(.a(gate303inter5), .b(gate303inter2), .O(gate303inter6));
  inv1  gate2120(.a(N1049), .O(gate303inter7));
  inv1  gate2121(.a(N1001), .O(gate303inter8));
  nand2 gate2122(.a(gate303inter8), .b(gate303inter7), .O(gate303inter9));
  nand2 gate2123(.a(s_177), .b(gate303inter3), .O(gate303inter10));
  nor2  gate2124(.a(gate303inter10), .b(gate303inter9), .O(gate303inter11));
  nor2  gate2125(.a(gate303inter11), .b(gate303inter6), .O(gate303inter12));
  nand2 gate2126(.a(gate303inter12), .b(gate303inter1), .O(N1242));
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );

  xor2  gate2757(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate2758(.a(gate316inter0), .b(s_268), .O(gate316inter1));
  and2  gate2759(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate2760(.a(s_268), .O(gate316inter3));
  inv1  gate2761(.a(s_269), .O(gate316inter4));
  nand2 gate2762(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate2763(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate2764(.a(N697), .O(gate316inter7));
  inv1  gate2765(.a(N1211), .O(gate316inter8));
  nand2 gate2766(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate2767(.a(s_269), .b(gate316inter3), .O(gate316inter10));
  nor2  gate2768(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate2769(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate2770(.a(gate316inter12), .b(gate316inter1), .O(N1312));
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );

  xor2  gate2491(.a(N1215), .b(N703), .O(gate318inter0));
  nand2 gate2492(.a(gate318inter0), .b(s_230), .O(gate318inter1));
  and2  gate2493(.a(N1215), .b(N703), .O(gate318inter2));
  inv1  gate2494(.a(s_230), .O(gate318inter3));
  inv1  gate2495(.a(s_231), .O(gate318inter4));
  nand2 gate2496(.a(gate318inter4), .b(gate318inter3), .O(gate318inter5));
  nor2  gate2497(.a(gate318inter5), .b(gate318inter2), .O(gate318inter6));
  inv1  gate2498(.a(N703), .O(gate318inter7));
  inv1  gate2499(.a(N1215), .O(gate318inter8));
  nand2 gate2500(.a(gate318inter8), .b(gate318inter7), .O(gate318inter9));
  nand2 gate2501(.a(s_231), .b(gate318inter3), .O(gate318inter10));
  nor2  gate2502(.a(gate318inter10), .b(gate318inter9), .O(gate318inter11));
  nor2  gate2503(.a(gate318inter11), .b(gate318inter6), .O(gate318inter12));
  nand2 gate2504(.a(gate318inter12), .b(gate318inter1), .O(N1314));

  xor2  gate1707(.a(N1220), .b(N706), .O(gate319inter0));
  nand2 gate1708(.a(gate319inter0), .b(s_118), .O(gate319inter1));
  and2  gate1709(.a(N1220), .b(N706), .O(gate319inter2));
  inv1  gate1710(.a(s_118), .O(gate319inter3));
  inv1  gate1711(.a(s_119), .O(gate319inter4));
  nand2 gate1712(.a(gate319inter4), .b(gate319inter3), .O(gate319inter5));
  nor2  gate1713(.a(gate319inter5), .b(gate319inter2), .O(gate319inter6));
  inv1  gate1714(.a(N706), .O(gate319inter7));
  inv1  gate1715(.a(N1220), .O(gate319inter8));
  nand2 gate1716(.a(gate319inter8), .b(gate319inter7), .O(gate319inter9));
  nand2 gate1717(.a(s_119), .b(gate319inter3), .O(gate319inter10));
  nor2  gate1718(.a(gate319inter10), .b(gate319inter9), .O(gate319inter11));
  nor2  gate1719(.a(gate319inter11), .b(gate319inter6), .O(gate319inter12));
  nand2 gate1720(.a(gate319inter12), .b(gate319inter1), .O(N1315));
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );

  xor2  gate2519(.a(N1225), .b(N712), .O(gate321inter0));
  nand2 gate2520(.a(gate321inter0), .b(s_234), .O(gate321inter1));
  and2  gate2521(.a(N1225), .b(N712), .O(gate321inter2));
  inv1  gate2522(.a(s_234), .O(gate321inter3));
  inv1  gate2523(.a(s_235), .O(gate321inter4));
  nand2 gate2524(.a(gate321inter4), .b(gate321inter3), .O(gate321inter5));
  nor2  gate2525(.a(gate321inter5), .b(gate321inter2), .O(gate321inter6));
  inv1  gate2526(.a(N712), .O(gate321inter7));
  inv1  gate2527(.a(N1225), .O(gate321inter8));
  nand2 gate2528(.a(gate321inter8), .b(gate321inter7), .O(gate321inter9));
  nand2 gate2529(.a(s_235), .b(gate321inter3), .O(gate321inter10));
  nor2  gate2530(.a(gate321inter10), .b(gate321inter9), .O(gate321inter11));
  nor2  gate2531(.a(gate321inter11), .b(gate321inter6), .O(gate321inter12));
  nand2 gate2532(.a(gate321inter12), .b(gate321inter1), .O(N1317));
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );

  xor2  gate2043(.a(N1230), .b(N628), .O(gate324inter0));
  nand2 gate2044(.a(gate324inter0), .b(s_166), .O(gate324inter1));
  and2  gate2045(.a(N1230), .b(N628), .O(gate324inter2));
  inv1  gate2046(.a(s_166), .O(gate324inter3));
  inv1  gate2047(.a(s_167), .O(gate324inter4));
  nand2 gate2048(.a(gate324inter4), .b(gate324inter3), .O(gate324inter5));
  nor2  gate2049(.a(gate324inter5), .b(gate324inter2), .O(gate324inter6));
  inv1  gate2050(.a(N628), .O(gate324inter7));
  inv1  gate2051(.a(N1230), .O(gate324inter8));
  nand2 gate2052(.a(gate324inter8), .b(gate324inter7), .O(gate324inter9));
  nand2 gate2053(.a(s_167), .b(gate324inter3), .O(gate324inter10));
  nor2  gate2054(.a(gate324inter10), .b(gate324inter9), .O(gate324inter11));
  nor2  gate2055(.a(gate324inter11), .b(gate324inter6), .O(gate324inter12));
  nand2 gate2056(.a(gate324inter12), .b(gate324inter1), .O(N1322));

  xor2  gate1693(.a(N1238), .b(N730), .O(gate325inter0));
  nand2 gate1694(.a(gate325inter0), .b(s_116), .O(gate325inter1));
  and2  gate1695(.a(N1238), .b(N730), .O(gate325inter2));
  inv1  gate1696(.a(s_116), .O(gate325inter3));
  inv1  gate1697(.a(s_117), .O(gate325inter4));
  nand2 gate1698(.a(gate325inter4), .b(gate325inter3), .O(gate325inter5));
  nor2  gate1699(.a(gate325inter5), .b(gate325inter2), .O(gate325inter6));
  inv1  gate1700(.a(N730), .O(gate325inter7));
  inv1  gate1701(.a(N1238), .O(gate325inter8));
  nand2 gate1702(.a(gate325inter8), .b(gate325inter7), .O(gate325inter9));
  nand2 gate1703(.a(s_117), .b(gate325inter3), .O(gate325inter10));
  nor2  gate1704(.a(gate325inter10), .b(gate325inter9), .O(gate325inter11));
  nor2  gate1705(.a(gate325inter11), .b(gate325inter6), .O(gate325inter12));
  nand2 gate1706(.a(gate325inter12), .b(gate325inter1), .O(N1327));
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );

  xor2  gate1791(.a(N1160), .b(N1267), .O(gate328inter0));
  nand2 gate1792(.a(gate328inter0), .b(s_130), .O(gate328inter1));
  and2  gate1793(.a(N1160), .b(N1267), .O(gate328inter2));
  inv1  gate1794(.a(s_130), .O(gate328inter3));
  inv1  gate1795(.a(s_131), .O(gate328inter4));
  nand2 gate1796(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate1797(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate1798(.a(N1267), .O(gate328inter7));
  inv1  gate1799(.a(N1160), .O(gate328inter8));
  nand2 gate1800(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate1801(.a(s_131), .b(gate328inter3), .O(gate328inter10));
  nor2  gate1802(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate1803(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate1804(.a(gate328inter12), .b(gate328inter1), .O(N1344));

  xor2  gate1749(.a(N894), .b(N1249), .O(gate329inter0));
  nand2 gate1750(.a(gate329inter0), .b(s_124), .O(gate329inter1));
  and2  gate1751(.a(N894), .b(N1249), .O(gate329inter2));
  inv1  gate1752(.a(s_124), .O(gate329inter3));
  inv1  gate1753(.a(s_125), .O(gate329inter4));
  nand2 gate1754(.a(gate329inter4), .b(gate329inter3), .O(gate329inter5));
  nor2  gate1755(.a(gate329inter5), .b(gate329inter2), .O(gate329inter6));
  inv1  gate1756(.a(N1249), .O(gate329inter7));
  inv1  gate1757(.a(N894), .O(gate329inter8));
  nand2 gate1758(.a(gate329inter8), .b(gate329inter7), .O(gate329inter9));
  nand2 gate1759(.a(s_125), .b(gate329inter3), .O(gate329inter10));
  nor2  gate1760(.a(gate329inter10), .b(gate329inter9), .O(gate329inter11));
  nor2  gate1761(.a(gate329inter11), .b(gate329inter6), .O(gate329inter12));
  nand2 gate1762(.a(gate329inter12), .b(gate329inter1), .O(N1345));
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );

  xor2  gate2253(.a(N1206), .b(N1309), .O(gate335inter0));
  nand2 gate2254(.a(gate335inter0), .b(s_196), .O(gate335inter1));
  and2  gate2255(.a(N1206), .b(N1309), .O(gate335inter2));
  inv1  gate2256(.a(s_196), .O(gate335inter3));
  inv1  gate2257(.a(s_197), .O(gate335inter4));
  nand2 gate2258(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate2259(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate2260(.a(N1309), .O(gate335inter7));
  inv1  gate2261(.a(N1206), .O(gate335inter8));
  nand2 gate2262(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate2263(.a(s_197), .b(gate335inter3), .O(gate335inter10));
  nor2  gate2264(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate2265(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate2266(.a(gate335inter12), .b(gate335inter1), .O(N1352));
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );

  xor2  gate2071(.a(N1212), .b(N1312), .O(gate338inter0));
  nand2 gate2072(.a(gate338inter0), .b(s_170), .O(gate338inter1));
  and2  gate2073(.a(N1212), .b(N1312), .O(gate338inter2));
  inv1  gate2074(.a(s_170), .O(gate338inter3));
  inv1  gate2075(.a(s_171), .O(gate338inter4));
  nand2 gate2076(.a(gate338inter4), .b(gate338inter3), .O(gate338inter5));
  nor2  gate2077(.a(gate338inter5), .b(gate338inter2), .O(gate338inter6));
  inv1  gate2078(.a(N1312), .O(gate338inter7));
  inv1  gate2079(.a(N1212), .O(gate338inter8));
  nand2 gate2080(.a(gate338inter8), .b(gate338inter7), .O(gate338inter9));
  nand2 gate2081(.a(s_171), .b(gate338inter3), .O(gate338inter10));
  nor2  gate2082(.a(gate338inter10), .b(gate338inter9), .O(gate338inter11));
  nor2  gate2083(.a(gate338inter11), .b(gate338inter6), .O(gate338inter12));
  nand2 gate2084(.a(gate338inter12), .b(gate338inter1), .O(N1361));
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );

  xor2  gate965(.a(N1216), .b(N1314), .O(gate340inter0));
  nand2 gate966(.a(gate340inter0), .b(s_12), .O(gate340inter1));
  and2  gate967(.a(N1216), .b(N1314), .O(gate340inter2));
  inv1  gate968(.a(s_12), .O(gate340inter3));
  inv1  gate969(.a(s_13), .O(gate340inter4));
  nand2 gate970(.a(gate340inter4), .b(gate340inter3), .O(gate340inter5));
  nor2  gate971(.a(gate340inter5), .b(gate340inter2), .O(gate340inter6));
  inv1  gate972(.a(N1314), .O(gate340inter7));
  inv1  gate973(.a(N1216), .O(gate340inter8));
  nand2 gate974(.a(gate340inter8), .b(gate340inter7), .O(gate340inter9));
  nand2 gate975(.a(s_13), .b(gate340inter3), .O(gate340inter10));
  nor2  gate976(.a(gate340inter10), .b(gate340inter9), .O(gate340inter11));
  nor2  gate977(.a(gate340inter11), .b(gate340inter6), .O(gate340inter12));
  nand2 gate978(.a(gate340inter12), .b(gate340inter1), .O(N1367));
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );

  xor2  gate1287(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate1288(.a(gate342inter0), .b(s_58), .O(gate342inter1));
  and2  gate1289(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate1290(.a(s_58), .O(gate342inter3));
  inv1  gate1291(.a(s_59), .O(gate342inter4));
  nand2 gate1292(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate1293(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate1294(.a(N1316), .O(gate342inter7));
  inv1  gate1295(.a(N1224), .O(gate342inter8));
  nand2 gate1296(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate1297(.a(s_59), .b(gate342inter3), .O(gate342inter10));
  nor2  gate1298(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate1299(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate1300(.a(gate342inter12), .b(gate342inter1), .O(N1373));
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate1539(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate1540(.a(gate347inter0), .b(s_94), .O(gate347inter1));
  and2  gate1541(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate1542(.a(s_94), .O(gate347inter3));
  inv1  gate1543(.a(s_95), .O(gate347inter4));
  nand2 gate1544(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate1545(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate1546(.a(N1232), .O(gate347inter7));
  inv1  gate1547(.a(N990), .O(gate347inter8));
  nand2 gate1548(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate1549(.a(s_95), .b(gate347inter3), .O(gate347inter10));
  nor2  gate1550(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate1551(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate1552(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );

  xor2  gate895(.a(N993), .b(N1235), .O(gate349inter0));
  nand2 gate896(.a(gate349inter0), .b(s_2), .O(gate349inter1));
  and2  gate897(.a(N993), .b(N1235), .O(gate349inter2));
  inv1  gate898(.a(s_2), .O(gate349inter3));
  inv1  gate899(.a(s_3), .O(gate349inter4));
  nand2 gate900(.a(gate349inter4), .b(gate349inter3), .O(gate349inter5));
  nor2  gate901(.a(gate349inter5), .b(gate349inter2), .O(gate349inter6));
  inv1  gate902(.a(N1235), .O(gate349inter7));
  inv1  gate903(.a(N993), .O(gate349inter8));
  nand2 gate904(.a(gate349inter8), .b(gate349inter7), .O(gate349inter9));
  nand2 gate905(.a(s_3), .b(gate349inter3), .O(gate349inter10));
  nor2  gate906(.a(gate349inter10), .b(gate349inter9), .O(gate349inter11));
  nor2  gate907(.a(gate349inter11), .b(gate349inter6), .O(gate349inter12));
  nand2 gate908(.a(gate349inter12), .b(gate349inter1), .O(N1389));
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );

  xor2  gate2533(.a(N1004), .b(N1243), .O(gate353inter0));
  nand2 gate2534(.a(gate353inter0), .b(s_236), .O(gate353inter1));
  and2  gate2535(.a(N1004), .b(N1243), .O(gate353inter2));
  inv1  gate2536(.a(s_236), .O(gate353inter3));
  inv1  gate2537(.a(s_237), .O(gate353inter4));
  nand2 gate2538(.a(gate353inter4), .b(gate353inter3), .O(gate353inter5));
  nor2  gate2539(.a(gate353inter5), .b(gate353inter2), .O(gate353inter6));
  inv1  gate2540(.a(N1243), .O(gate353inter7));
  inv1  gate2541(.a(N1004), .O(gate353inter8));
  nand2 gate2542(.a(gate353inter8), .b(gate353inter7), .O(gate353inter9));
  nand2 gate2543(.a(s_237), .b(gate353inter3), .O(gate353inter10));
  nor2  gate2544(.a(gate353inter10), .b(gate353inter9), .O(gate353inter11));
  nor2  gate2545(.a(gate353inter11), .b(gate353inter6), .O(gate353inter12));
  nand2 gate2546(.a(gate353inter12), .b(gate353inter1), .O(N1397));
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );

  xor2  gate2281(.a(N1346), .b(N649), .O(gate357inter0));
  nand2 gate2282(.a(gate357inter0), .b(s_200), .O(gate357inter1));
  and2  gate2283(.a(N1346), .b(N649), .O(gate357inter2));
  inv1  gate2284(.a(s_200), .O(gate357inter3));
  inv1  gate2285(.a(s_201), .O(gate357inter4));
  nand2 gate2286(.a(gate357inter4), .b(gate357inter3), .O(gate357inter5));
  nor2  gate2287(.a(gate357inter5), .b(gate357inter2), .O(gate357inter6));
  inv1  gate2288(.a(N649), .O(gate357inter7));
  inv1  gate2289(.a(N1346), .O(gate357inter8));
  nand2 gate2290(.a(gate357inter8), .b(gate357inter7), .O(gate357inter9));
  nand2 gate2291(.a(s_201), .b(gate357inter3), .O(gate357inter10));
  nor2  gate2292(.a(gate357inter10), .b(gate357inter9), .O(gate357inter11));
  nor2  gate2293(.a(gate357inter11), .b(gate357inter6), .O(gate357inter12));
  nand2 gate2294(.a(gate357inter12), .b(gate357inter1), .O(N1412));
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );

  xor2  gate1735(.a(N1388), .b(N637), .O(gate362inter0));
  nand2 gate1736(.a(gate362inter0), .b(s_122), .O(gate362inter1));
  and2  gate1737(.a(N1388), .b(N637), .O(gate362inter2));
  inv1  gate1738(.a(s_122), .O(gate362inter3));
  inv1  gate1739(.a(s_123), .O(gate362inter4));
  nand2 gate1740(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate1741(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate1742(.a(N637), .O(gate362inter7));
  inv1  gate1743(.a(N1388), .O(gate362inter8));
  nand2 gate1744(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate1745(.a(s_123), .b(gate362inter3), .O(gate362inter10));
  nor2  gate1746(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate1747(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate1748(.a(gate362inter12), .b(gate362inter1), .O(N1434));
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );

  xor2  gate937(.a(N1149), .b(N1352), .O(gate368inter0));
  nand2 gate938(.a(gate368inter0), .b(s_8), .O(gate368inter1));
  and2  gate939(.a(N1149), .b(N1352), .O(gate368inter2));
  inv1  gate940(.a(s_8), .O(gate368inter3));
  inv1  gate941(.a(s_9), .O(gate368inter4));
  nand2 gate942(.a(gate368inter4), .b(gate368inter3), .O(gate368inter5));
  nor2  gate943(.a(gate368inter5), .b(gate368inter2), .O(gate368inter6));
  inv1  gate944(.a(N1352), .O(gate368inter7));
  inv1  gate945(.a(N1149), .O(gate368inter8));
  nand2 gate946(.a(gate368inter8), .b(gate368inter7), .O(gate368inter9));
  nand2 gate947(.a(s_9), .b(gate368inter3), .O(gate368inter10));
  nor2  gate948(.a(gate368inter10), .b(gate368inter9), .O(gate368inter11));
  nor2  gate949(.a(gate368inter11), .b(gate368inter6), .O(gate368inter12));
  nand2 gate950(.a(gate368inter12), .b(gate368inter1), .O(N1445));
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );

  xor2  gate1497(.a(N1152), .b(N1361), .O(gate372inter0));
  nand2 gate1498(.a(gate372inter0), .b(s_88), .O(gate372inter1));
  and2  gate1499(.a(N1152), .b(N1361), .O(gate372inter2));
  inv1  gate1500(.a(s_88), .O(gate372inter3));
  inv1  gate1501(.a(s_89), .O(gate372inter4));
  nand2 gate1502(.a(gate372inter4), .b(gate372inter3), .O(gate372inter5));
  nor2  gate1503(.a(gate372inter5), .b(gate372inter2), .O(gate372inter6));
  inv1  gate1504(.a(N1361), .O(gate372inter7));
  inv1  gate1505(.a(N1152), .O(gate372inter8));
  nand2 gate1506(.a(gate372inter8), .b(gate372inter7), .O(gate372inter9));
  nand2 gate1507(.a(s_89), .b(gate372inter3), .O(gate372inter10));
  nor2  gate1508(.a(gate372inter10), .b(gate372inter9), .O(gate372inter11));
  nor2  gate1509(.a(gate372inter11), .b(gate372inter6), .O(gate372inter12));
  nand2 gate1510(.a(gate372inter12), .b(gate372inter1), .O(N1451));
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );

  xor2  gate1889(.a(N1156), .b(N1373), .O(gate378inter0));
  nand2 gate1890(.a(gate378inter0), .b(s_144), .O(gate378inter1));
  and2  gate1891(.a(N1156), .b(N1373), .O(gate378inter2));
  inv1  gate1892(.a(s_144), .O(gate378inter3));
  inv1  gate1893(.a(s_145), .O(gate378inter4));
  nand2 gate1894(.a(gate378inter4), .b(gate378inter3), .O(gate378inter5));
  nor2  gate1895(.a(gate378inter5), .b(gate378inter2), .O(gate378inter6));
  inv1  gate1896(.a(N1373), .O(gate378inter7));
  inv1  gate1897(.a(N1156), .O(gate378inter8));
  nand2 gate1898(.a(gate378inter8), .b(gate378inter7), .O(gate378inter9));
  nand2 gate1899(.a(s_145), .b(gate378inter3), .O(gate378inter10));
  nor2  gate1900(.a(gate378inter10), .b(gate378inter9), .O(gate378inter11));
  nor2  gate1901(.a(gate378inter11), .b(gate378inter6), .O(gate378inter12));
  nand2 gate1902(.a(gate378inter12), .b(gate378inter1), .O(N1457));
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate1945(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate1946(.a(gate383inter0), .b(s_152), .O(gate383inter1));
  and2  gate1947(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate1948(.a(s_152), .O(gate383inter3));
  inv1  gate1949(.a(s_153), .O(gate383inter4));
  nand2 gate1950(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate1951(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate1952(.a(N1393), .O(gate383inter7));
  inv1  gate1953(.a(N1161), .O(gate383inter8));
  nand2 gate1954(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate1955(.a(s_153), .b(gate383inter3), .O(gate383inter10));
  nor2  gate1956(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate1957(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate1958(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );

  xor2  gate1567(.a(N1227), .b(N1376), .O(gate389inter0));
  nand2 gate1568(.a(gate389inter0), .b(s_98), .O(gate389inter1));
  and2  gate1569(.a(N1227), .b(N1376), .O(gate389inter2));
  inv1  gate1570(.a(s_98), .O(gate389inter3));
  inv1  gate1571(.a(s_99), .O(gate389inter4));
  nand2 gate1572(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1573(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1574(.a(N1376), .O(gate389inter7));
  inv1  gate1575(.a(N1227), .O(gate389inter8));
  nand2 gate1576(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1577(.a(s_99), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1578(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1579(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1580(.a(gate389inter12), .b(gate389inter1), .O(N1471));
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );

  xor2  gate1021(.a(N1240), .b(N1390), .O(gate392inter0));
  nand2 gate1022(.a(gate392inter0), .b(s_20), .O(gate392inter1));
  and2  gate1023(.a(N1240), .b(N1390), .O(gate392inter2));
  inv1  gate1024(.a(s_20), .O(gate392inter3));
  inv1  gate1025(.a(s_21), .O(gate392inter4));
  nand2 gate1026(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1027(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1028(.a(N1390), .O(gate392inter7));
  inv1  gate1029(.a(N1240), .O(gate392inter8));
  nand2 gate1030(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1031(.a(s_21), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1032(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1033(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1034(.a(gate392inter12), .b(gate392inter1), .O(N1476));
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );

  xor2  gate1777(.a(N1439), .b(N1399), .O(gate394inter0));
  nand2 gate1778(.a(gate394inter0), .b(s_128), .O(gate394inter1));
  and2  gate1779(.a(N1439), .b(N1399), .O(gate394inter2));
  inv1  gate1780(.a(s_128), .O(gate394inter3));
  inv1  gate1781(.a(s_129), .O(gate394inter4));
  nand2 gate1782(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1783(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1784(.a(N1399), .O(gate394inter7));
  inv1  gate1785(.a(N1439), .O(gate394inter8));
  nand2 gate1786(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1787(.a(s_129), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1788(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1789(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1790(.a(gate394inter12), .b(gate394inter1), .O(N1481));
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );

  xor2  gate2603(.a(N1448), .b(N943), .O(gate398inter0));
  nand2 gate2604(.a(gate398inter0), .b(s_246), .O(gate398inter1));
  and2  gate2605(.a(N1448), .b(N943), .O(gate398inter2));
  inv1  gate2606(.a(s_246), .O(gate398inter3));
  inv1  gate2607(.a(s_247), .O(gate398inter4));
  nand2 gate2608(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2609(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2610(.a(N943), .O(gate398inter7));
  inv1  gate2611(.a(N1448), .O(gate398inter8));
  nand2 gate2612(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2613(.a(s_247), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2614(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2615(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2616(.a(gate398inter12), .b(gate398inter1), .O(N1489));
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );

  xor2  gate2715(.a(N1458), .b(N969), .O(gate404inter0));
  nand2 gate2716(.a(gate404inter0), .b(s_262), .O(gate404inter1));
  and2  gate2717(.a(N1458), .b(N969), .O(gate404inter2));
  inv1  gate2718(.a(s_262), .O(gate404inter3));
  inv1  gate2719(.a(s_263), .O(gate404inter4));
  nand2 gate2720(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2721(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2722(.a(N969), .O(gate404inter7));
  inv1  gate2723(.a(N1458), .O(gate404inter8));
  nand2 gate2724(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2725(.a(s_263), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2726(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2727(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2728(.a(gate404inter12), .b(gate404inter1), .O(N1495));
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );

  xor2  gate1301(.a(N1468), .b(N965), .O(gate408inter0));
  nand2 gate1302(.a(gate408inter0), .b(s_60), .O(gate408inter1));
  and2  gate1303(.a(N1468), .b(N965), .O(gate408inter2));
  inv1  gate1304(.a(s_60), .O(gate408inter3));
  inv1  gate1305(.a(s_61), .O(gate408inter4));
  nand2 gate1306(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1307(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1308(.a(N965), .O(gate408inter7));
  inv1  gate1309(.a(N1468), .O(gate408inter8));
  nand2 gate1310(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1311(.a(s_61), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1312(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1313(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1314(.a(gate408inter12), .b(gate408inter1), .O(N1500));

  xor2  gate2197(.a(N1470), .b(N973), .O(gate409inter0));
  nand2 gate2198(.a(gate409inter0), .b(s_188), .O(gate409inter1));
  and2  gate2199(.a(N1470), .b(N973), .O(gate409inter2));
  inv1  gate2200(.a(s_188), .O(gate409inter3));
  inv1  gate2201(.a(s_189), .O(gate409inter4));
  nand2 gate2202(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2203(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2204(.a(N973), .O(gate409inter7));
  inv1  gate2205(.a(N1470), .O(gate409inter8));
  nand2 gate2206(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2207(.a(s_189), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2208(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2209(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2210(.a(gate409inter12), .b(gate409inter1), .O(N1501));

  xor2  gate2743(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate2744(.a(gate410inter0), .b(s_266), .O(gate410inter1));
  and2  gate2745(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate2746(.a(s_266), .O(gate410inter3));
  inv1  gate2747(.a(s_267), .O(gate410inter4));
  nand2 gate2748(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2749(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2750(.a(N994), .O(gate410inter7));
  inv1  gate2751(.a(N1475), .O(gate410inter8));
  nand2 gate2752(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2753(.a(s_267), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2754(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2755(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2756(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );

  xor2  gate1049(.a(N1501), .b(N1471), .O(gate425inter0));
  nand2 gate1050(.a(gate425inter0), .b(s_24), .O(gate425inter1));
  and2  gate1051(.a(N1501), .b(N1471), .O(gate425inter2));
  inv1  gate1052(.a(s_24), .O(gate425inter3));
  inv1  gate1053(.a(s_25), .O(gate425inter4));
  nand2 gate1054(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1055(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1056(.a(N1471), .O(gate425inter7));
  inv1  gate1057(.a(N1501), .O(gate425inter8));
  nand2 gate1058(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1059(.a(s_25), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1060(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1061(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1062(.a(gate425inter12), .b(gate425inter1), .O(N1534));
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );

  xor2  gate2295(.a(N1530), .b(N1540), .O(gate440inter0));
  nand2 gate2296(.a(gate440inter0), .b(s_202), .O(gate440inter1));
  and2  gate2297(.a(N1530), .b(N1540), .O(gate440inter2));
  inv1  gate2298(.a(s_202), .O(gate440inter3));
  inv1  gate2299(.a(s_203), .O(gate440inter4));
  nand2 gate2300(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2301(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2302(.a(N1540), .O(gate440inter7));
  inv1  gate2303(.a(N1530), .O(gate440inter8));
  nand2 gate2304(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2305(.a(s_203), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2306(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2307(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2308(.a(gate440inter12), .b(gate440inter1), .O(N1594));
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );

  xor2  gate1273(.a(N893), .b(N1596), .O(gate462inter0));
  nand2 gate1274(.a(gate462inter0), .b(s_56), .O(gate462inter1));
  and2  gate1275(.a(N893), .b(N1596), .O(gate462inter2));
  inv1  gate1276(.a(s_56), .O(gate462inter3));
  inv1  gate1277(.a(s_57), .O(gate462inter4));
  nand2 gate1278(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1279(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1280(.a(N1596), .O(gate462inter7));
  inv1  gate1281(.a(N893), .O(gate462inter8));
  nand2 gate1282(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1283(.a(s_57), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1284(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1285(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1286(.a(gate462inter12), .b(gate462inter1), .O(N1671));
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );

  xor2  gate1595(.a(N1636), .b(N1594), .O(gate472inter0));
  nand2 gate1596(.a(gate472inter0), .b(s_102), .O(gate472inter1));
  and2  gate1597(.a(N1636), .b(N1594), .O(gate472inter2));
  inv1  gate1598(.a(s_102), .O(gate472inter3));
  inv1  gate1599(.a(s_103), .O(gate472inter4));
  nand2 gate1600(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1601(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1602(.a(N1594), .O(gate472inter7));
  inv1  gate1603(.a(N1636), .O(gate472inter8));
  nand2 gate1604(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1605(.a(s_103), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1606(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1607(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1608(.a(gate472inter12), .b(gate472inter1), .O(N1685));

  xor2  gate1259(.a(N1639), .b(N1510), .O(gate473inter0));
  nand2 gate1260(.a(gate473inter0), .b(s_54), .O(gate473inter1));
  and2  gate1261(.a(N1639), .b(N1510), .O(gate473inter2));
  inv1  gate1262(.a(s_54), .O(gate473inter3));
  inv1  gate1263(.a(s_55), .O(gate473inter4));
  nand2 gate1264(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1265(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1266(.a(N1510), .O(gate473inter7));
  inv1  gate1267(.a(N1639), .O(gate473inter8));
  nand2 gate1268(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1269(.a(s_55), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1270(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1271(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1272(.a(gate473inter12), .b(gate473inter1), .O(N1688));
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );

  xor2  gate2617(.a(N1681), .b(N1031), .O(gate483inter0));
  nand2 gate2618(.a(gate483inter0), .b(s_248), .O(gate483inter1));
  and2  gate2619(.a(N1681), .b(N1031), .O(gate483inter2));
  inv1  gate2620(.a(s_248), .O(gate483inter3));
  inv1  gate2621(.a(s_249), .O(gate483inter4));
  nand2 gate2622(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2623(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2624(.a(N1031), .O(gate483inter7));
  inv1  gate2625(.a(N1681), .O(gate483inter8));
  nand2 gate2626(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2627(.a(s_249), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2628(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2629(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2630(.a(gate483inter12), .b(gate483inter1), .O(N1713));
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );

  xor2  gate1931(.a(N1528), .b(N1685), .O(gate494inter0));
  nand2 gate1932(.a(gate494inter0), .b(s_150), .O(gate494inter1));
  and2  gate1933(.a(N1528), .b(N1685), .O(gate494inter2));
  inv1  gate1934(.a(s_150), .O(gate494inter3));
  inv1  gate1935(.a(s_151), .O(gate494inter4));
  nand2 gate1936(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1937(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1938(.a(N1685), .O(gate494inter7));
  inv1  gate1939(.a(N1528), .O(gate494inter8));
  nand2 gate1940(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1941(.a(s_151), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1942(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1943(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1944(.a(gate494inter12), .b(gate494inter1), .O(N1740));
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );

  xor2  gate2393(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate2394(.a(gate499inter0), .b(s_216), .O(gate499inter1));
  and2  gate2395(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate2396(.a(s_216), .O(gate499inter3));
  inv1  gate2397(.a(s_217), .O(gate499inter4));
  nand2 gate2398(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2399(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2400(.a(N1678), .O(gate499inter7));
  inv1  gate2401(.a(N1712), .O(gate499inter8));
  nand2 gate2402(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2403(.a(s_217), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2404(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2405(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2406(.a(gate499inter12), .b(gate499inter1), .O(N1748));

  xor2  gate2239(.a(N1713), .b(N1680), .O(gate500inter0));
  nand2 gate2240(.a(gate500inter0), .b(s_194), .O(gate500inter1));
  and2  gate2241(.a(N1713), .b(N1680), .O(gate500inter2));
  inv1  gate2242(.a(s_194), .O(gate500inter3));
  inv1  gate2243(.a(s_195), .O(gate500inter4));
  nand2 gate2244(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2245(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2246(.a(N1680), .O(gate500inter7));
  inv1  gate2247(.a(N1713), .O(gate500inter8));
  nand2 gate2248(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2249(.a(s_195), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2250(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2251(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2252(.a(gate500inter12), .b(gate500inter1), .O(N1751));
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );

  xor2  gate2155(.a(N1730), .b(N1701), .O(gate505inter0));
  nand2 gate2156(.a(gate505inter0), .b(s_182), .O(gate505inter1));
  and2  gate2157(.a(N1730), .b(N1701), .O(gate505inter2));
  inv1  gate2158(.a(s_182), .O(gate505inter3));
  inv1  gate2159(.a(s_183), .O(gate505inter4));
  nand2 gate2160(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2161(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2162(.a(N1701), .O(gate505inter7));
  inv1  gate2163(.a(N1730), .O(gate505inter8));
  nand2 gate2164(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2165(.a(s_183), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2166(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2167(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2168(.a(gate505inter12), .b(gate505inter1), .O(N1764));
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );

  xor2  gate1231(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate1232(.a(gate508inter0), .b(s_50), .O(gate508inter1));
  and2  gate1233(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate1234(.a(s_50), .O(gate508inter3));
  inv1  gate1235(.a(s_51), .O(gate508inter4));
  nand2 gate1236(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1237(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1238(.a(N1723), .O(gate508inter7));
  inv1  gate1239(.a(N1413), .O(gate508inter8));
  nand2 gate1240(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1241(.a(s_51), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1242(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1243(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1244(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );

  xor2  gate909(.a(N1746), .b(N1708), .O(gate510inter0));
  nand2 gate910(.a(gate510inter0), .b(s_4), .O(gate510inter1));
  and2  gate911(.a(N1746), .b(N1708), .O(gate510inter2));
  inv1  gate912(.a(s_4), .O(gate510inter3));
  inv1  gate913(.a(s_5), .O(gate510inter4));
  nand2 gate914(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate915(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate916(.a(N1708), .O(gate510inter7));
  inv1  gate917(.a(N1746), .O(gate510inter8));
  nand2 gate918(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate919(.a(s_5), .b(gate510inter3), .O(gate510inter10));
  nor2  gate920(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate921(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate922(.a(gate510inter12), .b(gate510inter1), .O(N1774));
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1245(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1246(.a(gate513inter0), .b(s_52), .O(gate513inter1));
  and2  gate1247(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1248(.a(s_52), .O(gate513inter3));
  inv1  gate1249(.a(s_53), .O(gate513inter4));
  nand2 gate1250(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1251(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1252(.a(N1731), .O(gate513inter7));
  inv1  gate1253(.a(N1682), .O(gate513inter8));
  nand2 gate1254(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1255(.a(s_53), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1256(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1257(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1258(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );

  xor2  gate2141(.a(N1759), .b(N1720), .O(gate517inter0));
  nand2 gate2142(.a(gate517inter0), .b(s_180), .O(gate517inter1));
  and2  gate2143(.a(N1759), .b(N1720), .O(gate517inter2));
  inv1  gate2144(.a(s_180), .O(gate517inter3));
  inv1  gate2145(.a(s_181), .O(gate517inter4));
  nand2 gate2146(.a(gate517inter4), .b(gate517inter3), .O(gate517inter5));
  nor2  gate2147(.a(gate517inter5), .b(gate517inter2), .O(gate517inter6));
  inv1  gate2148(.a(N1720), .O(gate517inter7));
  inv1  gate2149(.a(N1759), .O(gate517inter8));
  nand2 gate2150(.a(gate517inter8), .b(gate517inter7), .O(gate517inter9));
  nand2 gate2151(.a(s_181), .b(gate517inter3), .O(gate517inter10));
  nor2  gate2152(.a(gate517inter10), .b(gate517inter9), .O(gate517inter11));
  nor2  gate2153(.a(gate517inter11), .b(gate517inter6), .O(gate517inter12));
  nand2 gate2154(.a(gate517inter12), .b(gate517inter1), .O(N1788));
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );

  xor2  gate1035(.a(N1763), .b(N1664), .O(gate519inter0));
  nand2 gate1036(.a(gate519inter0), .b(s_22), .O(gate519inter1));
  and2  gate1037(.a(N1763), .b(N1664), .O(gate519inter2));
  inv1  gate1038(.a(s_22), .O(gate519inter3));
  inv1  gate1039(.a(s_23), .O(gate519inter4));
  nand2 gate1040(.a(gate519inter4), .b(gate519inter3), .O(gate519inter5));
  nor2  gate1041(.a(gate519inter5), .b(gate519inter2), .O(gate519inter6));
  inv1  gate1042(.a(N1664), .O(gate519inter7));
  inv1  gate1043(.a(N1763), .O(gate519inter8));
  nand2 gate1044(.a(gate519inter8), .b(gate519inter7), .O(gate519inter9));
  nand2 gate1045(.a(s_23), .b(gate519inter3), .O(gate519inter10));
  nor2  gate1046(.a(gate519inter10), .b(gate519inter9), .O(gate519inter11));
  nor2  gate1047(.a(gate519inter11), .b(gate519inter6), .O(gate519inter12));
  nand2 gate1048(.a(gate519inter12), .b(gate519inter1), .O(N1792));

  xor2  gate1217(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate1218(.a(gate520inter0), .b(s_48), .O(gate520inter1));
  and2  gate1219(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate1220(.a(s_48), .O(gate520inter3));
  inv1  gate1221(.a(s_49), .O(gate520inter4));
  nand2 gate1222(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate1223(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate1224(.a(N1751), .O(gate520inter7));
  inv1  gate1225(.a(N1155), .O(gate520inter8));
  nand2 gate1226(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate1227(.a(s_49), .b(gate520inter3), .O(gate520inter10));
  nor2  gate1228(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate1229(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate1230(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate1385(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate1386(.a(gate522inter0), .b(s_72), .O(gate522inter1));
  and2  gate1387(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate1388(.a(s_72), .O(gate522inter3));
  inv1  gate1389(.a(s_73), .O(gate522inter4));
  nand2 gate1390(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate1391(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate1392(.a(N1740), .O(gate522inter7));
  inv1  gate1393(.a(N1769), .O(gate522inter8));
  nand2 gate1394(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate1395(.a(s_73), .b(gate522inter3), .O(gate522inter10));
  nor2  gate1396(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate1397(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate1398(.a(gate522inter12), .b(gate522inter1), .O(N1798));
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );

  xor2  gate1175(.a(N1218), .b(N1748), .O(gate526inter0));
  nand2 gate1176(.a(gate526inter0), .b(s_42), .O(gate526inter1));
  and2  gate1177(.a(N1218), .b(N1748), .O(gate526inter2));
  inv1  gate1178(.a(s_42), .O(gate526inter3));
  inv1  gate1179(.a(s_43), .O(gate526inter4));
  nand2 gate1180(.a(gate526inter4), .b(gate526inter3), .O(gate526inter5));
  nor2  gate1181(.a(gate526inter5), .b(gate526inter2), .O(gate526inter6));
  inv1  gate1182(.a(N1748), .O(gate526inter7));
  inv1  gate1183(.a(N1218), .O(gate526inter8));
  nand2 gate1184(.a(gate526inter8), .b(gate526inter7), .O(gate526inter9));
  nand2 gate1185(.a(s_43), .b(gate526inter3), .O(gate526inter10));
  nor2  gate1186(.a(gate526inter10), .b(gate526inter9), .O(gate526inter11));
  nor2  gate1187(.a(gate526inter11), .b(gate526inter6), .O(gate526inter12));
  nand2 gate1188(.a(gate526inter12), .b(gate526inter1), .O(N1808));
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );

  xor2  gate1609(.a(N1786), .b(N1615), .O(gate528inter0));
  nand2 gate1610(.a(gate528inter0), .b(s_104), .O(gate528inter1));
  and2  gate1611(.a(N1786), .b(N1615), .O(gate528inter2));
  inv1  gate1612(.a(s_104), .O(gate528inter3));
  inv1  gate1613(.a(s_105), .O(gate528inter4));
  nand2 gate1614(.a(gate528inter4), .b(gate528inter3), .O(gate528inter5));
  nor2  gate1615(.a(gate528inter5), .b(gate528inter2), .O(gate528inter6));
  inv1  gate1616(.a(N1615), .O(gate528inter7));
  inv1  gate1617(.a(N1786), .O(gate528inter8));
  nand2 gate1618(.a(gate528inter8), .b(gate528inter7), .O(gate528inter9));
  nand2 gate1619(.a(s_105), .b(gate528inter3), .O(gate528inter10));
  nor2  gate1620(.a(gate528inter10), .b(gate528inter9), .O(gate528inter11));
  nor2  gate1621(.a(gate528inter11), .b(gate528inter6), .O(gate528inter12));
  nand2 gate1622(.a(gate528inter12), .b(gate528inter1), .O(N1810));
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate2029(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate2030(.a(gate532inter0), .b(s_164), .O(gate532inter1));
  and2  gate2031(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate2032(.a(s_164), .O(gate532inter3));
  inv1  gate2033(.a(s_165), .O(gate532inter4));
  nand2 gate2034(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate2035(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate2036(.a(N1777), .O(gate532inter7));
  inv1  gate2037(.a(N1490), .O(gate532inter8));
  nand2 gate2038(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate2039(.a(s_165), .b(gate532inter3), .O(gate532inter10));
  nor2  gate2040(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate2041(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate2042(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );

  xor2  gate1805(.a(N1796), .b(N962), .O(gate536inter0));
  nand2 gate1806(.a(gate536inter0), .b(s_132), .O(gate536inter1));
  and2  gate1807(.a(N1796), .b(N962), .O(gate536inter2));
  inv1  gate1808(.a(s_132), .O(gate536inter3));
  inv1  gate1809(.a(s_133), .O(gate536inter4));
  nand2 gate1810(.a(gate536inter4), .b(gate536inter3), .O(gate536inter5));
  nor2  gate1811(.a(gate536inter5), .b(gate536inter2), .O(gate536inter6));
  inv1  gate1812(.a(N962), .O(gate536inter7));
  inv1  gate1813(.a(N1796), .O(gate536inter8));
  nand2 gate1814(.a(gate536inter8), .b(gate536inter7), .O(gate536inter9));
  nand2 gate1815(.a(s_133), .b(gate536inter3), .O(gate536inter10));
  nor2  gate1816(.a(gate536inter10), .b(gate536inter9), .O(gate536inter11));
  nor2  gate1817(.a(gate536inter11), .b(gate536inter6), .O(gate536inter12));
  nand2 gate1818(.a(gate536inter12), .b(gate536inter1), .O(N1825));
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );

  xor2  gate1427(.a(N1784), .b(N1809), .O(gate541inter0));
  nand2 gate1428(.a(gate541inter0), .b(s_78), .O(gate541inter1));
  and2  gate1429(.a(N1784), .b(N1809), .O(gate541inter2));
  inv1  gate1430(.a(s_78), .O(gate541inter3));
  inv1  gate1431(.a(s_79), .O(gate541inter4));
  nand2 gate1432(.a(gate541inter4), .b(gate541inter3), .O(gate541inter5));
  nor2  gate1433(.a(gate541inter5), .b(gate541inter2), .O(gate541inter6));
  inv1  gate1434(.a(N1809), .O(gate541inter7));
  inv1  gate1435(.a(N1784), .O(gate541inter8));
  nand2 gate1436(.a(gate541inter8), .b(gate541inter7), .O(gate541inter9));
  nand2 gate1437(.a(s_79), .b(gate541inter3), .O(gate541inter10));
  nor2  gate1438(.a(gate541inter10), .b(gate541inter9), .O(gate541inter11));
  nor2  gate1439(.a(gate541inter11), .b(gate541inter6), .O(gate541inter12));
  nand2 gate1440(.a(gate541inter12), .b(gate541inter1), .O(N1838));
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );

  xor2  gate1721(.a(N1825), .b(N1795), .O(gate545inter0));
  nand2 gate1722(.a(gate545inter0), .b(s_120), .O(gate545inter1));
  and2  gate1723(.a(N1825), .b(N1795), .O(gate545inter2));
  inv1  gate1724(.a(s_120), .O(gate545inter3));
  inv1  gate1725(.a(s_121), .O(gate545inter4));
  nand2 gate1726(.a(gate545inter4), .b(gate545inter3), .O(gate545inter5));
  nor2  gate1727(.a(gate545inter5), .b(gate545inter2), .O(gate545inter6));
  inv1  gate1728(.a(N1795), .O(gate545inter7));
  inv1  gate1729(.a(N1825), .O(gate545inter8));
  nand2 gate1730(.a(gate545inter8), .b(gate545inter7), .O(gate545inter9));
  nand2 gate1731(.a(s_121), .b(gate545inter3), .O(gate545inter10));
  nor2  gate1732(.a(gate545inter10), .b(gate545inter9), .O(gate545inter11));
  nor2  gate1733(.a(gate545inter11), .b(gate545inter6), .O(gate545inter12));
  nand2 gate1734(.a(gate545inter12), .b(gate545inter1), .O(N1850));
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );

  xor2  gate1063(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate1064(.a(gate547inter0), .b(s_26), .O(gate547inter1));
  and2  gate1065(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate1066(.a(s_26), .O(gate547inter3));
  inv1  gate1067(.a(s_27), .O(gate547inter4));
  nand2 gate1068(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate1069(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate1070(.a(N1815), .O(gate547inter7));
  inv1  gate1071(.a(N1707), .O(gate547inter8));
  nand2 gate1072(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate1073(.a(s_27), .b(gate547inter3), .O(gate547inter10));
  nor2  gate1074(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate1075(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate1076(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );

  xor2  gate923(.a(N1728), .b(N1812), .O(gate552inter0));
  nand2 gate924(.a(gate552inter0), .b(s_6), .O(gate552inter1));
  and2  gate925(.a(N1728), .b(N1812), .O(gate552inter2));
  inv1  gate926(.a(s_6), .O(gate552inter3));
  inv1  gate927(.a(s_7), .O(gate552inter4));
  nand2 gate928(.a(gate552inter4), .b(gate552inter3), .O(gate552inter5));
  nor2  gate929(.a(gate552inter5), .b(gate552inter2), .O(gate552inter6));
  inv1  gate930(.a(N1812), .O(gate552inter7));
  inv1  gate931(.a(N1728), .O(gate552inter8));
  nand2 gate932(.a(gate552inter8), .b(gate552inter7), .O(gate552inter9));
  nand2 gate933(.a(s_7), .b(gate552inter3), .O(gate552inter10));
  nor2  gate934(.a(gate552inter10), .b(gate552inter9), .O(gate552inter11));
  nor2  gate935(.a(gate552inter11), .b(gate552inter6), .O(gate552inter12));
  nand2 gate936(.a(gate552inter12), .b(gate552inter1), .O(N1865));
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );

  xor2  gate951(.a(N1837), .b(N1808), .O(gate556inter0));
  nand2 gate952(.a(gate556inter0), .b(s_10), .O(gate556inter1));
  and2  gate953(.a(N1837), .b(N1808), .O(gate556inter2));
  inv1  gate954(.a(s_10), .O(gate556inter3));
  inv1  gate955(.a(s_11), .O(gate556inter4));
  nand2 gate956(.a(gate556inter4), .b(gate556inter3), .O(gate556inter5));
  nor2  gate957(.a(gate556inter5), .b(gate556inter2), .O(gate556inter6));
  inv1  gate958(.a(N1808), .O(gate556inter7));
  inv1  gate959(.a(N1837), .O(gate556inter8));
  nand2 gate960(.a(gate556inter8), .b(gate556inter7), .O(gate556inter9));
  nand2 gate961(.a(s_11), .b(gate556inter3), .O(gate556inter10));
  nor2  gate962(.a(gate556inter10), .b(gate556inter9), .O(gate556inter11));
  nor2  gate963(.a(gate556inter11), .b(gate556inter6), .O(gate556inter12));
  nand2 gate964(.a(gate556inter12), .b(gate556inter1), .O(N1875));

  xor2  gate1819(.a(N1848), .b(N1821), .O(gate557inter0));
  nand2 gate1820(.a(gate557inter0), .b(s_134), .O(gate557inter1));
  and2  gate1821(.a(N1848), .b(N1821), .O(gate557inter2));
  inv1  gate1822(.a(s_134), .O(gate557inter3));
  inv1  gate1823(.a(s_135), .O(gate557inter4));
  nand2 gate1824(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate1825(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate1826(.a(N1821), .O(gate557inter7));
  inv1  gate1827(.a(N1848), .O(gate557inter8));
  nand2 gate1828(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate1829(.a(s_135), .b(gate557inter3), .O(gate557inter10));
  nor2  gate1830(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate1831(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate1832(.a(gate557inter12), .b(gate557inter1), .O(N1878));
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );

  xor2  gate2589(.a(N1852), .b(N1826), .O(gate561inter0));
  nand2 gate2590(.a(gate561inter0), .b(s_244), .O(gate561inter1));
  and2  gate2591(.a(N1852), .b(N1826), .O(gate561inter2));
  inv1  gate2592(.a(s_244), .O(gate561inter3));
  inv1  gate2593(.a(s_245), .O(gate561inter4));
  nand2 gate2594(.a(gate561inter4), .b(gate561inter3), .O(gate561inter5));
  nor2  gate2595(.a(gate561inter5), .b(gate561inter2), .O(gate561inter6));
  inv1  gate2596(.a(N1826), .O(gate561inter7));
  inv1  gate2597(.a(N1852), .O(gate561inter8));
  nand2 gate2598(.a(gate561inter8), .b(gate561inter7), .O(gate561inter9));
  nand2 gate2599(.a(s_245), .b(gate561inter3), .O(gate561inter10));
  nor2  gate2600(.a(gate561inter10), .b(gate561inter9), .O(gate561inter11));
  nor2  gate2601(.a(gate561inter11), .b(gate561inter6), .O(gate561inter12));
  nand2 gate2602(.a(gate561inter12), .b(gate561inter1), .O(N1884));

  xor2  gate2659(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate2660(.a(gate562inter0), .b(s_254), .O(gate562inter1));
  and2  gate2661(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate2662(.a(s_254), .O(gate562inter3));
  inv1  gate2663(.a(s_255), .O(gate562inter4));
  nand2 gate2664(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate2665(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate2666(.a(N1643), .O(gate562inter7));
  inv1  gate2667(.a(N1856), .O(gate562inter8));
  nand2 gate2668(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate2669(.a(s_255), .b(gate562inter3), .O(gate562inter10));
  nor2  gate2670(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate2671(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate2672(.a(gate562inter12), .b(gate562inter1), .O(N1885));
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate1091(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate1092(.a(gate565inter0), .b(s_30), .O(gate565inter1));
  and2  gate1093(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate1094(.a(s_30), .O(gate565inter3));
  inv1  gate1095(.a(s_31), .O(gate565inter4));
  nand2 gate1096(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate1097(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate1098(.a(N1838), .O(gate565inter7));
  inv1  gate1099(.a(N1785), .O(gate565inter8));
  nand2 gate1100(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate1101(.a(s_31), .b(gate565inter3), .O(gate565inter10));
  nor2  gate1102(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate1103(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate1104(.a(gate565inter12), .b(gate565inter1), .O(N1896));

  xor2  gate2127(.a(N1864), .b(N1640), .O(gate566inter0));
  nand2 gate2128(.a(gate566inter0), .b(s_178), .O(gate566inter1));
  and2  gate2129(.a(N1864), .b(N1640), .O(gate566inter2));
  inv1  gate2130(.a(s_178), .O(gate566inter3));
  inv1  gate2131(.a(s_179), .O(gate566inter4));
  nand2 gate2132(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate2133(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate2134(.a(N1640), .O(gate566inter7));
  inv1  gate2135(.a(N1864), .O(gate566inter8));
  nand2 gate2136(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate2137(.a(s_179), .b(gate566inter3), .O(gate566inter10));
  nor2  gate2138(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate2139(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate2140(.a(gate566inter12), .b(gate566inter1), .O(N1897));
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );

  xor2  gate1637(.a(N1885), .b(N1855), .O(gate572inter0));
  nand2 gate1638(.a(gate572inter0), .b(s_108), .O(gate572inter1));
  and2  gate1639(.a(N1885), .b(N1855), .O(gate572inter2));
  inv1  gate1640(.a(s_108), .O(gate572inter3));
  inv1  gate1641(.a(s_109), .O(gate572inter4));
  nand2 gate1642(.a(gate572inter4), .b(gate572inter3), .O(gate572inter5));
  nor2  gate1643(.a(gate572inter5), .b(gate572inter2), .O(gate572inter6));
  inv1  gate1644(.a(N1855), .O(gate572inter7));
  inv1  gate1645(.a(N1885), .O(gate572inter8));
  nand2 gate1646(.a(gate572inter8), .b(gate572inter7), .O(gate572inter9));
  nand2 gate1647(.a(s_109), .b(gate572inter3), .O(gate572inter10));
  nor2  gate1648(.a(gate572inter10), .b(gate572inter9), .O(gate572inter11));
  nor2  gate1649(.a(gate572inter11), .b(gate572inter6), .O(gate572inter12));
  nand2 gate1650(.a(gate572inter12), .b(gate572inter1), .O(N1913));
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate2337(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate2338(.a(gate579inter0), .b(s_208), .O(gate579inter1));
  and2  gate2339(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate2340(.a(s_208), .O(gate579inter3));
  inv1  gate2341(.a(s_209), .O(gate579inter4));
  nand2 gate2342(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate2343(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate2344(.a(N1714), .O(gate579inter7));
  inv1  gate2345(.a(N1895), .O(gate579inter8));
  nand2 gate2346(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate2347(.a(s_209), .b(gate579inter3), .O(gate579inter10));
  nor2  gate2348(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate2349(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate2350(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );

  xor2  gate1861(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate1862(.a(gate601inter0), .b(s_140), .O(gate601inter1));
  and2  gate1863(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate1864(.a(s_140), .O(gate601inter3));
  inv1  gate1865(.a(s_141), .O(gate601inter4));
  nand2 gate1866(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate1867(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate1868(.a(N1921), .O(gate601inter7));
  inv1  gate1869(.a(N1942), .O(gate601inter8));
  nand2 gate1870(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate1871(.a(s_141), .b(gate601inter3), .O(gate601inter10));
  nor2  gate1872(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate1873(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate1874(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );

  xor2  gate2351(.a(N1499), .b(N1947), .O(gate607inter0));
  nand2 gate2352(.a(gate607inter0), .b(s_210), .O(gate607inter1));
  and2  gate2353(.a(N1499), .b(N1947), .O(gate607inter2));
  inv1  gate2354(.a(s_210), .O(gate607inter3));
  inv1  gate2355(.a(s_211), .O(gate607inter4));
  nand2 gate2356(.a(gate607inter4), .b(gate607inter3), .O(gate607inter5));
  nor2  gate2357(.a(gate607inter5), .b(gate607inter2), .O(gate607inter6));
  inv1  gate2358(.a(N1947), .O(gate607inter7));
  inv1  gate2359(.a(N1499), .O(gate607inter8));
  nand2 gate2360(.a(gate607inter8), .b(gate607inter7), .O(gate607inter9));
  nand2 gate2361(.a(s_211), .b(gate607inter3), .O(gate607inter10));
  nor2  gate2362(.a(gate607inter10), .b(gate607inter9), .O(gate607inter11));
  nor2  gate2363(.a(gate607inter11), .b(gate607inter6), .O(gate607inter12));
  nand2 gate2364(.a(gate607inter12), .b(gate607inter1), .O(N2003));

  xor2  gate1763(.a(N1350), .b(N1953), .O(gate608inter0));
  nand2 gate1764(.a(gate608inter0), .b(s_126), .O(gate608inter1));
  and2  gate1765(.a(N1350), .b(N1953), .O(gate608inter2));
  inv1  gate1766(.a(s_126), .O(gate608inter3));
  inv1  gate1767(.a(s_127), .O(gate608inter4));
  nand2 gate1768(.a(gate608inter4), .b(gate608inter3), .O(gate608inter5));
  nor2  gate1769(.a(gate608inter5), .b(gate608inter2), .O(gate608inter6));
  inv1  gate1770(.a(N1953), .O(gate608inter7));
  inv1  gate1771(.a(N1350), .O(gate608inter8));
  nand2 gate1772(.a(gate608inter8), .b(gate608inter7), .O(gate608inter9));
  nand2 gate1773(.a(s_127), .b(gate608inter3), .O(gate608inter10));
  nor2  gate1774(.a(gate608inter10), .b(gate608inter9), .O(gate608inter11));
  nor2  gate1775(.a(gate608inter11), .b(gate608inter6), .O(gate608inter12));
  nand2 gate1776(.a(gate608inter12), .b(gate608inter1), .O(N2004));
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );

  xor2  gate1203(.a(N1635), .b(N1961), .O(gate618inter0));
  nand2 gate1204(.a(gate618inter0), .b(s_46), .O(gate618inter1));
  and2  gate1205(.a(N1635), .b(N1961), .O(gate618inter2));
  inv1  gate1206(.a(s_46), .O(gate618inter3));
  inv1  gate1207(.a(s_47), .O(gate618inter4));
  nand2 gate1208(.a(gate618inter4), .b(gate618inter3), .O(gate618inter5));
  nor2  gate1209(.a(gate618inter5), .b(gate618inter2), .O(gate618inter6));
  inv1  gate1210(.a(N1961), .O(gate618inter7));
  inv1  gate1211(.a(N1635), .O(gate618inter8));
  nand2 gate1212(.a(gate618inter8), .b(gate618inter7), .O(gate618inter9));
  nand2 gate1213(.a(s_47), .b(gate618inter3), .O(gate618inter10));
  nor2  gate1214(.a(gate618inter10), .b(gate618inter9), .O(gate618inter11));
  nor2  gate1215(.a(gate618inter11), .b(gate618inter6), .O(gate618inter12));
  nand2 gate1216(.a(gate618inter12), .b(gate618inter1), .O(N2016));
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );

  xor2  gate2505(.a(N1999), .b(N1898), .O(gate621inter0));
  nand2 gate2506(.a(gate621inter0), .b(s_232), .O(gate621inter1));
  and2  gate2507(.a(N1999), .b(N1898), .O(gate621inter2));
  inv1  gate2508(.a(s_232), .O(gate621inter3));
  inv1  gate2509(.a(s_233), .O(gate621inter4));
  nand2 gate2510(.a(gate621inter4), .b(gate621inter3), .O(gate621inter5));
  nor2  gate2511(.a(gate621inter5), .b(gate621inter2), .O(gate621inter6));
  inv1  gate2512(.a(N1898), .O(gate621inter7));
  inv1  gate2513(.a(N1999), .O(gate621inter8));
  nand2 gate2514(.a(gate621inter8), .b(gate621inter7), .O(gate621inter9));
  nand2 gate2515(.a(s_233), .b(gate621inter3), .O(gate621inter10));
  nor2  gate2516(.a(gate621inter10), .b(gate621inter9), .O(gate621inter11));
  nor2  gate2517(.a(gate621inter11), .b(gate621inter6), .O(gate621inter12));
  nand2 gate2518(.a(gate621inter12), .b(gate621inter1), .O(N2020));
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );

  xor2  gate2771(.a(N2002), .b(N1440), .O(gate624inter0));
  nand2 gate2772(.a(gate624inter0), .b(s_270), .O(gate624inter1));
  and2  gate2773(.a(N2002), .b(N1440), .O(gate624inter2));
  inv1  gate2774(.a(s_270), .O(gate624inter3));
  inv1  gate2775(.a(s_271), .O(gate624inter4));
  nand2 gate2776(.a(gate624inter4), .b(gate624inter3), .O(gate624inter5));
  nor2  gate2777(.a(gate624inter5), .b(gate624inter2), .O(gate624inter6));
  inv1  gate2778(.a(N1440), .O(gate624inter7));
  inv1  gate2779(.a(N2002), .O(gate624inter8));
  nand2 gate2780(.a(gate624inter8), .b(gate624inter7), .O(gate624inter9));
  nand2 gate2781(.a(s_271), .b(gate624inter3), .O(gate624inter10));
  nor2  gate2782(.a(gate624inter10), .b(gate624inter9), .O(gate624inter11));
  nor2  gate2783(.a(gate624inter11), .b(gate624inter6), .O(gate624inter12));
  nand2 gate2784(.a(gate624inter12), .b(gate624inter1), .O(N2023));
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );

  xor2  gate2169(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate2170(.a(gate627inter0), .b(s_184), .O(gate627inter1));
  and2  gate2171(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate2172(.a(s_184), .O(gate627inter3));
  inv1  gate2173(.a(s_185), .O(gate627inter4));
  nand2 gate2174(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate2175(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate2176(.a(N1975), .O(gate627inter7));
  inv1  gate2177(.a(N2008), .O(gate627inter8));
  nand2 gate2178(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate2179(.a(s_185), .b(gate627inter3), .O(gate627inter10));
  nor2  gate2180(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate2181(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate2182(.a(gate627inter12), .b(gate627inter1), .O(N2026));
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );

  xor2  gate2687(.a(N2003), .b(N2023), .O(gate635inter0));
  nand2 gate2688(.a(gate635inter0), .b(s_258), .O(gate635inter1));
  and2  gate2689(.a(N2003), .b(N2023), .O(gate635inter2));
  inv1  gate2690(.a(s_258), .O(gate635inter3));
  inv1  gate2691(.a(s_259), .O(gate635inter4));
  nand2 gate2692(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate2693(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate2694(.a(N2023), .O(gate635inter7));
  inv1  gate2695(.a(N2003), .O(gate635inter8));
  nand2 gate2696(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate2697(.a(s_259), .b(gate635inter3), .O(gate635inter10));
  nor2  gate2698(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate2699(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate2700(.a(gate635inter12), .b(gate635inter1), .O(N2040));
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );

  xor2  gate1833(.a(N2025), .b(N2006), .O(gate637inter0));
  nand2 gate1834(.a(gate637inter0), .b(s_136), .O(gate637inter1));
  and2  gate1835(.a(N2025), .b(N2006), .O(gate637inter2));
  inv1  gate1836(.a(s_136), .O(gate637inter3));
  inv1  gate1837(.a(s_137), .O(gate637inter4));
  nand2 gate1838(.a(gate637inter4), .b(gate637inter3), .O(gate637inter5));
  nor2  gate1839(.a(gate637inter5), .b(gate637inter2), .O(gate637inter6));
  inv1  gate1840(.a(N2006), .O(gate637inter7));
  inv1  gate1841(.a(N2025), .O(gate637inter8));
  nand2 gate1842(.a(gate637inter8), .b(gate637inter7), .O(gate637inter9));
  nand2 gate1843(.a(s_137), .b(gate637inter3), .O(gate637inter10));
  nor2  gate1844(.a(gate637inter10), .b(gate637inter9), .O(gate637inter11));
  nor2  gate1845(.a(gate637inter11), .b(gate637inter6), .O(gate637inter12));
  nand2 gate1846(.a(gate637inter12), .b(gate637inter1), .O(N2042));
inv1 gate638( .a(N2026), .O(N2047) );

  xor2  gate1469(.a(N2014), .b(N2036), .O(gate639inter0));
  nand2 gate1470(.a(gate639inter0), .b(s_84), .O(gate639inter1));
  and2  gate1471(.a(N2014), .b(N2036), .O(gate639inter2));
  inv1  gate1472(.a(s_84), .O(gate639inter3));
  inv1  gate1473(.a(s_85), .O(gate639inter4));
  nand2 gate1474(.a(gate639inter4), .b(gate639inter3), .O(gate639inter5));
  nor2  gate1475(.a(gate639inter5), .b(gate639inter2), .O(gate639inter6));
  inv1  gate1476(.a(N2036), .O(gate639inter7));
  inv1  gate1477(.a(N2014), .O(gate639inter8));
  nand2 gate1478(.a(gate639inter8), .b(gate639inter7), .O(gate639inter9));
  nand2 gate1479(.a(s_85), .b(gate639inter3), .O(gate639inter10));
  nor2  gate1480(.a(gate639inter10), .b(gate639inter9), .O(gate639inter11));
  nor2  gate1481(.a(gate639inter11), .b(gate639inter6), .O(gate639inter12));
  nand2 gate1482(.a(gate639inter12), .b(gate639inter1), .O(N2052));

  xor2  gate2575(.a(N2016), .b(N2037), .O(gate640inter0));
  nand2 gate2576(.a(gate640inter0), .b(s_242), .O(gate640inter1));
  and2  gate2577(.a(N2016), .b(N2037), .O(gate640inter2));
  inv1  gate2578(.a(s_242), .O(gate640inter3));
  inv1  gate2579(.a(s_243), .O(gate640inter4));
  nand2 gate2580(.a(gate640inter4), .b(gate640inter3), .O(gate640inter5));
  nor2  gate2581(.a(gate640inter5), .b(gate640inter2), .O(gate640inter6));
  inv1  gate2582(.a(N2037), .O(gate640inter7));
  inv1  gate2583(.a(N2016), .O(gate640inter8));
  nand2 gate2584(.a(gate640inter8), .b(gate640inter7), .O(gate640inter9));
  nand2 gate2585(.a(s_243), .b(gate640inter3), .O(gate640inter10));
  nor2  gate2586(.a(gate640inter10), .b(gate640inter9), .O(gate640inter11));
  nor2  gate2587(.a(gate640inter11), .b(gate640inter6), .O(gate640inter12));
  nand2 gate2588(.a(gate640inter12), .b(gate640inter1), .O(N2055));
inv1 gate641( .a(N2038), .O(N2060) );

  xor2  gate2449(.a(N2022), .b(N2039), .O(gate642inter0));
  nand2 gate2450(.a(gate642inter0), .b(s_224), .O(gate642inter1));
  and2  gate2451(.a(N2022), .b(N2039), .O(gate642inter2));
  inv1  gate2452(.a(s_224), .O(gate642inter3));
  inv1  gate2453(.a(s_225), .O(gate642inter4));
  nand2 gate2454(.a(gate642inter4), .b(gate642inter3), .O(gate642inter5));
  nor2  gate2455(.a(gate642inter5), .b(gate642inter2), .O(gate642inter6));
  inv1  gate2456(.a(N2039), .O(gate642inter7));
  inv1  gate2457(.a(N2022), .O(gate642inter8));
  nand2 gate2458(.a(gate642inter8), .b(gate642inter7), .O(gate642inter9));
  nand2 gate2459(.a(s_225), .b(gate642inter3), .O(gate642inter10));
  nor2  gate2460(.a(gate642inter10), .b(gate642inter9), .O(gate642inter11));
  nor2  gate2461(.a(gate642inter11), .b(gate642inter6), .O(gate642inter12));
  nand2 gate2462(.a(gate642inter12), .b(gate642inter1), .O(N2061));

  xor2  gate2407(.a(N290), .b(N2040), .O(gate643inter0));
  nand2 gate2408(.a(gate643inter0), .b(s_218), .O(gate643inter1));
  and2  gate2409(.a(N290), .b(N2040), .O(gate643inter2));
  inv1  gate2410(.a(s_218), .O(gate643inter3));
  inv1  gate2411(.a(s_219), .O(gate643inter4));
  nand2 gate2412(.a(gate643inter4), .b(gate643inter3), .O(gate643inter5));
  nor2  gate2413(.a(gate643inter5), .b(gate643inter2), .O(gate643inter6));
  inv1  gate2414(.a(N2040), .O(gate643inter7));
  inv1  gate2415(.a(N290), .O(gate643inter8));
  nand2 gate2416(.a(gate643inter8), .b(gate643inter7), .O(gate643inter9));
  nand2 gate2417(.a(s_219), .b(gate643inter3), .O(gate643inter10));
  nor2  gate2418(.a(gate643inter10), .b(gate643inter9), .O(gate643inter11));
  nor2  gate2419(.a(gate643inter11), .b(gate643inter6), .O(gate643inter12));
  nand2 gate2420(.a(gate643inter12), .b(gate643inter1), .O(N2062));
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate2309(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate2310(.a(gate671inter0), .b(s_204), .O(gate671inter1));
  and2  gate2311(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate2312(.a(s_204), .O(gate671inter3));
  inv1  gate2313(.a(s_205), .O(gate671inter4));
  nand2 gate2314(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate2315(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate2316(.a(N2205), .O(gate671inter7));
  inv1  gate2317(.a(N913), .O(gate671inter8));
  nand2 gate2318(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate2319(.a(s_205), .b(gate671inter3), .O(gate671inter10));
  nor2  gate2320(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate2321(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate2322(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );

  xor2  gate1455(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate1456(.a(gate678inter0), .b(s_82), .O(gate678inter1));
  and2  gate1457(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate1458(.a(s_82), .O(gate678inter3));
  inv1  gate1459(.a(s_83), .O(gate678inter4));
  nand2 gate1460(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate1461(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate1462(.a(N1252), .O(gate678inter7));
  inv1  gate1463(.a(N2225), .O(gate678inter8));
  nand2 gate1464(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate1465(.a(s_83), .b(gate678inter3), .O(gate678inter10));
  nor2  gate1466(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate1467(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate1468(.a(gate678inter12), .b(gate678inter1), .O(N2233));

  xor2  gate1623(.a(N2227), .b(N661), .O(gate679inter0));
  nand2 gate1624(.a(gate679inter0), .b(s_106), .O(gate679inter1));
  and2  gate1625(.a(N2227), .b(N661), .O(gate679inter2));
  inv1  gate1626(.a(s_106), .O(gate679inter3));
  inv1  gate1627(.a(s_107), .O(gate679inter4));
  nand2 gate1628(.a(gate679inter4), .b(gate679inter3), .O(gate679inter5));
  nor2  gate1629(.a(gate679inter5), .b(gate679inter2), .O(gate679inter6));
  inv1  gate1630(.a(N661), .O(gate679inter7));
  inv1  gate1631(.a(N2227), .O(gate679inter8));
  nand2 gate1632(.a(gate679inter8), .b(gate679inter7), .O(gate679inter9));
  nand2 gate1633(.a(s_107), .b(gate679inter3), .O(gate679inter10));
  nor2  gate1634(.a(gate679inter10), .b(gate679inter9), .O(gate679inter11));
  nor2  gate1635(.a(gate679inter11), .b(gate679inter6), .O(gate679inter12));
  nand2 gate1636(.a(gate679inter12), .b(gate679inter1), .O(N2234));
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );

  xor2  gate1581(.a(N2230), .b(N2214), .O(gate681inter0));
  nand2 gate1582(.a(gate681inter0), .b(s_100), .O(gate681inter1));
  and2  gate1583(.a(N2230), .b(N2214), .O(gate681inter2));
  inv1  gate1584(.a(s_100), .O(gate681inter3));
  inv1  gate1585(.a(s_101), .O(gate681inter4));
  nand2 gate1586(.a(gate681inter4), .b(gate681inter3), .O(gate681inter5));
  nor2  gate1587(.a(gate681inter5), .b(gate681inter2), .O(gate681inter6));
  inv1  gate1588(.a(N2214), .O(gate681inter7));
  inv1  gate1589(.a(N2230), .O(gate681inter8));
  nand2 gate1590(.a(gate681inter8), .b(gate681inter7), .O(gate681inter9));
  nand2 gate1591(.a(s_101), .b(gate681inter3), .O(gate681inter10));
  nor2  gate1592(.a(gate681inter10), .b(gate681inter9), .O(gate681inter11));
  nor2  gate1593(.a(gate681inter11), .b(gate681inter6), .O(gate681inter12));
  nand2 gate1594(.a(gate681inter12), .b(gate681inter1), .O(N2236));

  xor2  gate1679(.a(N2231), .b(N2216), .O(gate682inter0));
  nand2 gate1680(.a(gate682inter0), .b(s_114), .O(gate682inter1));
  and2  gate1681(.a(N2231), .b(N2216), .O(gate682inter2));
  inv1  gate1682(.a(s_114), .O(gate682inter3));
  inv1  gate1683(.a(s_115), .O(gate682inter4));
  nand2 gate1684(.a(gate682inter4), .b(gate682inter3), .O(gate682inter5));
  nor2  gate1685(.a(gate682inter5), .b(gate682inter2), .O(gate682inter6));
  inv1  gate1686(.a(N2216), .O(gate682inter7));
  inv1  gate1687(.a(N2231), .O(gate682inter8));
  nand2 gate1688(.a(gate682inter8), .b(gate682inter7), .O(gate682inter9));
  nand2 gate1689(.a(s_115), .b(gate682inter3), .O(gate682inter10));
  nor2  gate1690(.a(gate682inter10), .b(gate682inter9), .O(gate682inter11));
  nor2  gate1691(.a(gate682inter11), .b(gate682inter6), .O(gate682inter12));
  nand2 gate1692(.a(gate682inter12), .b(gate682inter1), .O(N2237));
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );

  xor2  gate2701(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate2702(.a(gate684inter0), .b(s_260), .O(gate684inter1));
  and2  gate2703(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate2704(.a(s_260), .O(gate684inter3));
  inv1  gate2705(.a(s_261), .O(gate684inter4));
  nand2 gate2706(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate2707(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate2708(.a(N2224), .O(gate684inter7));
  inv1  gate2709(.a(N2233), .O(gate684inter8));
  nand2 gate2710(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate2711(.a(s_261), .b(gate684inter3), .O(gate684inter10));
  nor2  gate2712(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate2713(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate2714(.a(gate684inter12), .b(gate684inter1), .O(N2241));
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate1343(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate1344(.a(gate756inter0), .b(s_66), .O(gate756inter1));
  and2  gate1345(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate1346(.a(s_66), .O(gate756inter3));
  inv1  gate1347(.a(s_67), .O(gate756inter4));
  nand2 gate1348(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate1349(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate1350(.a(N2567), .O(gate756inter7));
  inv1  gate1351(.a(N537), .O(gate756inter8));
  nand2 gate1352(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate1353(.a(s_67), .b(gate756inter3), .O(gate756inter10));
  nor2  gate1354(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate1355(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate1356(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );

  xor2  gate1903(.a(N543), .b(N2570), .O(gate758inter0));
  nand2 gate1904(.a(gate758inter0), .b(s_146), .O(gate758inter1));
  and2  gate1905(.a(N543), .b(N2570), .O(gate758inter2));
  inv1  gate1906(.a(s_146), .O(gate758inter3));
  inv1  gate1907(.a(s_147), .O(gate758inter4));
  nand2 gate1908(.a(gate758inter4), .b(gate758inter3), .O(gate758inter5));
  nor2  gate1909(.a(gate758inter5), .b(gate758inter2), .O(gate758inter6));
  inv1  gate1910(.a(N2570), .O(gate758inter7));
  inv1  gate1911(.a(N543), .O(gate758inter8));
  nand2 gate1912(.a(gate758inter8), .b(gate758inter7), .O(gate758inter9));
  nand2 gate1913(.a(s_147), .b(gate758inter3), .O(gate758inter10));
  nor2  gate1914(.a(gate758inter10), .b(gate758inter9), .O(gate758inter11));
  nor2  gate1915(.a(gate758inter11), .b(gate758inter6), .O(gate758inter12));
  nand2 gate1916(.a(gate758inter12), .b(gate758inter1), .O(N2682));
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );

  xor2  gate2085(.a(N549), .b(N2576), .O(gate762inter0));
  nand2 gate2086(.a(gate762inter0), .b(s_172), .O(gate762inter1));
  and2  gate2087(.a(N549), .b(N2576), .O(gate762inter2));
  inv1  gate2088(.a(s_172), .O(gate762inter3));
  inv1  gate2089(.a(s_173), .O(gate762inter4));
  nand2 gate2090(.a(gate762inter4), .b(gate762inter3), .O(gate762inter5));
  nor2  gate2091(.a(gate762inter5), .b(gate762inter2), .O(gate762inter6));
  inv1  gate2092(.a(N2576), .O(gate762inter7));
  inv1  gate2093(.a(N549), .O(gate762inter8));
  nand2 gate2094(.a(gate762inter8), .b(gate762inter7), .O(gate762inter9));
  nand2 gate2095(.a(s_173), .b(gate762inter3), .O(gate762inter10));
  nor2  gate2096(.a(gate762inter10), .b(gate762inter9), .O(gate762inter11));
  nor2  gate2097(.a(gate762inter11), .b(gate762inter6), .O(gate762inter12));
  nand2 gate2098(.a(gate762inter12), .b(gate762inter1), .O(N2690));
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );

  xor2  gate1357(.a(N2672), .b(N346), .O(gate766inter0));
  nand2 gate1358(.a(gate766inter0), .b(s_68), .O(gate766inter1));
  and2  gate1359(.a(N2672), .b(N346), .O(gate766inter2));
  inv1  gate1360(.a(s_68), .O(gate766inter3));
  inv1  gate1361(.a(s_69), .O(gate766inter4));
  nand2 gate1362(.a(gate766inter4), .b(gate766inter3), .O(gate766inter5));
  nor2  gate1363(.a(gate766inter5), .b(gate766inter2), .O(gate766inter6));
  inv1  gate1364(.a(N346), .O(gate766inter7));
  inv1  gate1365(.a(N2672), .O(gate766inter8));
  nand2 gate1366(.a(gate766inter8), .b(gate766inter7), .O(gate766inter9));
  nand2 gate1367(.a(s_69), .b(gate766inter3), .O(gate766inter10));
  nor2  gate1368(.a(gate766inter10), .b(gate766inter9), .O(gate766inter11));
  nor2  gate1369(.a(gate766inter11), .b(gate766inter6), .O(gate766inter12));
  nand2 gate1370(.a(gate766inter12), .b(gate766inter1), .O(N2721));

  xor2  gate1315(.a(N2674), .b(N349), .O(gate767inter0));
  nand2 gate1316(.a(gate767inter0), .b(s_62), .O(gate767inter1));
  and2  gate1317(.a(N2674), .b(N349), .O(gate767inter2));
  inv1  gate1318(.a(s_62), .O(gate767inter3));
  inv1  gate1319(.a(s_63), .O(gate767inter4));
  nand2 gate1320(.a(gate767inter4), .b(gate767inter3), .O(gate767inter5));
  nor2  gate1321(.a(gate767inter5), .b(gate767inter2), .O(gate767inter6));
  inv1  gate1322(.a(N349), .O(gate767inter7));
  inv1  gate1323(.a(N2674), .O(gate767inter8));
  nand2 gate1324(.a(gate767inter8), .b(gate767inter7), .O(gate767inter9));
  nand2 gate1325(.a(s_63), .b(gate767inter3), .O(gate767inter10));
  nor2  gate1326(.a(gate767inter10), .b(gate767inter9), .O(gate767inter11));
  nor2  gate1327(.a(gate767inter11), .b(gate767inter6), .O(gate767inter12));
  nand2 gate1328(.a(gate767inter12), .b(gate767inter1), .O(N2722));

  xor2  gate1399(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate1400(.a(gate768inter0), .b(s_74), .O(gate768inter1));
  and2  gate1401(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate1402(.a(s_74), .O(gate768inter3));
  inv1  gate1403(.a(s_75), .O(gate768inter4));
  nand2 gate1404(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate1405(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate1406(.a(N352), .O(gate768inter7));
  inv1  gate1407(.a(N2676), .O(gate768inter8));
  nand2 gate1408(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate1409(.a(s_75), .b(gate768inter3), .O(gate768inter10));
  nor2  gate1410(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate1411(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate1412(.a(gate768inter12), .b(gate768inter1), .O(N2723));

  xor2  gate1553(.a(N538), .b(N2639), .O(gate769inter0));
  nand2 gate1554(.a(gate769inter0), .b(s_96), .O(gate769inter1));
  and2  gate1555(.a(N538), .b(N2639), .O(gate769inter2));
  inv1  gate1556(.a(s_96), .O(gate769inter3));
  inv1  gate1557(.a(s_97), .O(gate769inter4));
  nand2 gate1558(.a(gate769inter4), .b(gate769inter3), .O(gate769inter5));
  nor2  gate1559(.a(gate769inter5), .b(gate769inter2), .O(gate769inter6));
  inv1  gate1560(.a(N2639), .O(gate769inter7));
  inv1  gate1561(.a(N538), .O(gate769inter8));
  nand2 gate1562(.a(gate769inter8), .b(gate769inter7), .O(gate769inter9));
  nand2 gate1563(.a(s_97), .b(gate769inter3), .O(gate769inter10));
  nor2  gate1564(.a(gate769inter10), .b(gate769inter9), .O(gate769inter11));
  nor2  gate1565(.a(gate769inter11), .b(gate769inter6), .O(gate769inter12));
  nand2 gate1566(.a(gate769inter12), .b(gate769inter1), .O(N2724));
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );

  xor2  gate1371(.a(N541), .b(N2648), .O(gate775inter0));
  nand2 gate1372(.a(gate775inter0), .b(s_70), .O(gate775inter1));
  and2  gate1373(.a(N541), .b(N2648), .O(gate775inter2));
  inv1  gate1374(.a(s_70), .O(gate775inter3));
  inv1  gate1375(.a(s_71), .O(gate775inter4));
  nand2 gate1376(.a(gate775inter4), .b(gate775inter3), .O(gate775inter5));
  nor2  gate1377(.a(gate775inter5), .b(gate775inter2), .O(gate775inter6));
  inv1  gate1378(.a(N2648), .O(gate775inter7));
  inv1  gate1379(.a(N541), .O(gate775inter8));
  nand2 gate1380(.a(gate775inter8), .b(gate775inter7), .O(gate775inter9));
  nand2 gate1381(.a(s_71), .b(gate775inter3), .O(gate775inter10));
  nor2  gate1382(.a(gate775inter10), .b(gate775inter9), .O(gate775inter11));
  nor2  gate1383(.a(gate775inter11), .b(gate775inter6), .O(gate775inter12));
  nand2 gate1384(.a(gate775inter12), .b(gate775inter1), .O(N2730));
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );

  xor2  gate1847(.a(N544), .b(N2655), .O(gate780inter0));
  nand2 gate1848(.a(gate780inter0), .b(s_138), .O(gate780inter1));
  and2  gate1849(.a(N544), .b(N2655), .O(gate780inter2));
  inv1  gate1850(.a(s_138), .O(gate780inter3));
  inv1  gate1851(.a(s_139), .O(gate780inter4));
  nand2 gate1852(.a(gate780inter4), .b(gate780inter3), .O(gate780inter5));
  nor2  gate1853(.a(gate780inter5), .b(gate780inter2), .O(gate780inter6));
  inv1  gate1854(.a(N2655), .O(gate780inter7));
  inv1  gate1855(.a(N544), .O(gate780inter8));
  nand2 gate1856(.a(gate780inter8), .b(gate780inter7), .O(gate780inter9));
  nand2 gate1857(.a(s_139), .b(gate780inter3), .O(gate780inter10));
  nor2  gate1858(.a(gate780inter10), .b(gate780inter9), .O(gate780inter11));
  nor2  gate1859(.a(gate780inter11), .b(gate780inter6), .O(gate780inter12));
  nand2 gate1860(.a(gate780inter12), .b(gate780inter1), .O(N2735));
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );

  xor2  gate1105(.a(N546), .b(N2661), .O(gate784inter0));
  nand2 gate1106(.a(gate784inter0), .b(s_32), .O(gate784inter1));
  and2  gate1107(.a(N546), .b(N2661), .O(gate784inter2));
  inv1  gate1108(.a(s_32), .O(gate784inter3));
  inv1  gate1109(.a(s_33), .O(gate784inter4));
  nand2 gate1110(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate1111(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate1112(.a(N2661), .O(gate784inter7));
  inv1  gate1113(.a(N546), .O(gate784inter8));
  nand2 gate1114(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate1115(.a(s_33), .b(gate784inter3), .O(gate784inter10));
  nor2  gate1116(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate1117(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate1118(.a(gate784inter12), .b(gate784inter1), .O(N2739));
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate1525(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate1526(.a(gate788inter0), .b(s_92), .O(gate788inter1));
  and2  gate1527(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate1528(.a(s_92), .O(gate788inter3));
  inv1  gate1529(.a(s_93), .O(gate788inter4));
  nand2 gate1530(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate1531(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate1532(.a(N385), .O(gate788inter7));
  inv1  gate1533(.a(N2689), .O(gate788inter8));
  nand2 gate1534(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate1535(.a(s_93), .b(gate788inter3), .O(gate788inter10));
  nor2  gate1536(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate1537(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate1538(.a(gate788inter12), .b(gate788inter1), .O(N2743));
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );

  xor2  gate1987(.a(N2722), .b(N2673), .O(gate796inter0));
  nand2 gate1988(.a(gate796inter0), .b(s_158), .O(gate796inter1));
  and2  gate1989(.a(N2722), .b(N2673), .O(gate796inter2));
  inv1  gate1990(.a(s_158), .O(gate796inter3));
  inv1  gate1991(.a(s_159), .O(gate796inter4));
  nand2 gate1992(.a(gate796inter4), .b(gate796inter3), .O(gate796inter5));
  nor2  gate1993(.a(gate796inter5), .b(gate796inter2), .O(gate796inter6));
  inv1  gate1994(.a(N2673), .O(gate796inter7));
  inv1  gate1995(.a(N2722), .O(gate796inter8));
  nand2 gate1996(.a(gate796inter8), .b(gate796inter7), .O(gate796inter9));
  nand2 gate1997(.a(s_159), .b(gate796inter3), .O(gate796inter10));
  nor2  gate1998(.a(gate796inter10), .b(gate796inter9), .O(gate796inter11));
  nor2  gate1999(.a(gate796inter11), .b(gate796inter6), .O(gate796inter12));
  nand2 gate2000(.a(gate796inter12), .b(gate796inter1), .O(N2755));
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );

  xor2  gate2673(.a(N2725), .b(N355), .O(gate798inter0));
  nand2 gate2674(.a(gate798inter0), .b(s_256), .O(gate798inter1));
  and2  gate2675(.a(N2725), .b(N355), .O(gate798inter2));
  inv1  gate2676(.a(s_256), .O(gate798inter3));
  inv1  gate2677(.a(s_257), .O(gate798inter4));
  nand2 gate2678(.a(gate798inter4), .b(gate798inter3), .O(gate798inter5));
  nor2  gate2679(.a(gate798inter5), .b(gate798inter2), .O(gate798inter6));
  inv1  gate2680(.a(N355), .O(gate798inter7));
  inv1  gate2681(.a(N2725), .O(gate798inter8));
  nand2 gate2682(.a(gate798inter8), .b(gate798inter7), .O(gate798inter9));
  nand2 gate2683(.a(s_257), .b(gate798inter3), .O(gate798inter10));
  nor2  gate2684(.a(gate798inter10), .b(gate798inter9), .O(gate798inter11));
  nor2  gate2685(.a(gate798inter11), .b(gate798inter6), .O(gate798inter12));
  nand2 gate2686(.a(gate798inter12), .b(gate798inter1), .O(N2757));
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );

  xor2  gate1133(.a(N2731), .b(N364), .O(gate801inter0));
  nand2 gate1134(.a(gate801inter0), .b(s_36), .O(gate801inter1));
  and2  gate1135(.a(N2731), .b(N364), .O(gate801inter2));
  inv1  gate1136(.a(s_36), .O(gate801inter3));
  inv1  gate1137(.a(s_37), .O(gate801inter4));
  nand2 gate1138(.a(gate801inter4), .b(gate801inter3), .O(gate801inter5));
  nor2  gate1139(.a(gate801inter5), .b(gate801inter2), .O(gate801inter6));
  inv1  gate1140(.a(N364), .O(gate801inter7));
  inv1  gate1141(.a(N2731), .O(gate801inter8));
  nand2 gate1142(.a(gate801inter8), .b(gate801inter7), .O(gate801inter9));
  nand2 gate1143(.a(s_37), .b(gate801inter3), .O(gate801inter10));
  nor2  gate1144(.a(gate801inter10), .b(gate801inter9), .O(gate801inter11));
  nor2  gate1145(.a(gate801inter11), .b(gate801inter6), .O(gate801inter12));
  nand2 gate1146(.a(gate801inter12), .b(gate801inter1), .O(N2760));
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );

  xor2  gate1329(.a(N2738), .b(N376), .O(gate805inter0));
  nand2 gate1330(.a(gate805inter0), .b(s_64), .O(gate805inter1));
  and2  gate1331(.a(N2738), .b(N376), .O(gate805inter2));
  inv1  gate1332(.a(s_64), .O(gate805inter3));
  inv1  gate1333(.a(s_65), .O(gate805inter4));
  nand2 gate1334(.a(gate805inter4), .b(gate805inter3), .O(gate805inter5));
  nor2  gate1335(.a(gate805inter5), .b(gate805inter2), .O(gate805inter6));
  inv1  gate1336(.a(N376), .O(gate805inter7));
  inv1  gate1337(.a(N2738), .O(gate805inter8));
  nand2 gate1338(.a(gate805inter8), .b(gate805inter7), .O(gate805inter9));
  nand2 gate1339(.a(s_65), .b(gate805inter3), .O(gate805inter10));
  nor2  gate1340(.a(gate805inter10), .b(gate805inter9), .O(gate805inter11));
  nor2  gate1341(.a(gate805inter11), .b(gate805inter6), .O(gate805inter12));
  nand2 gate1342(.a(gate805inter12), .b(gate805inter1), .O(N2764));
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );

  xor2  gate1119(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate1120(.a(gate813inter0), .b(s_34), .O(gate813inter1));
  and2  gate1121(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate1122(.a(s_34), .O(gate813inter3));
  inv1  gate1123(.a(s_35), .O(gate813inter4));
  nand2 gate1124(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate1125(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate1126(.a(N2726), .O(gate813inter7));
  inv1  gate1127(.a(N2758), .O(gate813inter8));
  nand2 gate1128(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate1129(.a(s_35), .b(gate813inter3), .O(gate813inter10));
  nor2  gate1130(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate1131(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate1132(.a(gate813inter12), .b(gate813inter1), .O(N2780));

  xor2  gate2547(.a(N2759), .b(N2728), .O(gate814inter0));
  nand2 gate2548(.a(gate814inter0), .b(s_238), .O(gate814inter1));
  and2  gate2549(.a(N2759), .b(N2728), .O(gate814inter2));
  inv1  gate2550(.a(s_238), .O(gate814inter3));
  inv1  gate2551(.a(s_239), .O(gate814inter4));
  nand2 gate2552(.a(gate814inter4), .b(gate814inter3), .O(gate814inter5));
  nor2  gate2553(.a(gate814inter5), .b(gate814inter2), .O(gate814inter6));
  inv1  gate2554(.a(N2728), .O(gate814inter7));
  inv1  gate2555(.a(N2759), .O(gate814inter8));
  nand2 gate2556(.a(gate814inter8), .b(gate814inter7), .O(gate814inter9));
  nand2 gate2557(.a(s_239), .b(gate814inter3), .O(gate814inter10));
  nor2  gate2558(.a(gate814inter10), .b(gate814inter9), .O(gate814inter11));
  nor2  gate2559(.a(gate814inter11), .b(gate814inter6), .O(gate814inter12));
  nand2 gate2560(.a(gate814inter12), .b(gate814inter1), .O(N2781));

  xor2  gate1511(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate1512(.a(gate815inter0), .b(s_90), .O(gate815inter1));
  and2  gate1513(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate1514(.a(s_90), .O(gate815inter3));
  inv1  gate1515(.a(s_91), .O(gate815inter4));
  nand2 gate1516(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate1517(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate1518(.a(N2730), .O(gate815inter7));
  inv1  gate1519(.a(N2760), .O(gate815inter8));
  nand2 gate1520(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate1521(.a(s_91), .b(gate815inter3), .O(gate815inter10));
  nor2  gate1522(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate1523(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate1524(.a(gate815inter12), .b(gate815inter1), .O(N2782));

  xor2  gate993(.a(N2761), .b(N2732), .O(gate816inter0));
  nand2 gate994(.a(gate816inter0), .b(s_16), .O(gate816inter1));
  and2  gate995(.a(N2761), .b(N2732), .O(gate816inter2));
  inv1  gate996(.a(s_16), .O(gate816inter3));
  inv1  gate997(.a(s_17), .O(gate816inter4));
  nand2 gate998(.a(gate816inter4), .b(gate816inter3), .O(gate816inter5));
  nor2  gate999(.a(gate816inter5), .b(gate816inter2), .O(gate816inter6));
  inv1  gate1000(.a(N2732), .O(gate816inter7));
  inv1  gate1001(.a(N2761), .O(gate816inter8));
  nand2 gate1002(.a(gate816inter8), .b(gate816inter7), .O(gate816inter9));
  nand2 gate1003(.a(s_17), .b(gate816inter3), .O(gate816inter10));
  nor2  gate1004(.a(gate816inter10), .b(gate816inter9), .O(gate816inter11));
  nor2  gate1005(.a(gate816inter11), .b(gate816inter6), .O(gate816inter12));
  nand2 gate1006(.a(gate816inter12), .b(gate816inter1), .O(N2783));
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );

  xor2  gate1973(.a(N2764), .b(N2737), .O(gate818inter0));
  nand2 gate1974(.a(gate818inter0), .b(s_156), .O(gate818inter1));
  and2  gate1975(.a(N2764), .b(N2737), .O(gate818inter2));
  inv1  gate1976(.a(s_156), .O(gate818inter3));
  inv1  gate1977(.a(s_157), .O(gate818inter4));
  nand2 gate1978(.a(gate818inter4), .b(gate818inter3), .O(gate818inter5));
  nor2  gate1979(.a(gate818inter5), .b(gate818inter2), .O(gate818inter6));
  inv1  gate1980(.a(N2737), .O(gate818inter7));
  inv1  gate1981(.a(N2764), .O(gate818inter8));
  nand2 gate1982(.a(gate818inter8), .b(gate818inter7), .O(gate818inter9));
  nand2 gate1983(.a(s_157), .b(gate818inter3), .O(gate818inter10));
  nor2  gate1984(.a(gate818inter10), .b(gate818inter9), .O(gate818inter11));
  nor2  gate1985(.a(gate818inter11), .b(gate818inter6), .O(gate818inter12));
  nand2 gate1986(.a(gate818inter12), .b(gate818inter1), .O(N2785));
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );

  xor2  gate1441(.a(N2019), .b(N2776), .O(gate826inter0));
  nand2 gate1442(.a(gate826inter0), .b(s_80), .O(gate826inter1));
  and2  gate1443(.a(N2019), .b(N2776), .O(gate826inter2));
  inv1  gate1444(.a(s_80), .O(gate826inter3));
  inv1  gate1445(.a(s_81), .O(gate826inter4));
  nand2 gate1446(.a(gate826inter4), .b(gate826inter3), .O(gate826inter5));
  nor2  gate1447(.a(gate826inter5), .b(gate826inter2), .O(gate826inter6));
  inv1  gate1448(.a(N2776), .O(gate826inter7));
  inv1  gate1449(.a(N2019), .O(gate826inter8));
  nand2 gate1450(.a(gate826inter8), .b(gate826inter7), .O(gate826inter9));
  nand2 gate1451(.a(s_81), .b(gate826inter3), .O(gate826inter10));
  nor2  gate1452(.a(gate826inter10), .b(gate826inter9), .O(gate826inter11));
  nor2  gate1453(.a(gate826inter11), .b(gate826inter6), .O(gate826inter12));
  nand2 gate1454(.a(gate826inter12), .b(gate826inter1), .O(N2809));
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );

  xor2  gate2211(.a(N2827), .b(N2807), .O(gate837inter0));
  nand2 gate2212(.a(gate837inter0), .b(s_190), .O(gate837inter1));
  and2  gate2213(.a(N2827), .b(N2807), .O(gate837inter2));
  inv1  gate2214(.a(s_190), .O(gate837inter3));
  inv1  gate2215(.a(s_191), .O(gate837inter4));
  nand2 gate2216(.a(gate837inter4), .b(gate837inter3), .O(gate837inter5));
  nor2  gate2217(.a(gate837inter5), .b(gate837inter2), .O(gate837inter6));
  inv1  gate2218(.a(N2807), .O(gate837inter7));
  inv1  gate2219(.a(N2827), .O(gate837inter8));
  nand2 gate2220(.a(gate837inter8), .b(gate837inter7), .O(gate837inter9));
  nand2 gate2221(.a(s_191), .b(gate837inter3), .O(gate837inter10));
  nor2  gate2222(.a(gate837inter10), .b(gate837inter9), .O(gate837inter11));
  nor2  gate2223(.a(gate837inter11), .b(gate837inter6), .O(gate837inter12));
  nand2 gate2224(.a(gate837inter12), .b(gate837inter1), .O(N2843));
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );

  xor2  gate2421(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate2422(.a(gate840inter0), .b(s_220), .O(gate840inter1));
  and2  gate2423(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate2424(.a(s_220), .O(gate840inter3));
  inv1  gate2425(.a(s_221), .O(gate840inter4));
  nand2 gate2426(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate2427(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate2428(.a(N2815), .O(gate840inter7));
  inv1  gate2429(.a(N2077), .O(gate840inter8));
  nand2 gate2430(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate2431(.a(s_221), .b(gate840inter3), .O(gate840inter10));
  nor2  gate2432(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate2433(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate2434(.a(gate840inter12), .b(gate840inter1), .O(N2851));
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );

  xor2  gate2099(.a(N2857), .b(N2052), .O(gate851inter0));
  nand2 gate2100(.a(gate851inter0), .b(s_174), .O(gate851inter1));
  and2  gate2101(.a(N2857), .b(N2052), .O(gate851inter2));
  inv1  gate2102(.a(s_174), .O(gate851inter3));
  inv1  gate2103(.a(s_175), .O(gate851inter4));
  nand2 gate2104(.a(gate851inter4), .b(gate851inter3), .O(gate851inter5));
  nor2  gate2105(.a(gate851inter5), .b(gate851inter2), .O(gate851inter6));
  inv1  gate2106(.a(N2052), .O(gate851inter7));
  inv1  gate2107(.a(N2857), .O(gate851inter8));
  nand2 gate2108(.a(gate851inter8), .b(gate851inter7), .O(gate851inter9));
  nand2 gate2109(.a(s_175), .b(gate851inter3), .O(gate851inter10));
  nor2  gate2110(.a(gate851inter10), .b(gate851inter9), .O(gate851inter11));
  nor2  gate2111(.a(gate851inter11), .b(gate851inter6), .O(gate851inter12));
  nand2 gate2112(.a(gate851inter12), .b(gate851inter1), .O(N2866));

  xor2  gate2365(.a(N2858), .b(N2055), .O(gate852inter0));
  nand2 gate2366(.a(gate852inter0), .b(s_212), .O(gate852inter1));
  and2  gate2367(.a(N2858), .b(N2055), .O(gate852inter2));
  inv1  gate2368(.a(s_212), .O(gate852inter3));
  inv1  gate2369(.a(s_213), .O(gate852inter4));
  nand2 gate2370(.a(gate852inter4), .b(gate852inter3), .O(gate852inter5));
  nor2  gate2371(.a(gate852inter5), .b(gate852inter2), .O(gate852inter6));
  inv1  gate2372(.a(N2055), .O(gate852inter7));
  inv1  gate2373(.a(N2858), .O(gate852inter8));
  nand2 gate2374(.a(gate852inter8), .b(gate852inter7), .O(gate852inter9));
  nand2 gate2375(.a(s_213), .b(gate852inter3), .O(gate852inter10));
  nor2  gate2376(.a(gate852inter10), .b(gate852inter9), .O(gate852inter11));
  nor2  gate2377(.a(gate852inter11), .b(gate852inter6), .O(gate852inter12));
  nand2 gate2378(.a(gate852inter12), .b(gate852inter1), .O(N2867));

  xor2  gate881(.a(N2859), .b(N1866), .O(gate853inter0));
  nand2 gate882(.a(gate853inter0), .b(s_0), .O(gate853inter1));
  and2  gate883(.a(N2859), .b(N1866), .O(gate853inter2));
  inv1  gate884(.a(s_0), .O(gate853inter3));
  inv1  gate885(.a(s_1), .O(gate853inter4));
  nand2 gate886(.a(gate853inter4), .b(gate853inter3), .O(gate853inter5));
  nor2  gate887(.a(gate853inter5), .b(gate853inter2), .O(gate853inter6));
  inv1  gate888(.a(N1866), .O(gate853inter7));
  inv1  gate889(.a(N2859), .O(gate853inter8));
  nand2 gate890(.a(gate853inter8), .b(gate853inter7), .O(gate853inter9));
  nand2 gate891(.a(s_1), .b(gate853inter3), .O(gate853inter10));
  nor2  gate892(.a(gate853inter10), .b(gate853inter9), .O(gate853inter11));
  nor2  gate893(.a(gate853inter11), .b(gate853inter6), .O(gate853inter12));
  nand2 gate894(.a(gate853inter12), .b(gate853inter1), .O(N2868));

  xor2  gate2729(.a(N2860), .b(N1818), .O(gate854inter0));
  nand2 gate2730(.a(gate854inter0), .b(s_264), .O(gate854inter1));
  and2  gate2731(.a(N2860), .b(N1818), .O(gate854inter2));
  inv1  gate2732(.a(s_264), .O(gate854inter3));
  inv1  gate2733(.a(s_265), .O(gate854inter4));
  nand2 gate2734(.a(gate854inter4), .b(gate854inter3), .O(gate854inter5));
  nor2  gate2735(.a(gate854inter5), .b(gate854inter2), .O(gate854inter6));
  inv1  gate2736(.a(N1818), .O(gate854inter7));
  inv1  gate2737(.a(N2860), .O(gate854inter8));
  nand2 gate2738(.a(gate854inter8), .b(gate854inter7), .O(gate854inter9));
  nand2 gate2739(.a(s_265), .b(gate854inter3), .O(gate854inter10));
  nor2  gate2740(.a(gate854inter10), .b(gate854inter9), .O(gate854inter11));
  nor2  gate2741(.a(gate854inter11), .b(gate854inter6), .O(gate854inter12));
  nand2 gate2742(.a(gate854inter12), .b(gate854inter1), .O(N2869));

  xor2  gate2463(.a(N2861), .b(N1902), .O(gate855inter0));
  nand2 gate2464(.a(gate855inter0), .b(s_226), .O(gate855inter1));
  and2  gate2465(.a(N2861), .b(N1902), .O(gate855inter2));
  inv1  gate2466(.a(s_226), .O(gate855inter3));
  inv1  gate2467(.a(s_227), .O(gate855inter4));
  nand2 gate2468(.a(gate855inter4), .b(gate855inter3), .O(gate855inter5));
  nor2  gate2469(.a(gate855inter5), .b(gate855inter2), .O(gate855inter6));
  inv1  gate2470(.a(N1902), .O(gate855inter7));
  inv1  gate2471(.a(N2861), .O(gate855inter8));
  nand2 gate2472(.a(gate855inter8), .b(gate855inter7), .O(gate855inter9));
  nand2 gate2473(.a(s_227), .b(gate855inter3), .O(gate855inter10));
  nor2  gate2474(.a(gate855inter10), .b(gate855inter9), .O(gate855inter11));
  nor2  gate2475(.a(gate855inter11), .b(gate855inter6), .O(gate855inter12));
  nand2 gate2476(.a(gate855inter12), .b(gate855inter1), .O(N2870));
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate2057(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate2058(.a(gate860inter0), .b(s_168), .O(gate860inter1));
  and2  gate2059(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate2060(.a(s_168), .O(gate860inter3));
  inv1  gate2061(.a(s_169), .O(gate860inter4));
  nand2 gate2062(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate2063(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate2064(.a(N1933), .O(gate860inter7));
  inv1  gate2065(.a(N2862), .O(gate860inter8));
  nand2 gate2066(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate2067(.a(s_169), .b(gate860inter3), .O(gate860inter10));
  nor2  gate2068(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate2069(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate2070(.a(gate860inter12), .b(gate860inter1), .O(N2875));
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );

  xor2  gate1959(.a(N2852), .b(N2868), .O(gate863inter0));
  nand2 gate1960(.a(gate863inter0), .b(s_154), .O(gate863inter1));
  and2  gate1961(.a(N2852), .b(N2868), .O(gate863inter2));
  inv1  gate1962(.a(s_154), .O(gate863inter3));
  inv1  gate1963(.a(s_155), .O(gate863inter4));
  nand2 gate1964(.a(gate863inter4), .b(gate863inter3), .O(gate863inter5));
  nor2  gate1965(.a(gate863inter5), .b(gate863inter2), .O(gate863inter6));
  inv1  gate1966(.a(N2868), .O(gate863inter7));
  inv1  gate1967(.a(N2852), .O(gate863inter8));
  nand2 gate1968(.a(gate863inter8), .b(gate863inter7), .O(gate863inter9));
  nand2 gate1969(.a(s_155), .b(gate863inter3), .O(gate863inter10));
  nor2  gate1970(.a(gate863inter10), .b(gate863inter9), .O(gate863inter11));
  nor2  gate1971(.a(gate863inter11), .b(gate863inter6), .O(gate863inter12));
  nand2 gate1972(.a(gate863inter12), .b(gate863inter1), .O(N2878));

  xor2  gate2323(.a(N2853), .b(N2869), .O(gate864inter0));
  nand2 gate2324(.a(gate864inter0), .b(s_206), .O(gate864inter1));
  and2  gate2325(.a(N2853), .b(N2869), .O(gate864inter2));
  inv1  gate2326(.a(s_206), .O(gate864inter3));
  inv1  gate2327(.a(s_207), .O(gate864inter4));
  nand2 gate2328(.a(gate864inter4), .b(gate864inter3), .O(gate864inter5));
  nor2  gate2329(.a(gate864inter5), .b(gate864inter2), .O(gate864inter6));
  inv1  gate2330(.a(N2869), .O(gate864inter7));
  inv1  gate2331(.a(N2853), .O(gate864inter8));
  nand2 gate2332(.a(gate864inter8), .b(gate864inter7), .O(gate864inter9));
  nand2 gate2333(.a(s_207), .b(gate864inter3), .O(gate864inter10));
  nor2  gate2334(.a(gate864inter10), .b(gate864inter9), .O(gate864inter11));
  nor2  gate2335(.a(gate864inter11), .b(gate864inter6), .O(gate864inter12));
  nand2 gate2336(.a(gate864inter12), .b(gate864inter1), .O(N2879));

  xor2  gate1413(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate1414(.a(gate865inter0), .b(s_76), .O(gate865inter1));
  and2  gate1415(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate1416(.a(s_76), .O(gate865inter3));
  inv1  gate1417(.a(s_77), .O(gate865inter4));
  nand2 gate1418(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate1419(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate1420(.a(N2870), .O(gate865inter7));
  inv1  gate1421(.a(N2854), .O(gate865inter8));
  nand2 gate1422(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate1423(.a(s_77), .b(gate865inter3), .O(gate865inter10));
  nor2  gate1424(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate1425(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate1426(.a(gate865inter12), .b(gate865inter1), .O(N2880));

  xor2  gate979(.a(N2872), .b(N682), .O(gate866inter0));
  nand2 gate980(.a(gate866inter0), .b(s_14), .O(gate866inter1));
  and2  gate981(.a(N2872), .b(N682), .O(gate866inter2));
  inv1  gate982(.a(s_14), .O(gate866inter3));
  inv1  gate983(.a(s_15), .O(gate866inter4));
  nand2 gate984(.a(gate866inter4), .b(gate866inter3), .O(gate866inter5));
  nor2  gate985(.a(gate866inter5), .b(gate866inter2), .O(gate866inter6));
  inv1  gate986(.a(N682), .O(gate866inter7));
  inv1  gate987(.a(N2872), .O(gate866inter8));
  nand2 gate988(.a(gate866inter8), .b(gate866inter7), .O(gate866inter9));
  nand2 gate989(.a(s_15), .b(gate866inter3), .O(gate866inter10));
  nor2  gate990(.a(gate866inter10), .b(gate866inter9), .O(gate866inter11));
  nor2  gate991(.a(gate866inter11), .b(gate866inter6), .O(gate866inter12));
  nand2 gate992(.a(gate866inter12), .b(gate866inter1), .O(N2881));
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );

  xor2  gate1651(.a(N2897), .b(N2895), .O(gate879inter0));
  nand2 gate1652(.a(gate879inter0), .b(s_110), .O(gate879inter1));
  and2  gate1653(.a(N2897), .b(N2895), .O(gate879inter2));
  inv1  gate1654(.a(s_110), .O(gate879inter3));
  inv1  gate1655(.a(s_111), .O(gate879inter4));
  nand2 gate1656(.a(gate879inter4), .b(gate879inter3), .O(gate879inter5));
  nor2  gate1657(.a(gate879inter5), .b(gate879inter2), .O(gate879inter6));
  inv1  gate1658(.a(N2895), .O(gate879inter7));
  inv1  gate1659(.a(N2897), .O(gate879inter8));
  nand2 gate1660(.a(gate879inter8), .b(gate879inter7), .O(gate879inter9));
  nand2 gate1661(.a(s_111), .b(gate879inter3), .O(gate879inter10));
  nor2  gate1662(.a(gate879inter10), .b(gate879inter9), .O(gate879inter11));
  nor2  gate1663(.a(gate879inter11), .b(gate879inter6), .O(gate879inter12));
  nand2 gate1664(.a(gate879inter12), .b(gate879inter1), .O(N2898));
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule