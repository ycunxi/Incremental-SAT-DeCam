module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate7inter0, gate7inter1, gate7inter2, gate7inter3, gate7inter4, gate7inter5, gate7inter6, gate7inter7, gate7inter8, gate7inter9, gate7inter10, gate7inter11, gate7inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12;


  xor2  gate329(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate330(.a(gate1inter0), .b(s_18), .O(gate1inter1));
  and2  gate331(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate332(.a(s_18), .O(gate1inter3));
  inv1  gate333(.a(s_19), .O(gate1inter4));
  nand2 gate334(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate335(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate336(.a(N1), .O(gate1inter7));
  inv1  gate337(.a(N5), .O(gate1inter8));
  nand2 gate338(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate339(.a(s_19), .b(gate1inter3), .O(gate1inter10));
  nor2  gate340(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate341(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate342(.a(gate1inter12), .b(gate1inter1), .O(N250));
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate749(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate750(.a(gate4inter0), .b(s_78), .O(gate4inter1));
  and2  gate751(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate752(.a(s_78), .O(gate4inter3));
  inv1  gate753(.a(s_79), .O(gate4inter4));
  nand2 gate754(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate755(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate756(.a(N25), .O(gate4inter7));
  inv1  gate757(.a(N29), .O(gate4inter8));
  nand2 gate758(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate759(.a(s_79), .b(gate4inter3), .O(gate4inter10));
  nor2  gate760(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate761(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate762(.a(gate4inter12), .b(gate4inter1), .O(N253));

  xor2  gate427(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate428(.a(gate5inter0), .b(s_32), .O(gate5inter1));
  and2  gate429(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate430(.a(s_32), .O(gate5inter3));
  inv1  gate431(.a(s_33), .O(gate5inter4));
  nand2 gate432(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate433(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate434(.a(N33), .O(gate5inter7));
  inv1  gate435(.a(N37), .O(gate5inter8));
  nand2 gate436(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate437(.a(s_33), .b(gate5inter3), .O(gate5inter10));
  nor2  gate438(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate439(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate440(.a(gate5inter12), .b(gate5inter1), .O(N254));
xor2 gate6( .a(N41), .b(N45), .O(N255) );

  xor2  gate637(.a(N53), .b(N49), .O(gate7inter0));
  nand2 gate638(.a(gate7inter0), .b(s_62), .O(gate7inter1));
  and2  gate639(.a(N53), .b(N49), .O(gate7inter2));
  inv1  gate640(.a(s_62), .O(gate7inter3));
  inv1  gate641(.a(s_63), .O(gate7inter4));
  nand2 gate642(.a(gate7inter4), .b(gate7inter3), .O(gate7inter5));
  nor2  gate643(.a(gate7inter5), .b(gate7inter2), .O(gate7inter6));
  inv1  gate644(.a(N49), .O(gate7inter7));
  inv1  gate645(.a(N53), .O(gate7inter8));
  nand2 gate646(.a(gate7inter8), .b(gate7inter7), .O(gate7inter9));
  nand2 gate647(.a(s_63), .b(gate7inter3), .O(gate7inter10));
  nor2  gate648(.a(gate7inter10), .b(gate7inter9), .O(gate7inter11));
  nor2  gate649(.a(gate7inter11), .b(gate7inter6), .O(gate7inter12));
  nand2 gate650(.a(gate7inter12), .b(gate7inter1), .O(N256));
xor2 gate8( .a(N57), .b(N61), .O(N257) );

  xor2  gate735(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate736(.a(gate9inter0), .b(s_76), .O(gate9inter1));
  and2  gate737(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate738(.a(s_76), .O(gate9inter3));
  inv1  gate739(.a(s_77), .O(gate9inter4));
  nand2 gate740(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate741(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate742(.a(N65), .O(gate9inter7));
  inv1  gate743(.a(N69), .O(gate9inter8));
  nand2 gate744(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate745(.a(s_77), .b(gate9inter3), .O(gate9inter10));
  nor2  gate746(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate747(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate748(.a(gate9inter12), .b(gate9inter1), .O(N258));

  xor2  gate231(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate232(.a(gate10inter0), .b(s_4), .O(gate10inter1));
  and2  gate233(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate234(.a(s_4), .O(gate10inter3));
  inv1  gate235(.a(s_5), .O(gate10inter4));
  nand2 gate236(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate237(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate238(.a(N73), .O(gate10inter7));
  inv1  gate239(.a(N77), .O(gate10inter8));
  nand2 gate240(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate241(.a(s_5), .b(gate10inter3), .O(gate10inter10));
  nor2  gate242(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate243(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate244(.a(gate10inter12), .b(gate10inter1), .O(N259));
xor2 gate11( .a(N81), .b(N85), .O(N260) );

  xor2  gate217(.a(N93), .b(N89), .O(gate12inter0));
  nand2 gate218(.a(gate12inter0), .b(s_2), .O(gate12inter1));
  and2  gate219(.a(N93), .b(N89), .O(gate12inter2));
  inv1  gate220(.a(s_2), .O(gate12inter3));
  inv1  gate221(.a(s_3), .O(gate12inter4));
  nand2 gate222(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate223(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate224(.a(N89), .O(gate12inter7));
  inv1  gate225(.a(N93), .O(gate12inter8));
  nand2 gate226(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate227(.a(s_3), .b(gate12inter3), .O(gate12inter10));
  nor2  gate228(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate229(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate230(.a(gate12inter12), .b(gate12inter1), .O(N261));

  xor2  gate315(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate316(.a(gate13inter0), .b(s_16), .O(gate13inter1));
  and2  gate317(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate318(.a(s_16), .O(gate13inter3));
  inv1  gate319(.a(s_17), .O(gate13inter4));
  nand2 gate320(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate321(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate322(.a(N97), .O(gate13inter7));
  inv1  gate323(.a(N101), .O(gate13inter8));
  nand2 gate324(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate325(.a(s_17), .b(gate13inter3), .O(gate13inter10));
  nor2  gate326(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate327(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate328(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );

  xor2  gate441(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate442(.a(gate32inter0), .b(s_34), .O(gate32inter1));
  and2  gate443(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate444(.a(s_34), .O(gate32inter3));
  inv1  gate445(.a(s_35), .O(gate32inter4));
  nand2 gate446(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate447(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate448(.a(N45), .O(gate32inter7));
  inv1  gate449(.a(N61), .O(gate32inter8));
  nand2 gate450(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate451(.a(s_35), .b(gate32inter3), .O(gate32inter10));
  nor2  gate452(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate453(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate454(.a(gate32inter12), .b(gate32inter1), .O(N281));

  xor2  gate763(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate764(.a(gate33inter0), .b(s_80), .O(gate33inter1));
  and2  gate765(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate766(.a(s_80), .O(gate33inter3));
  inv1  gate767(.a(s_81), .O(gate33inter4));
  nand2 gate768(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate769(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate770(.a(N65), .O(gate33inter7));
  inv1  gate771(.a(N81), .O(gate33inter8));
  nand2 gate772(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate773(.a(s_81), .b(gate33inter3), .O(gate33inter10));
  nor2  gate774(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate775(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate776(.a(gate33inter12), .b(gate33inter1), .O(N282));
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );

  xor2  gate497(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate498(.a(gate38inter0), .b(s_42), .O(gate38inter1));
  and2  gate499(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate500(.a(s_42), .O(gate38inter3));
  inv1  gate501(.a(s_43), .O(gate38inter4));
  nand2 gate502(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate503(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate504(.a(N105), .O(gate38inter7));
  inv1  gate505(.a(N121), .O(gate38inter8));
  nand2 gate506(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate507(.a(s_43), .b(gate38inter3), .O(gate38inter10));
  nor2  gate508(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate509(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate510(.a(gate38inter12), .b(gate38inter1), .O(N287));
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate343(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate344(.a(gate42inter0), .b(s_20), .O(gate42inter1));
  and2  gate345(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate346(.a(s_20), .O(gate42inter3));
  inv1  gate347(.a(s_21), .O(gate42inter4));
  nand2 gate348(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate349(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate350(.a(N252), .O(gate42inter7));
  inv1  gate351(.a(N253), .O(gate42inter8));
  nand2 gate352(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate353(.a(s_21), .b(gate42inter3), .O(gate42inter10));
  nor2  gate354(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate355(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate356(.a(gate42inter12), .b(gate42inter1), .O(N293));

  xor2  gate623(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate624(.a(gate43inter0), .b(s_60), .O(gate43inter1));
  and2  gate625(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate626(.a(s_60), .O(gate43inter3));
  inv1  gate627(.a(s_61), .O(gate43inter4));
  nand2 gate628(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate629(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate630(.a(N254), .O(gate43inter7));
  inv1  gate631(.a(N255), .O(gate43inter8));
  nand2 gate632(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate633(.a(s_61), .b(gate43inter3), .O(gate43inter10));
  nor2  gate634(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate635(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate636(.a(gate43inter12), .b(gate43inter1), .O(N296));

  xor2  gate413(.a(N257), .b(N256), .O(gate44inter0));
  nand2 gate414(.a(gate44inter0), .b(s_30), .O(gate44inter1));
  and2  gate415(.a(N257), .b(N256), .O(gate44inter2));
  inv1  gate416(.a(s_30), .O(gate44inter3));
  inv1  gate417(.a(s_31), .O(gate44inter4));
  nand2 gate418(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate419(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate420(.a(N256), .O(gate44inter7));
  inv1  gate421(.a(N257), .O(gate44inter8));
  nand2 gate422(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate423(.a(s_31), .b(gate44inter3), .O(gate44inter10));
  nor2  gate424(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate425(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate426(.a(gate44inter12), .b(gate44inter1), .O(N299));

  xor2  gate371(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate372(.a(gate45inter0), .b(s_24), .O(gate45inter1));
  and2  gate373(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate374(.a(s_24), .O(gate45inter3));
  inv1  gate375(.a(s_25), .O(gate45inter4));
  nand2 gate376(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate377(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate378(.a(N258), .O(gate45inter7));
  inv1  gate379(.a(N259), .O(gate45inter8));
  nand2 gate380(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate381(.a(s_25), .b(gate45inter3), .O(gate45inter10));
  nor2  gate382(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate383(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate384(.a(gate45inter12), .b(gate45inter1), .O(N302));
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );

  xor2  gate693(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate694(.a(gate54inter0), .b(s_70), .O(gate54inter1));
  and2  gate695(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate696(.a(s_70), .O(gate54inter3));
  inv1  gate697(.a(s_71), .O(gate54inter4));
  nand2 gate698(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate699(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate700(.a(N284), .O(gate54inter7));
  inv1  gate701(.a(N285), .O(gate54inter8));
  nand2 gate702(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate703(.a(s_71), .b(gate54inter3), .O(gate54inter10));
  nor2  gate704(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate705(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate706(.a(gate54inter12), .b(gate54inter1), .O(N319));
xor2 gate55( .a(N286), .b(N287), .O(N320) );

  xor2  gate399(.a(N289), .b(N288), .O(gate56inter0));
  nand2 gate400(.a(gate56inter0), .b(s_28), .O(gate56inter1));
  and2  gate401(.a(N289), .b(N288), .O(gate56inter2));
  inv1  gate402(.a(s_28), .O(gate56inter3));
  inv1  gate403(.a(s_29), .O(gate56inter4));
  nand2 gate404(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate405(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate406(.a(N288), .O(gate56inter7));
  inv1  gate407(.a(N289), .O(gate56inter8));
  nand2 gate408(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate409(.a(s_29), .b(gate56inter3), .O(gate56inter10));
  nor2  gate410(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate411(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate412(.a(gate56inter12), .b(gate56inter1), .O(N321));

  xor2  gate203(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate204(.a(gate57inter0), .b(s_0), .O(gate57inter1));
  and2  gate205(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate206(.a(s_0), .O(gate57inter3));
  inv1  gate207(.a(s_1), .O(gate57inter4));
  nand2 gate208(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate209(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate210(.a(N290), .O(gate57inter7));
  inv1  gate211(.a(N293), .O(gate57inter8));
  nand2 gate212(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate213(.a(s_1), .b(gate57inter3), .O(gate57inter10));
  nor2  gate214(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate215(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate216(.a(gate57inter12), .b(gate57inter1), .O(N338));

  xor2  gate553(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate554(.a(gate58inter0), .b(s_50), .O(gate58inter1));
  and2  gate555(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate556(.a(s_50), .O(gate58inter3));
  inv1  gate557(.a(s_51), .O(gate58inter4));
  nand2 gate558(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate559(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate560(.a(N296), .O(gate58inter7));
  inv1  gate561(.a(N299), .O(gate58inter8));
  nand2 gate562(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate563(.a(s_51), .b(gate58inter3), .O(gate58inter10));
  nor2  gate564(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate565(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate566(.a(gate58inter12), .b(gate58inter1), .O(N339));

  xor2  gate567(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate568(.a(gate59inter0), .b(s_52), .O(gate59inter1));
  and2  gate569(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate570(.a(s_52), .O(gate59inter3));
  inv1  gate571(.a(s_53), .O(gate59inter4));
  nand2 gate572(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate573(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate574(.a(N290), .O(gate59inter7));
  inv1  gate575(.a(N296), .O(gate59inter8));
  nand2 gate576(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate577(.a(s_53), .b(gate59inter3), .O(gate59inter10));
  nor2  gate578(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate579(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate580(.a(gate59inter12), .b(gate59inter1), .O(N340));

  xor2  gate651(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate652(.a(gate60inter0), .b(s_64), .O(gate60inter1));
  and2  gate653(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate654(.a(s_64), .O(gate60inter3));
  inv1  gate655(.a(s_65), .O(gate60inter4));
  nand2 gate656(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate657(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate658(.a(N293), .O(gate60inter7));
  inv1  gate659(.a(N299), .O(gate60inter8));
  nand2 gate660(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate661(.a(s_65), .b(gate60inter3), .O(gate60inter10));
  nor2  gate662(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate663(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate664(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );

  xor2  gate301(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate302(.a(gate63inter0), .b(s_14), .O(gate63inter1));
  and2  gate303(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate304(.a(s_14), .O(gate63inter3));
  inv1  gate305(.a(s_15), .O(gate63inter4));
  nand2 gate306(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate307(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate308(.a(N302), .O(gate63inter7));
  inv1  gate309(.a(N308), .O(gate63inter8));
  nand2 gate310(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate311(.a(s_15), .b(gate63inter3), .O(gate63inter10));
  nor2  gate312(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate313(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate314(.a(gate63inter12), .b(gate63inter1), .O(N344));

  xor2  gate539(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate540(.a(gate64inter0), .b(s_48), .O(gate64inter1));
  and2  gate541(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate542(.a(s_48), .O(gate64inter3));
  inv1  gate543(.a(s_49), .O(gate64inter4));
  nand2 gate544(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate545(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate546(.a(N305), .O(gate64inter7));
  inv1  gate547(.a(N311), .O(gate64inter8));
  nand2 gate548(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate549(.a(s_49), .b(gate64inter3), .O(gate64inter10));
  nor2  gate550(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate551(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate552(.a(gate64inter12), .b(gate64inter1), .O(N345));
xor2 gate65( .a(N266), .b(N342), .O(N346) );

  xor2  gate483(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate484(.a(gate66inter0), .b(s_40), .O(gate66inter1));
  and2  gate485(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate486(.a(s_40), .O(gate66inter3));
  inv1  gate487(.a(s_41), .O(gate66inter4));
  nand2 gate488(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate489(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate490(.a(N267), .O(gate66inter7));
  inv1  gate491(.a(N343), .O(gate66inter8));
  nand2 gate492(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate493(.a(s_41), .b(gate66inter3), .O(gate66inter10));
  nor2  gate494(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate495(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate496(.a(gate66inter12), .b(gate66inter1), .O(N347));

  xor2  gate609(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate610(.a(gate67inter0), .b(s_58), .O(gate67inter1));
  and2  gate611(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate612(.a(s_58), .O(gate67inter3));
  inv1  gate613(.a(s_59), .O(gate67inter4));
  nand2 gate614(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate615(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate616(.a(N268), .O(gate67inter7));
  inv1  gate617(.a(N344), .O(gate67inter8));
  nand2 gate618(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate619(.a(s_59), .b(gate67inter3), .O(gate67inter10));
  nor2  gate620(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate621(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate622(.a(gate67inter12), .b(gate67inter1), .O(N348));
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );

  xor2  gate595(.a(N341), .b(N273), .O(gate72inter0));
  nand2 gate596(.a(gate72inter0), .b(s_56), .O(gate72inter1));
  and2  gate597(.a(N341), .b(N273), .O(gate72inter2));
  inv1  gate598(.a(s_56), .O(gate72inter3));
  inv1  gate599(.a(s_57), .O(gate72inter4));
  nand2 gate600(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate601(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate602(.a(N273), .O(gate72inter7));
  inv1  gate603(.a(N341), .O(gate72inter8));
  nand2 gate604(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate605(.a(s_57), .b(gate72inter3), .O(gate72inter10));
  nor2  gate606(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate607(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate608(.a(gate72inter12), .b(gate72inter1), .O(N353));
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate511(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate512(.a(gate75inter0), .b(s_44), .O(gate75inter1));
  and2  gate513(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate514(.a(s_44), .O(gate75inter3));
  inv1  gate515(.a(s_45), .O(gate75inter4));
  nand2 gate516(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate517(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate518(.a(N316), .O(gate75inter7));
  inv1  gate519(.a(N348), .O(gate75inter8));
  nand2 gate520(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate521(.a(s_45), .b(gate75inter3), .O(gate75inter10));
  nor2  gate522(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate523(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate524(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate287(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate288(.a(gate80inter0), .b(s_12), .O(gate80inter1));
  and2  gate289(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate290(.a(s_12), .O(gate80inter3));
  inv1  gate291(.a(s_13), .O(gate80inter4));
  nand2 gate292(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate293(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate294(.a(N321), .O(gate80inter7));
  inv1  gate295(.a(N353), .O(gate80inter8));
  nand2 gate296(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate297(.a(s_13), .b(gate80inter3), .O(gate80inter10));
  nor2  gate298(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate299(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate300(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );

  xor2  gate707(.a(N695), .b(N13), .O(gate174inter0));
  nand2 gate708(.a(gate174inter0), .b(s_72), .O(gate174inter1));
  and2  gate709(.a(N695), .b(N13), .O(gate174inter2));
  inv1  gate710(.a(s_72), .O(gate174inter3));
  inv1  gate711(.a(s_73), .O(gate174inter4));
  nand2 gate712(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate713(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate714(.a(N13), .O(gate174inter7));
  inv1  gate715(.a(N695), .O(gate174inter8));
  nand2 gate716(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate717(.a(s_73), .b(gate174inter3), .O(gate174inter10));
  nor2  gate718(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate719(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate720(.a(gate174inter12), .b(gate174inter1), .O(N727));
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );

  xor2  gate525(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate526(.a(gate179inter0), .b(s_46), .O(gate179inter1));
  and2  gate527(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate528(.a(s_46), .O(gate179inter3));
  inv1  gate529(.a(s_47), .O(gate179inter4));
  nand2 gate530(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate531(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate532(.a(N33), .O(gate179inter7));
  inv1  gate533(.a(N700), .O(gate179inter8));
  nand2 gate534(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate535(.a(s_47), .b(gate179inter3), .O(gate179inter10));
  nor2  gate536(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate537(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate538(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );

  xor2  gate357(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate358(.a(gate181inter0), .b(s_22), .O(gate181inter1));
  and2  gate359(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate360(.a(s_22), .O(gate181inter3));
  inv1  gate361(.a(s_23), .O(gate181inter4));
  nand2 gate362(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate363(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate364(.a(N41), .O(gate181inter7));
  inv1  gate365(.a(N702), .O(gate181inter8));
  nand2 gate366(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate367(.a(s_23), .b(gate181inter3), .O(gate181inter10));
  nor2  gate368(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate369(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate370(.a(gate181inter12), .b(gate181inter1), .O(N734));

  xor2  gate385(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate386(.a(gate182inter0), .b(s_26), .O(gate182inter1));
  and2  gate387(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate388(.a(s_26), .O(gate182inter3));
  inv1  gate389(.a(s_27), .O(gate182inter4));
  nand2 gate390(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate391(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate392(.a(N45), .O(gate182inter7));
  inv1  gate393(.a(N703), .O(gate182inter8));
  nand2 gate394(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate395(.a(s_27), .b(gate182inter3), .O(gate182inter10));
  nor2  gate396(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate397(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate398(.a(gate182inter12), .b(gate182inter1), .O(N735));
xor2 gate183( .a(N49), .b(N704), .O(N736) );

  xor2  gate245(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate246(.a(gate184inter0), .b(s_6), .O(gate184inter1));
  and2  gate247(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate248(.a(s_6), .O(gate184inter3));
  inv1  gate249(.a(s_7), .O(gate184inter4));
  nand2 gate250(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate251(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate252(.a(N53), .O(gate184inter7));
  inv1  gate253(.a(N705), .O(gate184inter8));
  nand2 gate254(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate255(.a(s_7), .b(gate184inter3), .O(gate184inter10));
  nor2  gate256(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate257(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate258(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate469(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate470(.a(gate186inter0), .b(s_38), .O(gate186inter1));
  and2  gate471(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate472(.a(s_38), .O(gate186inter3));
  inv1  gate473(.a(s_39), .O(gate186inter4));
  nand2 gate474(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate475(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate476(.a(N61), .O(gate186inter7));
  inv1  gate477(.a(N707), .O(gate186inter8));
  nand2 gate478(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate479(.a(s_39), .b(gate186inter3), .O(gate186inter10));
  nor2  gate480(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate481(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate482(.a(gate186inter12), .b(gate186inter1), .O(N739));

  xor2  gate721(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate722(.a(gate187inter0), .b(s_74), .O(gate187inter1));
  and2  gate723(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate724(.a(s_74), .O(gate187inter3));
  inv1  gate725(.a(s_75), .O(gate187inter4));
  nand2 gate726(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate727(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate728(.a(N65), .O(gate187inter7));
  inv1  gate729(.a(N708), .O(gate187inter8));
  nand2 gate730(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate731(.a(s_75), .b(gate187inter3), .O(gate187inter10));
  nor2  gate732(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate733(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate734(.a(gate187inter12), .b(gate187inter1), .O(N740));

  xor2  gate273(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate274(.a(gate188inter0), .b(s_10), .O(gate188inter1));
  and2  gate275(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate276(.a(s_10), .O(gate188inter3));
  inv1  gate277(.a(s_11), .O(gate188inter4));
  nand2 gate278(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate279(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate280(.a(N69), .O(gate188inter7));
  inv1  gate281(.a(N709), .O(gate188inter8));
  nand2 gate282(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate283(.a(s_11), .b(gate188inter3), .O(gate188inter10));
  nor2  gate284(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate285(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate286(.a(gate188inter12), .b(gate188inter1), .O(N741));
xor2 gate189( .a(N73), .b(N710), .O(N742) );

  xor2  gate455(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate456(.a(gate190inter0), .b(s_36), .O(gate190inter1));
  and2  gate457(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate458(.a(s_36), .O(gate190inter3));
  inv1  gate459(.a(s_37), .O(gate190inter4));
  nand2 gate460(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate461(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate462(.a(N77), .O(gate190inter7));
  inv1  gate463(.a(N711), .O(gate190inter8));
  nand2 gate464(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate465(.a(s_37), .b(gate190inter3), .O(gate190inter10));
  nor2  gate466(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate467(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate468(.a(gate190inter12), .b(gate190inter1), .O(N743));
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );

  xor2  gate259(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate260(.a(gate194inter0), .b(s_8), .O(gate194inter1));
  and2  gate261(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate262(.a(s_8), .O(gate194inter3));
  inv1  gate263(.a(s_9), .O(gate194inter4));
  nand2 gate264(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate265(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate266(.a(N93), .O(gate194inter7));
  inv1  gate267(.a(N715), .O(gate194inter8));
  nand2 gate268(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate269(.a(s_9), .b(gate194inter3), .O(gate194inter10));
  nor2  gate270(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate271(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate272(.a(gate194inter12), .b(gate194inter1), .O(N747));
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );

  xor2  gate581(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate582(.a(gate198inter0), .b(s_54), .O(gate198inter1));
  and2  gate583(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate584(.a(s_54), .O(gate198inter3));
  inv1  gate585(.a(s_55), .O(gate198inter4));
  nand2 gate586(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate587(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate588(.a(N109), .O(gate198inter7));
  inv1  gate589(.a(N719), .O(gate198inter8));
  nand2 gate590(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate591(.a(s_55), .b(gate198inter3), .O(gate198inter10));
  nor2  gate592(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate593(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate594(.a(gate198inter12), .b(gate198inter1), .O(N751));

  xor2  gate665(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate666(.a(gate199inter0), .b(s_66), .O(gate199inter1));
  and2  gate667(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate668(.a(s_66), .O(gate199inter3));
  inv1  gate669(.a(s_67), .O(gate199inter4));
  nand2 gate670(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate671(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate672(.a(N113), .O(gate199inter7));
  inv1  gate673(.a(N720), .O(gate199inter8));
  nand2 gate674(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate675(.a(s_67), .b(gate199inter3), .O(gate199inter10));
  nor2  gate676(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate677(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate678(.a(gate199inter12), .b(gate199inter1), .O(N752));
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate679(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate680(.a(gate201inter0), .b(s_68), .O(gate201inter1));
  and2  gate681(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate682(.a(s_68), .O(gate201inter3));
  inv1  gate683(.a(s_69), .O(gate201inter4));
  nand2 gate684(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate685(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate686(.a(N121), .O(gate201inter7));
  inv1  gate687(.a(N722), .O(gate201inter8));
  nand2 gate688(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate689(.a(s_69), .b(gate201inter3), .O(gate201inter10));
  nor2  gate690(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate691(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate692(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule