module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate357(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate358(.a(gate19inter0), .b(s_28), .O(gate19inter1));
  and2  gate359(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate360(.a(s_28), .O(gate19inter3));
  inv1  gate361(.a(s_29), .O(gate19inter4));
  nand2 gate362(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate363(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate364(.a(N118), .O(gate19inter7));
  inv1  gate365(.a(N4), .O(gate19inter8));
  nand2 gate366(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate367(.a(s_29), .b(gate19inter3), .O(gate19inter10));
  nor2  gate368(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate369(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate370(.a(gate19inter12), .b(gate19inter1), .O(N154));
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate329(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate330(.a(gate29inter0), .b(s_24), .O(gate29inter1));
  and2  gate331(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate332(.a(s_24), .O(gate29inter3));
  inv1  gate333(.a(s_25), .O(gate29inter4));
  nand2 gate334(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate335(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate336(.a(N150), .O(gate29inter7));
  inv1  gate337(.a(N108), .O(gate29inter8));
  nand2 gate338(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate339(.a(s_25), .b(gate29inter3), .O(gate29inter10));
  nor2  gate340(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate341(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate342(.a(gate29inter12), .b(gate29inter1), .O(N180));

  xor2  gate315(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate316(.a(gate30inter0), .b(s_22), .O(gate30inter1));
  and2  gate317(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate318(.a(s_22), .O(gate30inter3));
  inv1  gate319(.a(s_23), .O(gate30inter4));
  nand2 gate320(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate321(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate322(.a(N21), .O(gate30inter7));
  inv1  gate323(.a(N123), .O(gate30inter8));
  nand2 gate324(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate325(.a(s_23), .b(gate30inter3), .O(gate30inter10));
  nor2  gate326(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate327(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate328(.a(gate30inter12), .b(gate30inter1), .O(N183));
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );

  xor2  gate427(.a(N127), .b(N40), .O(gate33inter0));
  nand2 gate428(.a(gate33inter0), .b(s_38), .O(gate33inter1));
  and2  gate429(.a(N127), .b(N40), .O(gate33inter2));
  inv1  gate430(.a(s_38), .O(gate33inter3));
  inv1  gate431(.a(s_39), .O(gate33inter4));
  nand2 gate432(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate433(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate434(.a(N40), .O(gate33inter7));
  inv1  gate435(.a(N127), .O(gate33inter8));
  nand2 gate436(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate437(.a(s_39), .b(gate33inter3), .O(gate33inter10));
  nor2  gate438(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate439(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate440(.a(gate33inter12), .b(gate33inter1), .O(N186));
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate399(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate400(.a(gate37inter0), .b(s_34), .O(gate37inter1));
  and2  gate401(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate402(.a(s_34), .O(gate37inter3));
  inv1  gate403(.a(s_35), .O(gate37inter4));
  nand2 gate404(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate405(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate406(.a(N66), .O(gate37inter7));
  inv1  gate407(.a(N135), .O(gate37inter8));
  nand2 gate408(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate409(.a(s_35), .b(gate37inter3), .O(gate37inter10));
  nor2  gate410(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate411(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate412(.a(gate37inter12), .b(gate37inter1), .O(N190));
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate371(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate372(.a(gate52inter0), .b(s_30), .O(gate52inter1));
  and2  gate373(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate374(.a(s_30), .O(gate52inter3));
  inv1  gate375(.a(s_31), .O(gate52inter4));
  nand2 gate376(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate377(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate378(.a(N203), .O(gate52inter7));
  inv1  gate379(.a(N162), .O(gate52inter8));
  nand2 gate380(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate381(.a(s_31), .b(gate52inter3), .O(gate52inter10));
  nor2  gate382(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate383(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate384(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );

  xor2  gate217(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate218(.a(gate67inter0), .b(s_8), .O(gate67inter1));
  and2  gate219(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate220(.a(s_8), .O(gate67inter3));
  inv1  gate221(.a(s_9), .O(gate67inter4));
  nand2 gate222(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate223(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate224(.a(N213), .O(gate67inter7));
  inv1  gate225(.a(N102), .O(gate67inter8));
  nand2 gate226(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate227(.a(s_9), .b(gate67inter3), .O(gate67inter10));
  nor2  gate228(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate229(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate230(.a(gate67inter12), .b(gate67inter1), .O(N259));
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate189(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate190(.a(gate71inter0), .b(s_4), .O(gate71inter1));
  and2  gate191(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate192(.a(s_4), .O(gate71inter3));
  inv1  gate193(.a(s_5), .O(gate71inter4));
  nand2 gate194(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate195(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate196(.a(N230), .O(gate71inter7));
  inv1  gate197(.a(N185), .O(gate71inter8));
  nand2 gate198(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate199(.a(s_5), .b(gate71inter3), .O(gate71inter10));
  nor2  gate200(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate201(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate202(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate273(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate274(.a(gate73inter0), .b(s_16), .O(gate73inter1));
  and2  gate275(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate276(.a(s_16), .O(gate73inter3));
  inv1  gate277(.a(s_17), .O(gate73inter4));
  nand2 gate278(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate279(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate280(.a(N236), .O(gate73inter7));
  inv1  gate281(.a(N189), .O(gate73inter8));
  nand2 gate282(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate283(.a(s_17), .b(gate73inter3), .O(gate73inter10));
  nor2  gate284(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate285(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate286(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );

  xor2  gate413(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate414(.a(gate84inter0), .b(s_36), .O(gate84inter1));
  and2  gate415(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate416(.a(s_36), .O(gate84inter3));
  inv1  gate417(.a(s_37), .O(gate84inter4));
  nand2 gate418(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate419(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate420(.a(N247), .O(gate84inter7));
  inv1  gate421(.a(N196), .O(gate84inter8));
  nand2 gate422(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate423(.a(s_37), .b(gate84inter3), .O(gate84inter10));
  nor2  gate424(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate425(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate426(.a(gate84inter12), .b(gate84inter1), .O(N294));
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate385(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate386(.a(gate99inter0), .b(s_32), .O(gate99inter1));
  and2  gate387(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate388(.a(s_32), .O(gate99inter3));
  inv1  gate389(.a(s_33), .O(gate99inter4));
  nand2 gate390(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate391(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate392(.a(N309), .O(gate99inter7));
  inv1  gate393(.a(N260), .O(gate99inter8));
  nand2 gate394(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate395(.a(s_33), .b(gate99inter3), .O(gate99inter10));
  nor2  gate396(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate397(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate398(.a(gate99inter12), .b(gate99inter1), .O(N330));
xor2 gate100( .a(N309), .b(N264), .O(N331) );

  xor2  gate259(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate260(.a(gate101inter0), .b(s_14), .O(gate101inter1));
  and2  gate261(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate262(.a(s_14), .O(gate101inter3));
  inv1  gate263(.a(s_15), .O(gate101inter4));
  nand2 gate264(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate265(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate266(.a(N309), .O(gate101inter7));
  inv1  gate267(.a(N267), .O(gate101inter8));
  nand2 gate268(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate269(.a(s_15), .b(gate101inter3), .O(gate101inter10));
  nor2  gate270(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate271(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate272(.a(gate101inter12), .b(gate101inter1), .O(N332));
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate203(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate204(.a(gate111inter0), .b(s_6), .O(gate111inter1));
  and2  gate205(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate206(.a(s_6), .O(gate111inter3));
  inv1  gate207(.a(s_7), .O(gate111inter4));
  nand2 gate208(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate209(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate210(.a(N319), .O(gate111inter7));
  inv1  gate211(.a(N60), .O(gate111inter8));
  nand2 gate212(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate213(.a(s_7), .b(gate111inter3), .O(gate111inter10));
  nor2  gate214(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate215(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate216(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );

  xor2  gate161(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate162(.a(gate114inter0), .b(s_0), .O(gate114inter1));
  and2  gate163(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate164(.a(s_0), .O(gate114inter3));
  inv1  gate165(.a(s_1), .O(gate114inter4));
  nand2 gate166(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate167(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate168(.a(N319), .O(gate114inter7));
  inv1  gate169(.a(N86), .O(gate114inter8));
  nand2 gate170(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate171(.a(s_1), .b(gate114inter3), .O(gate114inter10));
  nor2  gate172(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate173(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate174(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );

  xor2  gate231(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate232(.a(gate117inter0), .b(s_10), .O(gate117inter1));
  and2  gate233(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate234(.a(s_10), .O(gate117inter3));
  inv1  gate235(.a(s_11), .O(gate117inter4));
  nand2 gate236(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate237(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate238(.a(N330), .O(gate117inter7));
  inv1  gate239(.a(N300), .O(gate117inter8));
  nand2 gate240(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate241(.a(s_11), .b(gate117inter3), .O(gate117inter10));
  nor2  gate242(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate243(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate244(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate441(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate442(.a(gate119inter0), .b(s_40), .O(gate119inter1));
  and2  gate443(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate444(.a(s_40), .O(gate119inter3));
  inv1  gate445(.a(s_41), .O(gate119inter4));
  nand2 gate446(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate447(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate448(.a(N332), .O(gate119inter7));
  inv1  gate449(.a(N302), .O(gate119inter8));
  nand2 gate450(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate451(.a(s_41), .b(gate119inter3), .O(gate119inter10));
  nor2  gate452(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate453(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate454(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate175(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate176(.a(gate121inter0), .b(s_2), .O(gate121inter1));
  and2  gate177(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate178(.a(s_2), .O(gate121inter3));
  inv1  gate179(.a(s_3), .O(gate121inter4));
  nand2 gate180(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate181(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate182(.a(N335), .O(gate121inter7));
  inv1  gate183(.a(N304), .O(gate121inter8));
  nand2 gate184(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate185(.a(s_3), .b(gate121inter3), .O(gate121inter10));
  nor2  gate186(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate187(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate188(.a(gate121inter12), .b(gate121inter1), .O(N352));
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate287(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate288(.a(gate131inter0), .b(s_18), .O(gate131inter1));
  and2  gate289(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate290(.a(s_18), .O(gate131inter3));
  inv1  gate291(.a(s_19), .O(gate131inter4));
  nand2 gate292(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate293(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate294(.a(N360), .O(gate131inter7));
  inv1  gate295(.a(N40), .O(gate131inter8));
  nand2 gate296(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate297(.a(s_19), .b(gate131inter3), .O(gate131inter10));
  nor2  gate298(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate299(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate300(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate301(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate302(.a(gate136inter0), .b(s_20), .O(gate136inter1));
  and2  gate303(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate304(.a(s_20), .O(gate136inter3));
  inv1  gate305(.a(s_21), .O(gate136inter4));
  nand2 gate306(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate307(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate308(.a(N360), .O(gate136inter7));
  inv1  gate309(.a(N105), .O(gate136inter8));
  nand2 gate310(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate311(.a(s_21), .b(gate136inter3), .O(gate136inter10));
  nor2  gate312(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate313(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate314(.a(gate136inter12), .b(gate136inter1), .O(N378));

  xor2  gate343(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate344(.a(gate137inter0), .b(s_26), .O(gate137inter1));
  and2  gate345(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate346(.a(s_26), .O(gate137inter3));
  inv1  gate347(.a(s_27), .O(gate137inter4));
  nand2 gate348(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate349(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate350(.a(N360), .O(gate137inter7));
  inv1  gate351(.a(N115), .O(gate137inter8));
  nand2 gate352(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate353(.a(s_27), .b(gate137inter3), .O(gate137inter10));
  nor2  gate354(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate355(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate356(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate245(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate246(.a(gate153inter0), .b(s_12), .O(gate153inter1));
  and2  gate247(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate248(.a(s_12), .O(gate153inter3));
  inv1  gate249(.a(s_13), .O(gate153inter4));
  nand2 gate250(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate251(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate252(.a(N415), .O(gate153inter7));
  inv1  gate253(.a(N416), .O(gate153inter8));
  nand2 gate254(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate255(.a(s_13), .b(gate153inter3), .O(gate153inter10));
  nor2  gate256(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate257(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate258(.a(gate153inter12), .b(gate153inter1), .O(N421));
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule