module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1555(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1556(.a(gate9inter0), .b(s_144), .O(gate9inter1));
  and2  gate1557(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1558(.a(s_144), .O(gate9inter3));
  inv1  gate1559(.a(s_145), .O(gate9inter4));
  nand2 gate1560(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1561(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1562(.a(G1), .O(gate9inter7));
  inv1  gate1563(.a(G2), .O(gate9inter8));
  nand2 gate1564(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1565(.a(s_145), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1566(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1567(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1568(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate729(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate730(.a(gate12inter0), .b(s_26), .O(gate12inter1));
  and2  gate731(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate732(.a(s_26), .O(gate12inter3));
  inv1  gate733(.a(s_27), .O(gate12inter4));
  nand2 gate734(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate735(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate736(.a(G7), .O(gate12inter7));
  inv1  gate737(.a(G8), .O(gate12inter8));
  nand2 gate738(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate739(.a(s_27), .b(gate12inter3), .O(gate12inter10));
  nor2  gate740(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate741(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate742(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1247(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1248(.a(gate28inter0), .b(s_100), .O(gate28inter1));
  and2  gate1249(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1250(.a(s_100), .O(gate28inter3));
  inv1  gate1251(.a(s_101), .O(gate28inter4));
  nand2 gate1252(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1253(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1254(.a(G10), .O(gate28inter7));
  inv1  gate1255(.a(G14), .O(gate28inter8));
  nand2 gate1256(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1257(.a(s_101), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1258(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1259(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1260(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1345(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1346(.a(gate29inter0), .b(s_114), .O(gate29inter1));
  and2  gate1347(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1348(.a(s_114), .O(gate29inter3));
  inv1  gate1349(.a(s_115), .O(gate29inter4));
  nand2 gate1350(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1351(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1352(.a(G3), .O(gate29inter7));
  inv1  gate1353(.a(G7), .O(gate29inter8));
  nand2 gate1354(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1355(.a(s_115), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1356(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1357(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1358(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1275(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1276(.a(gate30inter0), .b(s_104), .O(gate30inter1));
  and2  gate1277(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1278(.a(s_104), .O(gate30inter3));
  inv1  gate1279(.a(s_105), .O(gate30inter4));
  nand2 gate1280(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1281(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1282(.a(G11), .O(gate30inter7));
  inv1  gate1283(.a(G15), .O(gate30inter8));
  nand2 gate1284(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1285(.a(s_105), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1286(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1287(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1288(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate715(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate716(.a(gate33inter0), .b(s_24), .O(gate33inter1));
  and2  gate717(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate718(.a(s_24), .O(gate33inter3));
  inv1  gate719(.a(s_25), .O(gate33inter4));
  nand2 gate720(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate721(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate722(.a(G17), .O(gate33inter7));
  inv1  gate723(.a(G21), .O(gate33inter8));
  nand2 gate724(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate725(.a(s_25), .b(gate33inter3), .O(gate33inter10));
  nor2  gate726(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate727(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate728(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1877(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1878(.a(gate37inter0), .b(s_190), .O(gate37inter1));
  and2  gate1879(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1880(.a(s_190), .O(gate37inter3));
  inv1  gate1881(.a(s_191), .O(gate37inter4));
  nand2 gate1882(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1883(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1884(.a(G19), .O(gate37inter7));
  inv1  gate1885(.a(G23), .O(gate37inter8));
  nand2 gate1886(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1887(.a(s_191), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1888(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1889(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1890(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1653(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1654(.a(gate41inter0), .b(s_158), .O(gate41inter1));
  and2  gate1655(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1656(.a(s_158), .O(gate41inter3));
  inv1  gate1657(.a(s_159), .O(gate41inter4));
  nand2 gate1658(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1659(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1660(.a(G1), .O(gate41inter7));
  inv1  gate1661(.a(G266), .O(gate41inter8));
  nand2 gate1662(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1663(.a(s_159), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1664(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1665(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1666(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate981(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate982(.a(gate49inter0), .b(s_62), .O(gate49inter1));
  and2  gate983(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate984(.a(s_62), .O(gate49inter3));
  inv1  gate985(.a(s_63), .O(gate49inter4));
  nand2 gate986(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate987(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate988(.a(G9), .O(gate49inter7));
  inv1  gate989(.a(G278), .O(gate49inter8));
  nand2 gate990(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate991(.a(s_63), .b(gate49inter3), .O(gate49inter10));
  nor2  gate992(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate993(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate994(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1233(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1234(.a(gate51inter0), .b(s_98), .O(gate51inter1));
  and2  gate1235(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1236(.a(s_98), .O(gate51inter3));
  inv1  gate1237(.a(s_99), .O(gate51inter4));
  nand2 gate1238(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1239(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1240(.a(G11), .O(gate51inter7));
  inv1  gate1241(.a(G281), .O(gate51inter8));
  nand2 gate1242(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1243(.a(s_99), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1244(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1245(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1246(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate799(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate800(.a(gate52inter0), .b(s_36), .O(gate52inter1));
  and2  gate801(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate802(.a(s_36), .O(gate52inter3));
  inv1  gate803(.a(s_37), .O(gate52inter4));
  nand2 gate804(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate805(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate806(.a(G12), .O(gate52inter7));
  inv1  gate807(.a(G281), .O(gate52inter8));
  nand2 gate808(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate809(.a(s_37), .b(gate52inter3), .O(gate52inter10));
  nor2  gate810(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate811(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate812(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1415(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1416(.a(gate55inter0), .b(s_124), .O(gate55inter1));
  and2  gate1417(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1418(.a(s_124), .O(gate55inter3));
  inv1  gate1419(.a(s_125), .O(gate55inter4));
  nand2 gate1420(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1421(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1422(.a(G15), .O(gate55inter7));
  inv1  gate1423(.a(G287), .O(gate55inter8));
  nand2 gate1424(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1425(.a(s_125), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1426(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1427(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1428(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1667(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1668(.a(gate65inter0), .b(s_160), .O(gate65inter1));
  and2  gate1669(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1670(.a(s_160), .O(gate65inter3));
  inv1  gate1671(.a(s_161), .O(gate65inter4));
  nand2 gate1672(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1673(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1674(.a(G25), .O(gate65inter7));
  inv1  gate1675(.a(G302), .O(gate65inter8));
  nand2 gate1676(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1677(.a(s_161), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1678(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1679(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1680(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1359(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1360(.a(gate71inter0), .b(s_116), .O(gate71inter1));
  and2  gate1361(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1362(.a(s_116), .O(gate71inter3));
  inv1  gate1363(.a(s_117), .O(gate71inter4));
  nand2 gate1364(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1365(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1366(.a(G31), .O(gate71inter7));
  inv1  gate1367(.a(G311), .O(gate71inter8));
  nand2 gate1368(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1369(.a(s_117), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1370(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1371(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1372(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1429(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1430(.a(gate80inter0), .b(s_126), .O(gate80inter1));
  and2  gate1431(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1432(.a(s_126), .O(gate80inter3));
  inv1  gate1433(.a(s_127), .O(gate80inter4));
  nand2 gate1434(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1435(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1436(.a(G14), .O(gate80inter7));
  inv1  gate1437(.a(G323), .O(gate80inter8));
  nand2 gate1438(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1439(.a(s_127), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1440(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1441(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1442(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate589(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate590(.a(gate82inter0), .b(s_6), .O(gate82inter1));
  and2  gate591(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate592(.a(s_6), .O(gate82inter3));
  inv1  gate593(.a(s_7), .O(gate82inter4));
  nand2 gate594(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate595(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate596(.a(G7), .O(gate82inter7));
  inv1  gate597(.a(G326), .O(gate82inter8));
  nand2 gate598(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate599(.a(s_7), .b(gate82inter3), .O(gate82inter10));
  nor2  gate600(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate601(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate602(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1583(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1584(.a(gate83inter0), .b(s_148), .O(gate83inter1));
  and2  gate1585(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1586(.a(s_148), .O(gate83inter3));
  inv1  gate1587(.a(s_149), .O(gate83inter4));
  nand2 gate1588(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1589(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1590(.a(G11), .O(gate83inter7));
  inv1  gate1591(.a(G329), .O(gate83inter8));
  nand2 gate1592(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1593(.a(s_149), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1594(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1595(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1596(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate855(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate856(.a(gate102inter0), .b(s_44), .O(gate102inter1));
  and2  gate857(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate858(.a(s_44), .O(gate102inter3));
  inv1  gate859(.a(s_45), .O(gate102inter4));
  nand2 gate860(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate861(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate862(.a(G24), .O(gate102inter7));
  inv1  gate863(.a(G356), .O(gate102inter8));
  nand2 gate864(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate865(.a(s_45), .b(gate102inter3), .O(gate102inter10));
  nor2  gate866(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate867(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate868(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate869(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate870(.a(gate104inter0), .b(s_46), .O(gate104inter1));
  and2  gate871(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate872(.a(s_46), .O(gate104inter3));
  inv1  gate873(.a(s_47), .O(gate104inter4));
  nand2 gate874(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate875(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate876(.a(G32), .O(gate104inter7));
  inv1  gate877(.a(G359), .O(gate104inter8));
  nand2 gate878(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate879(.a(s_47), .b(gate104inter3), .O(gate104inter10));
  nor2  gate880(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate881(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate882(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1849(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1850(.a(gate106inter0), .b(s_186), .O(gate106inter1));
  and2  gate1851(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1852(.a(s_186), .O(gate106inter3));
  inv1  gate1853(.a(s_187), .O(gate106inter4));
  nand2 gate1854(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1855(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1856(.a(G364), .O(gate106inter7));
  inv1  gate1857(.a(G365), .O(gate106inter8));
  nand2 gate1858(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1859(.a(s_187), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1860(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1861(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1862(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1373(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1374(.a(gate107inter0), .b(s_118), .O(gate107inter1));
  and2  gate1375(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1376(.a(s_118), .O(gate107inter3));
  inv1  gate1377(.a(s_119), .O(gate107inter4));
  nand2 gate1378(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1379(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1380(.a(G366), .O(gate107inter7));
  inv1  gate1381(.a(G367), .O(gate107inter8));
  nand2 gate1382(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1383(.a(s_119), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1384(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1385(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1386(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1541(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1542(.a(gate116inter0), .b(s_142), .O(gate116inter1));
  and2  gate1543(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1544(.a(s_142), .O(gate116inter3));
  inv1  gate1545(.a(s_143), .O(gate116inter4));
  nand2 gate1546(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1547(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1548(.a(G384), .O(gate116inter7));
  inv1  gate1549(.a(G385), .O(gate116inter8));
  nand2 gate1550(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1551(.a(s_143), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1552(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1553(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1554(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1527(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1528(.a(gate125inter0), .b(s_140), .O(gate125inter1));
  and2  gate1529(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1530(.a(s_140), .O(gate125inter3));
  inv1  gate1531(.a(s_141), .O(gate125inter4));
  nand2 gate1532(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1533(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1534(.a(G402), .O(gate125inter7));
  inv1  gate1535(.a(G403), .O(gate125inter8));
  nand2 gate1536(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1537(.a(s_141), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1538(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1539(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1540(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate911(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate912(.a(gate131inter0), .b(s_52), .O(gate131inter1));
  and2  gate913(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate914(.a(s_52), .O(gate131inter3));
  inv1  gate915(.a(s_53), .O(gate131inter4));
  nand2 gate916(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate917(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate918(.a(G414), .O(gate131inter7));
  inv1  gate919(.a(G415), .O(gate131inter8));
  nand2 gate920(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate921(.a(s_53), .b(gate131inter3), .O(gate131inter10));
  nor2  gate922(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate923(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate924(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1023(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1024(.a(gate137inter0), .b(s_68), .O(gate137inter1));
  and2  gate1025(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1026(.a(s_68), .O(gate137inter3));
  inv1  gate1027(.a(s_69), .O(gate137inter4));
  nand2 gate1028(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1029(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1030(.a(G426), .O(gate137inter7));
  inv1  gate1031(.a(G429), .O(gate137inter8));
  nand2 gate1032(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1033(.a(s_69), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1034(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1035(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1036(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1079(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1080(.a(gate138inter0), .b(s_76), .O(gate138inter1));
  and2  gate1081(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1082(.a(s_76), .O(gate138inter3));
  inv1  gate1083(.a(s_77), .O(gate138inter4));
  nand2 gate1084(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1085(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1086(.a(G432), .O(gate138inter7));
  inv1  gate1087(.a(G435), .O(gate138inter8));
  nand2 gate1088(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1089(.a(s_77), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1090(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1091(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1092(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1639(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1640(.a(gate143inter0), .b(s_156), .O(gate143inter1));
  and2  gate1641(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1642(.a(s_156), .O(gate143inter3));
  inv1  gate1643(.a(s_157), .O(gate143inter4));
  nand2 gate1644(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1645(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1646(.a(G462), .O(gate143inter7));
  inv1  gate1647(.a(G465), .O(gate143inter8));
  nand2 gate1648(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1649(.a(s_157), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1650(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1651(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1652(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1443(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1444(.a(gate145inter0), .b(s_128), .O(gate145inter1));
  and2  gate1445(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1446(.a(s_128), .O(gate145inter3));
  inv1  gate1447(.a(s_129), .O(gate145inter4));
  nand2 gate1448(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1449(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1450(.a(G474), .O(gate145inter7));
  inv1  gate1451(.a(G477), .O(gate145inter8));
  nand2 gate1452(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1453(.a(s_129), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1454(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1455(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1456(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1765(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1766(.a(gate148inter0), .b(s_174), .O(gate148inter1));
  and2  gate1767(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1768(.a(s_174), .O(gate148inter3));
  inv1  gate1769(.a(s_175), .O(gate148inter4));
  nand2 gate1770(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1771(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1772(.a(G492), .O(gate148inter7));
  inv1  gate1773(.a(G495), .O(gate148inter8));
  nand2 gate1774(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1775(.a(s_175), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1776(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1777(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1778(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1485(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1486(.a(gate161inter0), .b(s_134), .O(gate161inter1));
  and2  gate1487(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1488(.a(s_134), .O(gate161inter3));
  inv1  gate1489(.a(s_135), .O(gate161inter4));
  nand2 gate1490(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1491(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1492(.a(G450), .O(gate161inter7));
  inv1  gate1493(.a(G534), .O(gate161inter8));
  nand2 gate1494(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1495(.a(s_135), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1496(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1497(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1498(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1401(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1402(.a(gate175inter0), .b(s_122), .O(gate175inter1));
  and2  gate1403(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1404(.a(s_122), .O(gate175inter3));
  inv1  gate1405(.a(s_123), .O(gate175inter4));
  nand2 gate1406(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1407(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1408(.a(G492), .O(gate175inter7));
  inv1  gate1409(.a(G555), .O(gate175inter8));
  nand2 gate1410(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1411(.a(s_123), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1412(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1413(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1414(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1107(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1108(.a(gate178inter0), .b(s_80), .O(gate178inter1));
  and2  gate1109(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1110(.a(s_80), .O(gate178inter3));
  inv1  gate1111(.a(s_81), .O(gate178inter4));
  nand2 gate1112(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1113(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1114(.a(G501), .O(gate178inter7));
  inv1  gate1115(.a(G558), .O(gate178inter8));
  nand2 gate1116(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1117(.a(s_81), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1118(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1119(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1120(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1191(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1192(.a(gate180inter0), .b(s_92), .O(gate180inter1));
  and2  gate1193(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1194(.a(s_92), .O(gate180inter3));
  inv1  gate1195(.a(s_93), .O(gate180inter4));
  nand2 gate1196(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1197(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1198(.a(G507), .O(gate180inter7));
  inv1  gate1199(.a(G561), .O(gate180inter8));
  nand2 gate1200(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1201(.a(s_93), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1202(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1203(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1204(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate673(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate674(.a(gate181inter0), .b(s_18), .O(gate181inter1));
  and2  gate675(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate676(.a(s_18), .O(gate181inter3));
  inv1  gate677(.a(s_19), .O(gate181inter4));
  nand2 gate678(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate679(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate680(.a(G510), .O(gate181inter7));
  inv1  gate681(.a(G564), .O(gate181inter8));
  nand2 gate682(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate683(.a(s_19), .b(gate181inter3), .O(gate181inter10));
  nor2  gate684(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate685(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate686(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1219(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1220(.a(gate182inter0), .b(s_96), .O(gate182inter1));
  and2  gate1221(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1222(.a(s_96), .O(gate182inter3));
  inv1  gate1223(.a(s_97), .O(gate182inter4));
  nand2 gate1224(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1225(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1226(.a(G513), .O(gate182inter7));
  inv1  gate1227(.a(G564), .O(gate182inter8));
  nand2 gate1228(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1229(.a(s_97), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1230(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1231(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1232(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1737(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1738(.a(gate184inter0), .b(s_170), .O(gate184inter1));
  and2  gate1739(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1740(.a(s_170), .O(gate184inter3));
  inv1  gate1741(.a(s_171), .O(gate184inter4));
  nand2 gate1742(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1743(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1744(.a(G519), .O(gate184inter7));
  inv1  gate1745(.a(G567), .O(gate184inter8));
  nand2 gate1746(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1747(.a(s_171), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1748(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1749(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1750(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1499(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1500(.a(gate188inter0), .b(s_136), .O(gate188inter1));
  and2  gate1501(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1502(.a(s_136), .O(gate188inter3));
  inv1  gate1503(.a(s_137), .O(gate188inter4));
  nand2 gate1504(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1505(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1506(.a(G576), .O(gate188inter7));
  inv1  gate1507(.a(G577), .O(gate188inter8));
  nand2 gate1508(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1509(.a(s_137), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1510(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1511(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1512(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate659(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate660(.a(gate194inter0), .b(s_16), .O(gate194inter1));
  and2  gate661(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate662(.a(s_16), .O(gate194inter3));
  inv1  gate663(.a(s_17), .O(gate194inter4));
  nand2 gate664(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate665(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate666(.a(G588), .O(gate194inter7));
  inv1  gate667(.a(G589), .O(gate194inter8));
  nand2 gate668(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate669(.a(s_17), .b(gate194inter3), .O(gate194inter10));
  nor2  gate670(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate671(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate672(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate617(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate618(.a(gate196inter0), .b(s_10), .O(gate196inter1));
  and2  gate619(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate620(.a(s_10), .O(gate196inter3));
  inv1  gate621(.a(s_11), .O(gate196inter4));
  nand2 gate622(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate623(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate624(.a(G592), .O(gate196inter7));
  inv1  gate625(.a(G593), .O(gate196inter8));
  nand2 gate626(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate627(.a(s_11), .b(gate196inter3), .O(gate196inter10));
  nor2  gate628(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate629(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate630(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1681(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1682(.a(gate197inter0), .b(s_162), .O(gate197inter1));
  and2  gate1683(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1684(.a(s_162), .O(gate197inter3));
  inv1  gate1685(.a(s_163), .O(gate197inter4));
  nand2 gate1686(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1687(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1688(.a(G594), .O(gate197inter7));
  inv1  gate1689(.a(G595), .O(gate197inter8));
  nand2 gate1690(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1691(.a(s_163), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1692(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1693(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1694(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate645(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate646(.a(gate198inter0), .b(s_14), .O(gate198inter1));
  and2  gate647(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate648(.a(s_14), .O(gate198inter3));
  inv1  gate649(.a(s_15), .O(gate198inter4));
  nand2 gate650(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate651(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate652(.a(G596), .O(gate198inter7));
  inv1  gate653(.a(G597), .O(gate198inter8));
  nand2 gate654(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate655(.a(s_15), .b(gate198inter3), .O(gate198inter10));
  nor2  gate656(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate657(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate658(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1037(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1038(.a(gate205inter0), .b(s_70), .O(gate205inter1));
  and2  gate1039(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1040(.a(s_70), .O(gate205inter3));
  inv1  gate1041(.a(s_71), .O(gate205inter4));
  nand2 gate1042(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1043(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1044(.a(G622), .O(gate205inter7));
  inv1  gate1045(.a(G627), .O(gate205inter8));
  nand2 gate1046(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1047(.a(s_71), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1048(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1049(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1050(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1779(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1780(.a(gate209inter0), .b(s_176), .O(gate209inter1));
  and2  gate1781(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1782(.a(s_176), .O(gate209inter3));
  inv1  gate1783(.a(s_177), .O(gate209inter4));
  nand2 gate1784(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1785(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1786(.a(G602), .O(gate209inter7));
  inv1  gate1787(.a(G666), .O(gate209inter8));
  nand2 gate1788(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1789(.a(s_177), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1790(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1791(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1792(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1807(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1808(.a(gate212inter0), .b(s_180), .O(gate212inter1));
  and2  gate1809(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1810(.a(s_180), .O(gate212inter3));
  inv1  gate1811(.a(s_181), .O(gate212inter4));
  nand2 gate1812(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1813(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1814(.a(G617), .O(gate212inter7));
  inv1  gate1815(.a(G669), .O(gate212inter8));
  nand2 gate1816(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1817(.a(s_181), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1818(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1819(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1820(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1205(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1206(.a(gate221inter0), .b(s_94), .O(gate221inter1));
  and2  gate1207(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1208(.a(s_94), .O(gate221inter3));
  inv1  gate1209(.a(s_95), .O(gate221inter4));
  nand2 gate1210(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1211(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1212(.a(G622), .O(gate221inter7));
  inv1  gate1213(.a(G684), .O(gate221inter8));
  nand2 gate1214(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1215(.a(s_95), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1216(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1217(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1218(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate743(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate744(.a(gate223inter0), .b(s_28), .O(gate223inter1));
  and2  gate745(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate746(.a(s_28), .O(gate223inter3));
  inv1  gate747(.a(s_29), .O(gate223inter4));
  nand2 gate748(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate749(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate750(.a(G627), .O(gate223inter7));
  inv1  gate751(.a(G687), .O(gate223inter8));
  nand2 gate752(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate753(.a(s_29), .b(gate223inter3), .O(gate223inter10));
  nor2  gate754(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate755(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate756(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1051(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1052(.a(gate226inter0), .b(s_72), .O(gate226inter1));
  and2  gate1053(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1054(.a(s_72), .O(gate226inter3));
  inv1  gate1055(.a(s_73), .O(gate226inter4));
  nand2 gate1056(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1057(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1058(.a(G692), .O(gate226inter7));
  inv1  gate1059(.a(G693), .O(gate226inter8));
  nand2 gate1060(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1061(.a(s_73), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1062(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1063(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1064(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate939(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate940(.a(gate228inter0), .b(s_56), .O(gate228inter1));
  and2  gate941(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate942(.a(s_56), .O(gate228inter3));
  inv1  gate943(.a(s_57), .O(gate228inter4));
  nand2 gate944(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate945(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate946(.a(G696), .O(gate228inter7));
  inv1  gate947(.a(G697), .O(gate228inter8));
  nand2 gate948(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate949(.a(s_57), .b(gate228inter3), .O(gate228inter10));
  nor2  gate950(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate951(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate952(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1303(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1304(.a(gate233inter0), .b(s_108), .O(gate233inter1));
  and2  gate1305(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1306(.a(s_108), .O(gate233inter3));
  inv1  gate1307(.a(s_109), .O(gate233inter4));
  nand2 gate1308(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1309(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1310(.a(G242), .O(gate233inter7));
  inv1  gate1311(.a(G718), .O(gate233inter8));
  nand2 gate1312(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1313(.a(s_109), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1314(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1315(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1316(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate813(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate814(.a(gate235inter0), .b(s_38), .O(gate235inter1));
  and2  gate815(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate816(.a(s_38), .O(gate235inter3));
  inv1  gate817(.a(s_39), .O(gate235inter4));
  nand2 gate818(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate819(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate820(.a(G248), .O(gate235inter7));
  inv1  gate821(.a(G724), .O(gate235inter8));
  nand2 gate822(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate823(.a(s_39), .b(gate235inter3), .O(gate235inter10));
  nor2  gate824(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate825(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate826(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate1835(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1836(.a(gate236inter0), .b(s_184), .O(gate236inter1));
  and2  gate1837(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1838(.a(s_184), .O(gate236inter3));
  inv1  gate1839(.a(s_185), .O(gate236inter4));
  nand2 gate1840(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1841(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1842(.a(G251), .O(gate236inter7));
  inv1  gate1843(.a(G727), .O(gate236inter8));
  nand2 gate1844(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1845(.a(s_185), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1846(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1847(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1848(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1009(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1010(.a(gate245inter0), .b(s_66), .O(gate245inter1));
  and2  gate1011(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1012(.a(s_66), .O(gate245inter3));
  inv1  gate1013(.a(s_67), .O(gate245inter4));
  nand2 gate1014(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1015(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1016(.a(G248), .O(gate245inter7));
  inv1  gate1017(.a(G736), .O(gate245inter8));
  nand2 gate1018(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1019(.a(s_67), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1020(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1021(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1022(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate771(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate772(.a(gate248inter0), .b(s_32), .O(gate248inter1));
  and2  gate773(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate774(.a(s_32), .O(gate248inter3));
  inv1  gate775(.a(s_33), .O(gate248inter4));
  nand2 gate776(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate777(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate778(.a(G727), .O(gate248inter7));
  inv1  gate779(.a(G739), .O(gate248inter8));
  nand2 gate780(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate781(.a(s_33), .b(gate248inter3), .O(gate248inter10));
  nor2  gate782(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate783(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate784(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1513(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1514(.a(gate251inter0), .b(s_138), .O(gate251inter1));
  and2  gate1515(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1516(.a(s_138), .O(gate251inter3));
  inv1  gate1517(.a(s_139), .O(gate251inter4));
  nand2 gate1518(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1519(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1520(.a(G257), .O(gate251inter7));
  inv1  gate1521(.a(G745), .O(gate251inter8));
  nand2 gate1522(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1523(.a(s_139), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1524(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1525(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1526(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1709(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1710(.a(gate253inter0), .b(s_166), .O(gate253inter1));
  and2  gate1711(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1712(.a(s_166), .O(gate253inter3));
  inv1  gate1713(.a(s_167), .O(gate253inter4));
  nand2 gate1714(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1715(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1716(.a(G260), .O(gate253inter7));
  inv1  gate1717(.a(G748), .O(gate253inter8));
  nand2 gate1718(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1719(.a(s_167), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1720(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1721(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1722(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1387(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1388(.a(gate256inter0), .b(s_120), .O(gate256inter1));
  and2  gate1389(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1390(.a(s_120), .O(gate256inter3));
  inv1  gate1391(.a(s_121), .O(gate256inter4));
  nand2 gate1392(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1393(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1394(.a(G715), .O(gate256inter7));
  inv1  gate1395(.a(G751), .O(gate256inter8));
  nand2 gate1396(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1397(.a(s_121), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1398(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1399(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1400(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate827(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate828(.a(gate262inter0), .b(s_40), .O(gate262inter1));
  and2  gate829(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate830(.a(s_40), .O(gate262inter3));
  inv1  gate831(.a(s_41), .O(gate262inter4));
  nand2 gate832(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate833(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate834(.a(G764), .O(gate262inter7));
  inv1  gate835(.a(G765), .O(gate262inter8));
  nand2 gate836(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate837(.a(s_41), .b(gate262inter3), .O(gate262inter10));
  nor2  gate838(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate839(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate840(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1625(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1626(.a(gate263inter0), .b(s_154), .O(gate263inter1));
  and2  gate1627(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1628(.a(s_154), .O(gate263inter3));
  inv1  gate1629(.a(s_155), .O(gate263inter4));
  nand2 gate1630(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1631(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1632(.a(G766), .O(gate263inter7));
  inv1  gate1633(.a(G767), .O(gate263inter8));
  nand2 gate1634(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1635(.a(s_155), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1636(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1637(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1638(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1331(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1332(.a(gate266inter0), .b(s_112), .O(gate266inter1));
  and2  gate1333(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1334(.a(s_112), .O(gate266inter3));
  inv1  gate1335(.a(s_113), .O(gate266inter4));
  nand2 gate1336(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1337(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1338(.a(G645), .O(gate266inter7));
  inv1  gate1339(.a(G773), .O(gate266inter8));
  nand2 gate1340(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1341(.a(s_113), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1342(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1343(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1344(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate757(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate758(.a(gate269inter0), .b(s_30), .O(gate269inter1));
  and2  gate759(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate760(.a(s_30), .O(gate269inter3));
  inv1  gate761(.a(s_31), .O(gate269inter4));
  nand2 gate762(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate763(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate764(.a(G654), .O(gate269inter7));
  inv1  gate765(.a(G782), .O(gate269inter8));
  nand2 gate766(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate767(.a(s_31), .b(gate269inter3), .O(gate269inter10));
  nor2  gate768(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate769(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate770(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1163(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1164(.a(gate274inter0), .b(s_88), .O(gate274inter1));
  and2  gate1165(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1166(.a(s_88), .O(gate274inter3));
  inv1  gate1167(.a(s_89), .O(gate274inter4));
  nand2 gate1168(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1169(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1170(.a(G770), .O(gate274inter7));
  inv1  gate1171(.a(G794), .O(gate274inter8));
  nand2 gate1172(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1173(.a(s_89), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1174(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1175(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1176(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate575(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate576(.a(gate286inter0), .b(s_4), .O(gate286inter1));
  and2  gate577(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate578(.a(s_4), .O(gate286inter3));
  inv1  gate579(.a(s_5), .O(gate286inter4));
  nand2 gate580(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate581(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate582(.a(G788), .O(gate286inter7));
  inv1  gate583(.a(G812), .O(gate286inter8));
  nand2 gate584(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate585(.a(s_5), .b(gate286inter3), .O(gate286inter10));
  nor2  gate586(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate587(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate588(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1695(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1696(.a(gate292inter0), .b(s_164), .O(gate292inter1));
  and2  gate1697(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1698(.a(s_164), .O(gate292inter3));
  inv1  gate1699(.a(s_165), .O(gate292inter4));
  nand2 gate1700(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1701(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1702(.a(G824), .O(gate292inter7));
  inv1  gate1703(.a(G825), .O(gate292inter8));
  nand2 gate1704(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1705(.a(s_165), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1706(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1707(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1708(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate967(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate968(.a(gate293inter0), .b(s_60), .O(gate293inter1));
  and2  gate969(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate970(.a(s_60), .O(gate293inter3));
  inv1  gate971(.a(s_61), .O(gate293inter4));
  nand2 gate972(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate973(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate974(.a(G828), .O(gate293inter7));
  inv1  gate975(.a(G829), .O(gate293inter8));
  nand2 gate976(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate977(.a(s_61), .b(gate293inter3), .O(gate293inter10));
  nor2  gate978(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate979(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate980(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate603(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate604(.a(gate294inter0), .b(s_8), .O(gate294inter1));
  and2  gate605(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate606(.a(s_8), .O(gate294inter3));
  inv1  gate607(.a(s_9), .O(gate294inter4));
  nand2 gate608(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate609(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate610(.a(G832), .O(gate294inter7));
  inv1  gate611(.a(G833), .O(gate294inter8));
  nand2 gate612(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate613(.a(s_9), .b(gate294inter3), .O(gate294inter10));
  nor2  gate614(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate615(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate616(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1471(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1472(.a(gate387inter0), .b(s_132), .O(gate387inter1));
  and2  gate1473(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1474(.a(s_132), .O(gate387inter3));
  inv1  gate1475(.a(s_133), .O(gate387inter4));
  nand2 gate1476(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1477(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1478(.a(G1), .O(gate387inter7));
  inv1  gate1479(.a(G1036), .O(gate387inter8));
  nand2 gate1480(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1481(.a(s_133), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1482(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1483(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1484(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate897(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate898(.a(gate392inter0), .b(s_50), .O(gate392inter1));
  and2  gate899(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate900(.a(s_50), .O(gate392inter3));
  inv1  gate901(.a(s_51), .O(gate392inter4));
  nand2 gate902(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate903(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate904(.a(G6), .O(gate392inter7));
  inv1  gate905(.a(G1051), .O(gate392inter8));
  nand2 gate906(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate907(.a(s_51), .b(gate392inter3), .O(gate392inter10));
  nor2  gate908(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate909(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate910(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1821(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1822(.a(gate394inter0), .b(s_182), .O(gate394inter1));
  and2  gate1823(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1824(.a(s_182), .O(gate394inter3));
  inv1  gate1825(.a(s_183), .O(gate394inter4));
  nand2 gate1826(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1827(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1828(.a(G8), .O(gate394inter7));
  inv1  gate1829(.a(G1057), .O(gate394inter8));
  nand2 gate1830(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1831(.a(s_183), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1832(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1833(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1834(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate925(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate926(.a(gate400inter0), .b(s_54), .O(gate400inter1));
  and2  gate927(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate928(.a(s_54), .O(gate400inter3));
  inv1  gate929(.a(s_55), .O(gate400inter4));
  nand2 gate930(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate931(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate932(.a(G14), .O(gate400inter7));
  inv1  gate933(.a(G1075), .O(gate400inter8));
  nand2 gate934(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate935(.a(s_55), .b(gate400inter3), .O(gate400inter10));
  nor2  gate936(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate937(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate938(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate631(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate632(.a(gate407inter0), .b(s_12), .O(gate407inter1));
  and2  gate633(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate634(.a(s_12), .O(gate407inter3));
  inv1  gate635(.a(s_13), .O(gate407inter4));
  nand2 gate636(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate637(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate638(.a(G21), .O(gate407inter7));
  inv1  gate639(.a(G1096), .O(gate407inter8));
  nand2 gate640(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate641(.a(s_13), .b(gate407inter3), .O(gate407inter10));
  nor2  gate642(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate643(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate644(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1135(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1136(.a(gate414inter0), .b(s_84), .O(gate414inter1));
  and2  gate1137(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1138(.a(s_84), .O(gate414inter3));
  inv1  gate1139(.a(s_85), .O(gate414inter4));
  nand2 gate1140(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1141(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1142(.a(G28), .O(gate414inter7));
  inv1  gate1143(.a(G1117), .O(gate414inter8));
  nand2 gate1144(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1145(.a(s_85), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1146(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1147(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1148(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1569(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1570(.a(gate417inter0), .b(s_146), .O(gate417inter1));
  and2  gate1571(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1572(.a(s_146), .O(gate417inter3));
  inv1  gate1573(.a(s_147), .O(gate417inter4));
  nand2 gate1574(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1575(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1576(.a(G31), .O(gate417inter7));
  inv1  gate1577(.a(G1126), .O(gate417inter8));
  nand2 gate1578(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1579(.a(s_147), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1580(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1581(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1582(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1723(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1724(.a(gate418inter0), .b(s_168), .O(gate418inter1));
  and2  gate1725(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1726(.a(s_168), .O(gate418inter3));
  inv1  gate1727(.a(s_169), .O(gate418inter4));
  nand2 gate1728(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1729(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1730(.a(G32), .O(gate418inter7));
  inv1  gate1731(.a(G1129), .O(gate418inter8));
  nand2 gate1732(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1733(.a(s_169), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1734(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1735(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1736(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1177(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1178(.a(gate419inter0), .b(s_90), .O(gate419inter1));
  and2  gate1179(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1180(.a(s_90), .O(gate419inter3));
  inv1  gate1181(.a(s_91), .O(gate419inter4));
  nand2 gate1182(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1183(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1184(.a(G1), .O(gate419inter7));
  inv1  gate1185(.a(G1132), .O(gate419inter8));
  nand2 gate1186(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1187(.a(s_91), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1188(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1189(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1190(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate841(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate842(.a(gate421inter0), .b(s_42), .O(gate421inter1));
  and2  gate843(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate844(.a(s_42), .O(gate421inter3));
  inv1  gate845(.a(s_43), .O(gate421inter4));
  nand2 gate846(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate847(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate848(.a(G2), .O(gate421inter7));
  inv1  gate849(.a(G1135), .O(gate421inter8));
  nand2 gate850(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate851(.a(s_43), .b(gate421inter3), .O(gate421inter10));
  nor2  gate852(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate853(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate854(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1597(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1598(.a(gate425inter0), .b(s_150), .O(gate425inter1));
  and2  gate1599(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1600(.a(s_150), .O(gate425inter3));
  inv1  gate1601(.a(s_151), .O(gate425inter4));
  nand2 gate1602(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1603(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1604(.a(G4), .O(gate425inter7));
  inv1  gate1605(.a(G1141), .O(gate425inter8));
  nand2 gate1606(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1607(.a(s_151), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1608(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1609(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1610(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1793(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1794(.a(gate428inter0), .b(s_178), .O(gate428inter1));
  and2  gate1795(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1796(.a(s_178), .O(gate428inter3));
  inv1  gate1797(.a(s_179), .O(gate428inter4));
  nand2 gate1798(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1799(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1800(.a(G1048), .O(gate428inter7));
  inv1  gate1801(.a(G1144), .O(gate428inter8));
  nand2 gate1802(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1803(.a(s_179), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1804(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1805(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1806(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1611(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1612(.a(gate429inter0), .b(s_152), .O(gate429inter1));
  and2  gate1613(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1614(.a(s_152), .O(gate429inter3));
  inv1  gate1615(.a(s_153), .O(gate429inter4));
  nand2 gate1616(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1617(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1618(.a(G6), .O(gate429inter7));
  inv1  gate1619(.a(G1147), .O(gate429inter8));
  nand2 gate1620(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1621(.a(s_153), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1622(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1623(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1624(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1149(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1150(.a(gate434inter0), .b(s_86), .O(gate434inter1));
  and2  gate1151(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1152(.a(s_86), .O(gate434inter3));
  inv1  gate1153(.a(s_87), .O(gate434inter4));
  nand2 gate1154(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1155(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1156(.a(G1057), .O(gate434inter7));
  inv1  gate1157(.a(G1153), .O(gate434inter8));
  nand2 gate1158(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1159(.a(s_87), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1160(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1161(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1162(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate953(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate954(.a(gate440inter0), .b(s_58), .O(gate440inter1));
  and2  gate955(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate956(.a(s_58), .O(gate440inter3));
  inv1  gate957(.a(s_59), .O(gate440inter4));
  nand2 gate958(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate959(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate960(.a(G1066), .O(gate440inter7));
  inv1  gate961(.a(G1162), .O(gate440inter8));
  nand2 gate962(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate963(.a(s_59), .b(gate440inter3), .O(gate440inter10));
  nor2  gate964(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate965(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate966(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1121(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1122(.a(gate441inter0), .b(s_82), .O(gate441inter1));
  and2  gate1123(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1124(.a(s_82), .O(gate441inter3));
  inv1  gate1125(.a(s_83), .O(gate441inter4));
  nand2 gate1126(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1127(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1128(.a(G12), .O(gate441inter7));
  inv1  gate1129(.a(G1165), .O(gate441inter8));
  nand2 gate1130(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1131(.a(s_83), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1132(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1133(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1134(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1261(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1262(.a(gate446inter0), .b(s_102), .O(gate446inter1));
  and2  gate1263(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1264(.a(s_102), .O(gate446inter3));
  inv1  gate1265(.a(s_103), .O(gate446inter4));
  nand2 gate1266(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1267(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1268(.a(G1075), .O(gate446inter7));
  inv1  gate1269(.a(G1171), .O(gate446inter8));
  nand2 gate1270(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1271(.a(s_103), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1272(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1273(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1274(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate561(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate562(.a(gate448inter0), .b(s_2), .O(gate448inter1));
  and2  gate563(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate564(.a(s_2), .O(gate448inter3));
  inv1  gate565(.a(s_3), .O(gate448inter4));
  nand2 gate566(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate567(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate568(.a(G1078), .O(gate448inter7));
  inv1  gate569(.a(G1174), .O(gate448inter8));
  nand2 gate570(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate571(.a(s_3), .b(gate448inter3), .O(gate448inter10));
  nor2  gate572(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate573(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate574(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate995(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate996(.a(gate452inter0), .b(s_64), .O(gate452inter1));
  and2  gate997(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate998(.a(s_64), .O(gate452inter3));
  inv1  gate999(.a(s_65), .O(gate452inter4));
  nand2 gate1000(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1001(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1002(.a(G1084), .O(gate452inter7));
  inv1  gate1003(.a(G1180), .O(gate452inter8));
  nand2 gate1004(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1005(.a(s_65), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1006(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1007(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1008(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1289(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1290(.a(gate457inter0), .b(s_106), .O(gate457inter1));
  and2  gate1291(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1292(.a(s_106), .O(gate457inter3));
  inv1  gate1293(.a(s_107), .O(gate457inter4));
  nand2 gate1294(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1295(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1296(.a(G20), .O(gate457inter7));
  inv1  gate1297(.a(G1189), .O(gate457inter8));
  nand2 gate1298(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1299(.a(s_107), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1300(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1301(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1302(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate687(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate688(.a(gate458inter0), .b(s_20), .O(gate458inter1));
  and2  gate689(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate690(.a(s_20), .O(gate458inter3));
  inv1  gate691(.a(s_21), .O(gate458inter4));
  nand2 gate692(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate693(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate694(.a(G1093), .O(gate458inter7));
  inv1  gate695(.a(G1189), .O(gate458inter8));
  nand2 gate696(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate697(.a(s_21), .b(gate458inter3), .O(gate458inter10));
  nor2  gate698(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate699(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate700(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1065(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1066(.a(gate459inter0), .b(s_74), .O(gate459inter1));
  and2  gate1067(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1068(.a(s_74), .O(gate459inter3));
  inv1  gate1069(.a(s_75), .O(gate459inter4));
  nand2 gate1070(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1071(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1072(.a(G21), .O(gate459inter7));
  inv1  gate1073(.a(G1192), .O(gate459inter8));
  nand2 gate1074(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1075(.a(s_75), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1076(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1077(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1078(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate547(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate548(.a(gate464inter0), .b(s_0), .O(gate464inter1));
  and2  gate549(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate550(.a(s_0), .O(gate464inter3));
  inv1  gate551(.a(s_1), .O(gate464inter4));
  nand2 gate552(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate553(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate554(.a(G1102), .O(gate464inter7));
  inv1  gate555(.a(G1198), .O(gate464inter8));
  nand2 gate556(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate557(.a(s_1), .b(gate464inter3), .O(gate464inter10));
  nor2  gate558(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate559(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate560(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1863(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1864(.a(gate465inter0), .b(s_188), .O(gate465inter1));
  and2  gate1865(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1866(.a(s_188), .O(gate465inter3));
  inv1  gate1867(.a(s_189), .O(gate465inter4));
  nand2 gate1868(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1869(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1870(.a(G24), .O(gate465inter7));
  inv1  gate1871(.a(G1201), .O(gate465inter8));
  nand2 gate1872(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1873(.a(s_189), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1874(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1875(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1876(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1457(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1458(.a(gate467inter0), .b(s_130), .O(gate467inter1));
  and2  gate1459(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1460(.a(s_130), .O(gate467inter3));
  inv1  gate1461(.a(s_131), .O(gate467inter4));
  nand2 gate1462(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1463(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1464(.a(G25), .O(gate467inter7));
  inv1  gate1465(.a(G1204), .O(gate467inter8));
  nand2 gate1466(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1467(.a(s_131), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1468(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1469(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1470(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate701(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate702(.a(gate472inter0), .b(s_22), .O(gate472inter1));
  and2  gate703(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate704(.a(s_22), .O(gate472inter3));
  inv1  gate705(.a(s_23), .O(gate472inter4));
  nand2 gate706(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate707(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate708(.a(G1114), .O(gate472inter7));
  inv1  gate709(.a(G1210), .O(gate472inter8));
  nand2 gate710(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate711(.a(s_23), .b(gate472inter3), .O(gate472inter10));
  nor2  gate712(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate713(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate714(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1093(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1094(.a(gate474inter0), .b(s_78), .O(gate474inter1));
  and2  gate1095(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1096(.a(s_78), .O(gate474inter3));
  inv1  gate1097(.a(s_79), .O(gate474inter4));
  nand2 gate1098(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1099(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1100(.a(G1117), .O(gate474inter7));
  inv1  gate1101(.a(G1213), .O(gate474inter8));
  nand2 gate1102(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1103(.a(s_79), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1104(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1105(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1106(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate785(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate786(.a(gate482inter0), .b(s_34), .O(gate482inter1));
  and2  gate787(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate788(.a(s_34), .O(gate482inter3));
  inv1  gate789(.a(s_35), .O(gate482inter4));
  nand2 gate790(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate791(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate792(.a(G1129), .O(gate482inter7));
  inv1  gate793(.a(G1225), .O(gate482inter8));
  nand2 gate794(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate795(.a(s_35), .b(gate482inter3), .O(gate482inter10));
  nor2  gate796(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate797(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate798(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1317(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1318(.a(gate492inter0), .b(s_110), .O(gate492inter1));
  and2  gate1319(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1320(.a(s_110), .O(gate492inter3));
  inv1  gate1321(.a(s_111), .O(gate492inter4));
  nand2 gate1322(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1323(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1324(.a(G1246), .O(gate492inter7));
  inv1  gate1325(.a(G1247), .O(gate492inter8));
  nand2 gate1326(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1327(.a(s_111), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1328(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1329(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1330(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1751(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1752(.a(gate504inter0), .b(s_172), .O(gate504inter1));
  and2  gate1753(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1754(.a(s_172), .O(gate504inter3));
  inv1  gate1755(.a(s_173), .O(gate504inter4));
  nand2 gate1756(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1757(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1758(.a(G1270), .O(gate504inter7));
  inv1  gate1759(.a(G1271), .O(gate504inter8));
  nand2 gate1760(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1761(.a(s_173), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1762(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1763(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1764(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate883(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate884(.a(gate510inter0), .b(s_48), .O(gate510inter1));
  and2  gate885(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate886(.a(s_48), .O(gate510inter3));
  inv1  gate887(.a(s_49), .O(gate510inter4));
  nand2 gate888(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate889(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate890(.a(G1282), .O(gate510inter7));
  inv1  gate891(.a(G1283), .O(gate510inter8));
  nand2 gate892(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate893(.a(s_49), .b(gate510inter3), .O(gate510inter10));
  nor2  gate894(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate895(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate896(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule