module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2171(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2172(.a(gate9inter0), .b(s_232), .O(gate9inter1));
  and2  gate2173(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2174(.a(s_232), .O(gate9inter3));
  inv1  gate2175(.a(s_233), .O(gate9inter4));
  nand2 gate2176(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2177(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2178(.a(G1), .O(gate9inter7));
  inv1  gate2179(.a(G2), .O(gate9inter8));
  nand2 gate2180(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2181(.a(s_233), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2182(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2183(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2184(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2997(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2998(.a(gate10inter0), .b(s_350), .O(gate10inter1));
  and2  gate2999(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate3000(.a(s_350), .O(gate10inter3));
  inv1  gate3001(.a(s_351), .O(gate10inter4));
  nand2 gate3002(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate3003(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate3004(.a(G3), .O(gate10inter7));
  inv1  gate3005(.a(G4), .O(gate10inter8));
  nand2 gate3006(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate3007(.a(s_351), .b(gate10inter3), .O(gate10inter10));
  nor2  gate3008(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate3009(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate3010(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate1107(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1108(.a(gate11inter0), .b(s_80), .O(gate11inter1));
  and2  gate1109(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1110(.a(s_80), .O(gate11inter3));
  inv1  gate1111(.a(s_81), .O(gate11inter4));
  nand2 gate1112(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1113(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1114(.a(G5), .O(gate11inter7));
  inv1  gate1115(.a(G6), .O(gate11inter8));
  nand2 gate1116(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1117(.a(s_81), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1118(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1119(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1120(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2619(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2620(.a(gate13inter0), .b(s_296), .O(gate13inter1));
  and2  gate2621(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2622(.a(s_296), .O(gate13inter3));
  inv1  gate2623(.a(s_297), .O(gate13inter4));
  nand2 gate2624(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2625(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2626(.a(G9), .O(gate13inter7));
  inv1  gate2627(.a(G10), .O(gate13inter8));
  nand2 gate2628(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2629(.a(s_297), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2630(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2631(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2632(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1695(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1696(.a(gate15inter0), .b(s_164), .O(gate15inter1));
  and2  gate1697(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1698(.a(s_164), .O(gate15inter3));
  inv1  gate1699(.a(s_165), .O(gate15inter4));
  nand2 gate1700(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1701(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1702(.a(G13), .O(gate15inter7));
  inv1  gate1703(.a(G14), .O(gate15inter8));
  nand2 gate1704(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1705(.a(s_165), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1706(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1707(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1708(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate813(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate814(.a(gate16inter0), .b(s_38), .O(gate16inter1));
  and2  gate815(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate816(.a(s_38), .O(gate16inter3));
  inv1  gate817(.a(s_39), .O(gate16inter4));
  nand2 gate818(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate819(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate820(.a(G15), .O(gate16inter7));
  inv1  gate821(.a(G16), .O(gate16inter8));
  nand2 gate822(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate823(.a(s_39), .b(gate16inter3), .O(gate16inter10));
  nor2  gate824(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate825(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate826(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1163(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1164(.a(gate17inter0), .b(s_88), .O(gate17inter1));
  and2  gate1165(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1166(.a(s_88), .O(gate17inter3));
  inv1  gate1167(.a(s_89), .O(gate17inter4));
  nand2 gate1168(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1169(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1170(.a(G17), .O(gate17inter7));
  inv1  gate1171(.a(G18), .O(gate17inter8));
  nand2 gate1172(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1173(.a(s_89), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1174(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1175(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1176(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1807(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1808(.a(gate18inter0), .b(s_180), .O(gate18inter1));
  and2  gate1809(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1810(.a(s_180), .O(gate18inter3));
  inv1  gate1811(.a(s_181), .O(gate18inter4));
  nand2 gate1812(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1813(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1814(.a(G19), .O(gate18inter7));
  inv1  gate1815(.a(G20), .O(gate18inter8));
  nand2 gate1816(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1817(.a(s_181), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1818(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1819(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1820(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate3039(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate3040(.a(gate21inter0), .b(s_356), .O(gate21inter1));
  and2  gate3041(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate3042(.a(s_356), .O(gate21inter3));
  inv1  gate3043(.a(s_357), .O(gate21inter4));
  nand2 gate3044(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate3045(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate3046(.a(G25), .O(gate21inter7));
  inv1  gate3047(.a(G26), .O(gate21inter8));
  nand2 gate3048(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate3049(.a(s_357), .b(gate21inter3), .O(gate21inter10));
  nor2  gate3050(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate3051(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate3052(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2255(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2256(.a(gate23inter0), .b(s_244), .O(gate23inter1));
  and2  gate2257(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2258(.a(s_244), .O(gate23inter3));
  inv1  gate2259(.a(s_245), .O(gate23inter4));
  nand2 gate2260(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2261(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2262(.a(G29), .O(gate23inter7));
  inv1  gate2263(.a(G30), .O(gate23inter8));
  nand2 gate2264(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2265(.a(s_245), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2266(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2267(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2268(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2311(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2312(.a(gate24inter0), .b(s_252), .O(gate24inter1));
  and2  gate2313(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2314(.a(s_252), .O(gate24inter3));
  inv1  gate2315(.a(s_253), .O(gate24inter4));
  nand2 gate2316(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2317(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2318(.a(G31), .O(gate24inter7));
  inv1  gate2319(.a(G32), .O(gate24inter8));
  nand2 gate2320(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2321(.a(s_253), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2322(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2323(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2324(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1345(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1346(.a(gate27inter0), .b(s_114), .O(gate27inter1));
  and2  gate1347(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1348(.a(s_114), .O(gate27inter3));
  inv1  gate1349(.a(s_115), .O(gate27inter4));
  nand2 gate1350(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1351(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1352(.a(G2), .O(gate27inter7));
  inv1  gate1353(.a(G6), .O(gate27inter8));
  nand2 gate1354(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1355(.a(s_115), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1356(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1357(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1358(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1933(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1934(.a(gate28inter0), .b(s_198), .O(gate28inter1));
  and2  gate1935(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1936(.a(s_198), .O(gate28inter3));
  inv1  gate1937(.a(s_199), .O(gate28inter4));
  nand2 gate1938(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1939(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1940(.a(G10), .O(gate28inter7));
  inv1  gate1941(.a(G14), .O(gate28inter8));
  nand2 gate1942(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1943(.a(s_199), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1944(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1945(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1946(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate3151(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate3152(.a(gate30inter0), .b(s_372), .O(gate30inter1));
  and2  gate3153(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate3154(.a(s_372), .O(gate30inter3));
  inv1  gate3155(.a(s_373), .O(gate30inter4));
  nand2 gate3156(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate3157(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate3158(.a(G11), .O(gate30inter7));
  inv1  gate3159(.a(G15), .O(gate30inter8));
  nand2 gate3160(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate3161(.a(s_373), .b(gate30inter3), .O(gate30inter10));
  nor2  gate3162(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate3163(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate3164(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate2549(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2550(.a(gate31inter0), .b(s_286), .O(gate31inter1));
  and2  gate2551(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2552(.a(s_286), .O(gate31inter3));
  inv1  gate2553(.a(s_287), .O(gate31inter4));
  nand2 gate2554(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2555(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2556(.a(G4), .O(gate31inter7));
  inv1  gate2557(.a(G8), .O(gate31inter8));
  nand2 gate2558(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2559(.a(s_287), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2560(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2561(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2562(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate2759(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2760(.a(gate32inter0), .b(s_316), .O(gate32inter1));
  and2  gate2761(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2762(.a(s_316), .O(gate32inter3));
  inv1  gate2763(.a(s_317), .O(gate32inter4));
  nand2 gate2764(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2765(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2766(.a(G12), .O(gate32inter7));
  inv1  gate2767(.a(G16), .O(gate32inter8));
  nand2 gate2768(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2769(.a(s_317), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2770(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2771(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2772(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1723(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1724(.a(gate35inter0), .b(s_168), .O(gate35inter1));
  and2  gate1725(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1726(.a(s_168), .O(gate35inter3));
  inv1  gate1727(.a(s_169), .O(gate35inter4));
  nand2 gate1728(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1729(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1730(.a(G18), .O(gate35inter7));
  inv1  gate1731(.a(G22), .O(gate35inter8));
  nand2 gate1732(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1733(.a(s_169), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1734(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1735(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1736(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2423(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2424(.a(gate40inter0), .b(s_268), .O(gate40inter1));
  and2  gate2425(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2426(.a(s_268), .O(gate40inter3));
  inv1  gate2427(.a(s_269), .O(gate40inter4));
  nand2 gate2428(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2429(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2430(.a(G28), .O(gate40inter7));
  inv1  gate2431(.a(G32), .O(gate40inter8));
  nand2 gate2432(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2433(.a(s_269), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2434(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2435(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2436(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2843(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2844(.a(gate44inter0), .b(s_328), .O(gate44inter1));
  and2  gate2845(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2846(.a(s_328), .O(gate44inter3));
  inv1  gate2847(.a(s_329), .O(gate44inter4));
  nand2 gate2848(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2849(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2850(.a(G4), .O(gate44inter7));
  inv1  gate2851(.a(G269), .O(gate44inter8));
  nand2 gate2852(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2853(.a(s_329), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2854(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2855(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2856(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate827(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate828(.a(gate45inter0), .b(s_40), .O(gate45inter1));
  and2  gate829(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate830(.a(s_40), .O(gate45inter3));
  inv1  gate831(.a(s_41), .O(gate45inter4));
  nand2 gate832(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate833(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate834(.a(G5), .O(gate45inter7));
  inv1  gate835(.a(G272), .O(gate45inter8));
  nand2 gate836(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate837(.a(s_41), .b(gate45inter3), .O(gate45inter10));
  nor2  gate838(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate839(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate840(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1961(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1962(.a(gate47inter0), .b(s_202), .O(gate47inter1));
  and2  gate1963(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1964(.a(s_202), .O(gate47inter3));
  inv1  gate1965(.a(s_203), .O(gate47inter4));
  nand2 gate1966(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1967(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1968(.a(G7), .O(gate47inter7));
  inv1  gate1969(.a(G275), .O(gate47inter8));
  nand2 gate1970(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1971(.a(s_203), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1972(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1973(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1974(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1079(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1080(.a(gate50inter0), .b(s_76), .O(gate50inter1));
  and2  gate1081(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1082(.a(s_76), .O(gate50inter3));
  inv1  gate1083(.a(s_77), .O(gate50inter4));
  nand2 gate1084(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1085(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1086(.a(G10), .O(gate50inter7));
  inv1  gate1087(.a(G278), .O(gate50inter8));
  nand2 gate1088(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1089(.a(s_77), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1090(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1091(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1092(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1121(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1122(.a(gate51inter0), .b(s_82), .O(gate51inter1));
  and2  gate1123(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1124(.a(s_82), .O(gate51inter3));
  inv1  gate1125(.a(s_83), .O(gate51inter4));
  nand2 gate1126(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1127(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1128(.a(G11), .O(gate51inter7));
  inv1  gate1129(.a(G281), .O(gate51inter8));
  nand2 gate1130(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1131(.a(s_83), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1132(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1133(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1134(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2829(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2830(.a(gate53inter0), .b(s_326), .O(gate53inter1));
  and2  gate2831(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2832(.a(s_326), .O(gate53inter3));
  inv1  gate2833(.a(s_327), .O(gate53inter4));
  nand2 gate2834(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2835(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2836(.a(G13), .O(gate53inter7));
  inv1  gate2837(.a(G284), .O(gate53inter8));
  nand2 gate2838(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2839(.a(s_327), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2840(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2841(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2842(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1331(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1332(.a(gate55inter0), .b(s_112), .O(gate55inter1));
  and2  gate1333(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1334(.a(s_112), .O(gate55inter3));
  inv1  gate1335(.a(s_113), .O(gate55inter4));
  nand2 gate1336(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1337(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1338(.a(G15), .O(gate55inter7));
  inv1  gate1339(.a(G287), .O(gate55inter8));
  nand2 gate1340(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1341(.a(s_113), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1342(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1343(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1344(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2451(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2452(.a(gate56inter0), .b(s_272), .O(gate56inter1));
  and2  gate2453(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2454(.a(s_272), .O(gate56inter3));
  inv1  gate2455(.a(s_273), .O(gate56inter4));
  nand2 gate2456(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2457(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2458(.a(G16), .O(gate56inter7));
  inv1  gate2459(.a(G287), .O(gate56inter8));
  nand2 gate2460(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2461(.a(s_273), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2462(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2463(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2464(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1863(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1864(.a(gate57inter0), .b(s_188), .O(gate57inter1));
  and2  gate1865(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1866(.a(s_188), .O(gate57inter3));
  inv1  gate1867(.a(s_189), .O(gate57inter4));
  nand2 gate1868(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1869(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1870(.a(G17), .O(gate57inter7));
  inv1  gate1871(.a(G290), .O(gate57inter8));
  nand2 gate1872(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1873(.a(s_189), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1874(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1875(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1876(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1569(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1570(.a(gate58inter0), .b(s_146), .O(gate58inter1));
  and2  gate1571(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1572(.a(s_146), .O(gate58inter3));
  inv1  gate1573(.a(s_147), .O(gate58inter4));
  nand2 gate1574(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1575(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1576(.a(G18), .O(gate58inter7));
  inv1  gate1577(.a(G290), .O(gate58inter8));
  nand2 gate1578(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1579(.a(s_147), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1580(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1581(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1582(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate659(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate660(.a(gate60inter0), .b(s_16), .O(gate60inter1));
  and2  gate661(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate662(.a(s_16), .O(gate60inter3));
  inv1  gate663(.a(s_17), .O(gate60inter4));
  nand2 gate664(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate665(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate666(.a(G20), .O(gate60inter7));
  inv1  gate667(.a(G293), .O(gate60inter8));
  nand2 gate668(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate669(.a(s_17), .b(gate60inter3), .O(gate60inter10));
  nor2  gate670(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate671(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate672(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1583(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1584(.a(gate63inter0), .b(s_148), .O(gate63inter1));
  and2  gate1585(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1586(.a(s_148), .O(gate63inter3));
  inv1  gate1587(.a(s_149), .O(gate63inter4));
  nand2 gate1588(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1589(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1590(.a(G23), .O(gate63inter7));
  inv1  gate1591(.a(G299), .O(gate63inter8));
  nand2 gate1592(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1593(.a(s_149), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1594(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1595(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1596(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2479(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2480(.a(gate64inter0), .b(s_276), .O(gate64inter1));
  and2  gate2481(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2482(.a(s_276), .O(gate64inter3));
  inv1  gate2483(.a(s_277), .O(gate64inter4));
  nand2 gate2484(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2485(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2486(.a(G24), .O(gate64inter7));
  inv1  gate2487(.a(G299), .O(gate64inter8));
  nand2 gate2488(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2489(.a(s_277), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2490(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2491(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2492(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1051(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1052(.a(gate66inter0), .b(s_72), .O(gate66inter1));
  and2  gate1053(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1054(.a(s_72), .O(gate66inter3));
  inv1  gate1055(.a(s_73), .O(gate66inter4));
  nand2 gate1056(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1057(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1058(.a(G26), .O(gate66inter7));
  inv1  gate1059(.a(G302), .O(gate66inter8));
  nand2 gate1060(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1061(.a(s_73), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1062(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1063(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1064(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1905(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1906(.a(gate67inter0), .b(s_194), .O(gate67inter1));
  and2  gate1907(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1908(.a(s_194), .O(gate67inter3));
  inv1  gate1909(.a(s_195), .O(gate67inter4));
  nand2 gate1910(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1911(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1912(.a(G27), .O(gate67inter7));
  inv1  gate1913(.a(G305), .O(gate67inter8));
  nand2 gate1914(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1915(.a(s_195), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1916(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1917(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1918(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate855(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate856(.a(gate69inter0), .b(s_44), .O(gate69inter1));
  and2  gate857(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate858(.a(s_44), .O(gate69inter3));
  inv1  gate859(.a(s_45), .O(gate69inter4));
  nand2 gate860(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate861(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate862(.a(G29), .O(gate69inter7));
  inv1  gate863(.a(G308), .O(gate69inter8));
  nand2 gate864(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate865(.a(s_45), .b(gate69inter3), .O(gate69inter10));
  nor2  gate866(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate867(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate868(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate785(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate786(.a(gate71inter0), .b(s_34), .O(gate71inter1));
  and2  gate787(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate788(.a(s_34), .O(gate71inter3));
  inv1  gate789(.a(s_35), .O(gate71inter4));
  nand2 gate790(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate791(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate792(.a(G31), .O(gate71inter7));
  inv1  gate793(.a(G311), .O(gate71inter8));
  nand2 gate794(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate795(.a(s_35), .b(gate71inter3), .O(gate71inter10));
  nor2  gate796(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate797(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate798(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1597(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1598(.a(gate72inter0), .b(s_150), .O(gate72inter1));
  and2  gate1599(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1600(.a(s_150), .O(gate72inter3));
  inv1  gate1601(.a(s_151), .O(gate72inter4));
  nand2 gate1602(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1603(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1604(.a(G32), .O(gate72inter7));
  inv1  gate1605(.a(G311), .O(gate72inter8));
  nand2 gate1606(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1607(.a(s_151), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1608(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1609(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1610(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2367(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2368(.a(gate78inter0), .b(s_260), .O(gate78inter1));
  and2  gate2369(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2370(.a(s_260), .O(gate78inter3));
  inv1  gate2371(.a(s_261), .O(gate78inter4));
  nand2 gate2372(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2373(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2374(.a(G6), .O(gate78inter7));
  inv1  gate2375(.a(G320), .O(gate78inter8));
  nand2 gate2376(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2377(.a(s_261), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2378(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2379(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2380(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1247(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1248(.a(gate82inter0), .b(s_100), .O(gate82inter1));
  and2  gate1249(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1250(.a(s_100), .O(gate82inter3));
  inv1  gate1251(.a(s_101), .O(gate82inter4));
  nand2 gate1252(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1253(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1254(.a(G7), .O(gate82inter7));
  inv1  gate1255(.a(G326), .O(gate82inter8));
  nand2 gate1256(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1257(.a(s_101), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1258(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1259(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1260(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2675(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2676(.a(gate86inter0), .b(s_304), .O(gate86inter1));
  and2  gate2677(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2678(.a(s_304), .O(gate86inter3));
  inv1  gate2679(.a(s_305), .O(gate86inter4));
  nand2 gate2680(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2681(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2682(.a(G8), .O(gate86inter7));
  inv1  gate2683(.a(G332), .O(gate86inter8));
  nand2 gate2684(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2685(.a(s_305), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2686(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2687(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2688(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2087(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2088(.a(gate87inter0), .b(s_220), .O(gate87inter1));
  and2  gate2089(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2090(.a(s_220), .O(gate87inter3));
  inv1  gate2091(.a(s_221), .O(gate87inter4));
  nand2 gate2092(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2093(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2094(.a(G12), .O(gate87inter7));
  inv1  gate2095(.a(G335), .O(gate87inter8));
  nand2 gate2096(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2097(.a(s_221), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2098(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2099(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2100(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate2465(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2466(.a(gate88inter0), .b(s_274), .O(gate88inter1));
  and2  gate2467(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2468(.a(s_274), .O(gate88inter3));
  inv1  gate2469(.a(s_275), .O(gate88inter4));
  nand2 gate2470(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2471(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2472(.a(G16), .O(gate88inter7));
  inv1  gate2473(.a(G335), .O(gate88inter8));
  nand2 gate2474(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2475(.a(s_275), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2476(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2477(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2478(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate953(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate954(.a(gate89inter0), .b(s_58), .O(gate89inter1));
  and2  gate955(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate956(.a(s_58), .O(gate89inter3));
  inv1  gate957(.a(s_59), .O(gate89inter4));
  nand2 gate958(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate959(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate960(.a(G17), .O(gate89inter7));
  inv1  gate961(.a(G338), .O(gate89inter8));
  nand2 gate962(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate963(.a(s_59), .b(gate89inter3), .O(gate89inter10));
  nor2  gate964(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate965(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate966(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1289(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1290(.a(gate91inter0), .b(s_106), .O(gate91inter1));
  and2  gate1291(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1292(.a(s_106), .O(gate91inter3));
  inv1  gate1293(.a(s_107), .O(gate91inter4));
  nand2 gate1294(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1295(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1296(.a(G25), .O(gate91inter7));
  inv1  gate1297(.a(G341), .O(gate91inter8));
  nand2 gate1298(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1299(.a(s_107), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1300(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1301(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1302(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1233(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1234(.a(gate92inter0), .b(s_98), .O(gate92inter1));
  and2  gate1235(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1236(.a(s_98), .O(gate92inter3));
  inv1  gate1237(.a(s_99), .O(gate92inter4));
  nand2 gate1238(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1239(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1240(.a(G29), .O(gate92inter7));
  inv1  gate1241(.a(G341), .O(gate92inter8));
  nand2 gate1242(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1243(.a(s_99), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1244(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1245(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1246(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2129(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2130(.a(gate94inter0), .b(s_226), .O(gate94inter1));
  and2  gate2131(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2132(.a(s_226), .O(gate94inter3));
  inv1  gate2133(.a(s_227), .O(gate94inter4));
  nand2 gate2134(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2135(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2136(.a(G22), .O(gate94inter7));
  inv1  gate2137(.a(G344), .O(gate94inter8));
  nand2 gate2138(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2139(.a(s_227), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2140(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2141(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2142(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate2199(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2200(.a(gate95inter0), .b(s_236), .O(gate95inter1));
  and2  gate2201(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2202(.a(s_236), .O(gate95inter3));
  inv1  gate2203(.a(s_237), .O(gate95inter4));
  nand2 gate2204(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2205(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2206(.a(G26), .O(gate95inter7));
  inv1  gate2207(.a(G347), .O(gate95inter8));
  nand2 gate2208(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2209(.a(s_237), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2210(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2211(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2212(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1359(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1360(.a(gate97inter0), .b(s_116), .O(gate97inter1));
  and2  gate1361(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1362(.a(s_116), .O(gate97inter3));
  inv1  gate1363(.a(s_117), .O(gate97inter4));
  nand2 gate1364(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1365(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1366(.a(G19), .O(gate97inter7));
  inv1  gate1367(.a(G350), .O(gate97inter8));
  nand2 gate1368(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1369(.a(s_117), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1370(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1371(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1372(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2703(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2704(.a(gate99inter0), .b(s_308), .O(gate99inter1));
  and2  gate2705(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2706(.a(s_308), .O(gate99inter3));
  inv1  gate2707(.a(s_309), .O(gate99inter4));
  nand2 gate2708(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2709(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2710(.a(G27), .O(gate99inter7));
  inv1  gate2711(.a(G353), .O(gate99inter8));
  nand2 gate2712(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2713(.a(s_309), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2714(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2715(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2716(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2927(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2928(.a(gate102inter0), .b(s_340), .O(gate102inter1));
  and2  gate2929(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2930(.a(s_340), .O(gate102inter3));
  inv1  gate2931(.a(s_341), .O(gate102inter4));
  nand2 gate2932(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2933(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2934(.a(G24), .O(gate102inter7));
  inv1  gate2935(.a(G356), .O(gate102inter8));
  nand2 gate2936(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2937(.a(s_341), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2938(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2939(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2940(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2395(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2396(.a(gate104inter0), .b(s_264), .O(gate104inter1));
  and2  gate2397(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2398(.a(s_264), .O(gate104inter3));
  inv1  gate2399(.a(s_265), .O(gate104inter4));
  nand2 gate2400(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2401(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2402(.a(G32), .O(gate104inter7));
  inv1  gate2403(.a(G359), .O(gate104inter8));
  nand2 gate2404(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2405(.a(s_265), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2406(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2407(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2408(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1023(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1024(.a(gate106inter0), .b(s_68), .O(gate106inter1));
  and2  gate1025(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1026(.a(s_68), .O(gate106inter3));
  inv1  gate1027(.a(s_69), .O(gate106inter4));
  nand2 gate1028(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1029(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1030(.a(G364), .O(gate106inter7));
  inv1  gate1031(.a(G365), .O(gate106inter8));
  nand2 gate1032(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1033(.a(s_69), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1034(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1035(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1036(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1205(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1206(.a(gate107inter0), .b(s_94), .O(gate107inter1));
  and2  gate1207(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1208(.a(s_94), .O(gate107inter3));
  inv1  gate1209(.a(s_95), .O(gate107inter4));
  nand2 gate1210(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1211(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1212(.a(G366), .O(gate107inter7));
  inv1  gate1213(.a(G367), .O(gate107inter8));
  nand2 gate1214(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1215(.a(s_95), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1216(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1217(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1218(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate2521(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2522(.a(gate108inter0), .b(s_282), .O(gate108inter1));
  and2  gate2523(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2524(.a(s_282), .O(gate108inter3));
  inv1  gate2525(.a(s_283), .O(gate108inter4));
  nand2 gate2526(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2527(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2528(.a(G368), .O(gate108inter7));
  inv1  gate2529(.a(G369), .O(gate108inter8));
  nand2 gate2530(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2531(.a(s_283), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2532(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2533(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2534(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1653(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1654(.a(gate112inter0), .b(s_158), .O(gate112inter1));
  and2  gate1655(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1656(.a(s_158), .O(gate112inter3));
  inv1  gate1657(.a(s_159), .O(gate112inter4));
  nand2 gate1658(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1659(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1660(.a(G376), .O(gate112inter7));
  inv1  gate1661(.a(G377), .O(gate112inter8));
  nand2 gate1662(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1663(.a(s_159), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1664(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1665(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1666(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2227(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2228(.a(gate115inter0), .b(s_240), .O(gate115inter1));
  and2  gate2229(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2230(.a(s_240), .O(gate115inter3));
  inv1  gate2231(.a(s_241), .O(gate115inter4));
  nand2 gate2232(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2233(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2234(.a(G382), .O(gate115inter7));
  inv1  gate2235(.a(G383), .O(gate115inter8));
  nand2 gate2236(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2237(.a(s_241), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2238(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2239(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2240(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2003(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2004(.a(gate117inter0), .b(s_208), .O(gate117inter1));
  and2  gate2005(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2006(.a(s_208), .O(gate117inter3));
  inv1  gate2007(.a(s_209), .O(gate117inter4));
  nand2 gate2008(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2009(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2010(.a(G386), .O(gate117inter7));
  inv1  gate2011(.a(G387), .O(gate117inter8));
  nand2 gate2012(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2013(.a(s_209), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2014(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2015(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2016(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1009(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1010(.a(gate120inter0), .b(s_66), .O(gate120inter1));
  and2  gate1011(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1012(.a(s_66), .O(gate120inter3));
  inv1  gate1013(.a(s_67), .O(gate120inter4));
  nand2 gate1014(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1015(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1016(.a(G392), .O(gate120inter7));
  inv1  gate1017(.a(G393), .O(gate120inter8));
  nand2 gate1018(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1019(.a(s_67), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1020(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1021(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1022(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2241(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2242(.a(gate123inter0), .b(s_242), .O(gate123inter1));
  and2  gate2243(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2244(.a(s_242), .O(gate123inter3));
  inv1  gate2245(.a(s_243), .O(gate123inter4));
  nand2 gate2246(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2247(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2248(.a(G398), .O(gate123inter7));
  inv1  gate2249(.a(G399), .O(gate123inter8));
  nand2 gate2250(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2251(.a(s_243), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2252(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2253(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2254(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2507(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2508(.a(gate125inter0), .b(s_280), .O(gate125inter1));
  and2  gate2509(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2510(.a(s_280), .O(gate125inter3));
  inv1  gate2511(.a(s_281), .O(gate125inter4));
  nand2 gate2512(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2513(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2514(.a(G402), .O(gate125inter7));
  inv1  gate2515(.a(G403), .O(gate125inter8));
  nand2 gate2516(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2517(.a(s_281), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2518(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2519(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2520(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2941(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2942(.a(gate127inter0), .b(s_342), .O(gate127inter1));
  and2  gate2943(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2944(.a(s_342), .O(gate127inter3));
  inv1  gate2945(.a(s_343), .O(gate127inter4));
  nand2 gate2946(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2947(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2948(.a(G406), .O(gate127inter7));
  inv1  gate2949(.a(G407), .O(gate127inter8));
  nand2 gate2950(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2951(.a(s_343), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2952(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2953(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2954(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate561(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate562(.a(gate128inter0), .b(s_2), .O(gate128inter1));
  and2  gate563(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate564(.a(s_2), .O(gate128inter3));
  inv1  gate565(.a(s_3), .O(gate128inter4));
  nand2 gate566(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate567(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate568(.a(G408), .O(gate128inter7));
  inv1  gate569(.a(G409), .O(gate128inter8));
  nand2 gate570(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate571(.a(s_3), .b(gate128inter3), .O(gate128inter10));
  nor2  gate572(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate573(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate574(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2563(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2564(.a(gate135inter0), .b(s_288), .O(gate135inter1));
  and2  gate2565(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2566(.a(s_288), .O(gate135inter3));
  inv1  gate2567(.a(s_289), .O(gate135inter4));
  nand2 gate2568(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2569(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2570(.a(G422), .O(gate135inter7));
  inv1  gate2571(.a(G423), .O(gate135inter8));
  nand2 gate2572(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2573(.a(s_289), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2574(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2575(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2576(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2787(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2788(.a(gate139inter0), .b(s_320), .O(gate139inter1));
  and2  gate2789(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2790(.a(s_320), .O(gate139inter3));
  inv1  gate2791(.a(s_321), .O(gate139inter4));
  nand2 gate2792(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2793(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2794(.a(G438), .O(gate139inter7));
  inv1  gate2795(.a(G441), .O(gate139inter8));
  nand2 gate2796(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2797(.a(s_321), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2798(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2799(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2800(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2045(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2046(.a(gate141inter0), .b(s_214), .O(gate141inter1));
  and2  gate2047(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2048(.a(s_214), .O(gate141inter3));
  inv1  gate2049(.a(s_215), .O(gate141inter4));
  nand2 gate2050(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2051(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2052(.a(G450), .O(gate141inter7));
  inv1  gate2053(.a(G453), .O(gate141inter8));
  nand2 gate2054(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2055(.a(s_215), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2056(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2057(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2058(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate3165(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate3166(.a(gate143inter0), .b(s_374), .O(gate143inter1));
  and2  gate3167(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate3168(.a(s_374), .O(gate143inter3));
  inv1  gate3169(.a(s_375), .O(gate143inter4));
  nand2 gate3170(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate3171(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate3172(.a(G462), .O(gate143inter7));
  inv1  gate3173(.a(G465), .O(gate143inter8));
  nand2 gate3174(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate3175(.a(s_375), .b(gate143inter3), .O(gate143inter10));
  nor2  gate3176(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate3177(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate3178(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1149(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1150(.a(gate144inter0), .b(s_86), .O(gate144inter1));
  and2  gate1151(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1152(.a(s_86), .O(gate144inter3));
  inv1  gate1153(.a(s_87), .O(gate144inter4));
  nand2 gate1154(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1155(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1156(.a(G468), .O(gate144inter7));
  inv1  gate1157(.a(G471), .O(gate144inter8));
  nand2 gate1158(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1159(.a(s_87), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1160(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1161(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1162(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2493(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2494(.a(gate147inter0), .b(s_278), .O(gate147inter1));
  and2  gate2495(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2496(.a(s_278), .O(gate147inter3));
  inv1  gate2497(.a(s_279), .O(gate147inter4));
  nand2 gate2498(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2499(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2500(.a(G486), .O(gate147inter7));
  inv1  gate2501(.a(G489), .O(gate147inter8));
  nand2 gate2502(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2503(.a(s_279), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2504(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2505(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2506(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2381(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2382(.a(gate149inter0), .b(s_262), .O(gate149inter1));
  and2  gate2383(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2384(.a(s_262), .O(gate149inter3));
  inv1  gate2385(.a(s_263), .O(gate149inter4));
  nand2 gate2386(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2387(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2388(.a(G498), .O(gate149inter7));
  inv1  gate2389(.a(G501), .O(gate149inter8));
  nand2 gate2390(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2391(.a(s_263), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2392(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2393(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2394(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1681(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1682(.a(gate150inter0), .b(s_162), .O(gate150inter1));
  and2  gate1683(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1684(.a(s_162), .O(gate150inter3));
  inv1  gate1685(.a(s_163), .O(gate150inter4));
  nand2 gate1686(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1687(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1688(.a(G504), .O(gate150inter7));
  inv1  gate1689(.a(G507), .O(gate150inter8));
  nand2 gate1690(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1691(.a(s_163), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1692(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1693(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1694(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1317(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1318(.a(gate151inter0), .b(s_110), .O(gate151inter1));
  and2  gate1319(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1320(.a(s_110), .O(gate151inter3));
  inv1  gate1321(.a(s_111), .O(gate151inter4));
  nand2 gate1322(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1323(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1324(.a(G510), .O(gate151inter7));
  inv1  gate1325(.a(G513), .O(gate151inter8));
  nand2 gate1326(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1327(.a(s_111), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1328(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1329(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1330(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1303(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1304(.a(gate152inter0), .b(s_108), .O(gate152inter1));
  and2  gate1305(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1306(.a(s_108), .O(gate152inter3));
  inv1  gate1307(.a(s_109), .O(gate152inter4));
  nand2 gate1308(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1309(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1310(.a(G516), .O(gate152inter7));
  inv1  gate1311(.a(G519), .O(gate152inter8));
  nand2 gate1312(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1313(.a(s_109), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1314(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1315(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1316(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2689(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2690(.a(gate156inter0), .b(s_306), .O(gate156inter1));
  and2  gate2691(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2692(.a(s_306), .O(gate156inter3));
  inv1  gate2693(.a(s_307), .O(gate156inter4));
  nand2 gate2694(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2695(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2696(.a(G435), .O(gate156inter7));
  inv1  gate2697(.a(G525), .O(gate156inter8));
  nand2 gate2698(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2699(.a(s_307), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2700(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2701(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2702(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1891(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1892(.a(gate161inter0), .b(s_192), .O(gate161inter1));
  and2  gate1893(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1894(.a(s_192), .O(gate161inter3));
  inv1  gate1895(.a(s_193), .O(gate161inter4));
  nand2 gate1896(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1897(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1898(.a(G450), .O(gate161inter7));
  inv1  gate1899(.a(G534), .O(gate161inter8));
  nand2 gate1900(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1901(.a(s_193), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1902(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1903(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1904(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate743(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate744(.a(gate163inter0), .b(s_28), .O(gate163inter1));
  and2  gate745(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate746(.a(s_28), .O(gate163inter3));
  inv1  gate747(.a(s_29), .O(gate163inter4));
  nand2 gate748(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate749(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate750(.a(G456), .O(gate163inter7));
  inv1  gate751(.a(G537), .O(gate163inter8));
  nand2 gate752(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate753(.a(s_29), .b(gate163inter3), .O(gate163inter10));
  nor2  gate754(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate755(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate756(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1219(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1220(.a(gate165inter0), .b(s_96), .O(gate165inter1));
  and2  gate1221(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1222(.a(s_96), .O(gate165inter3));
  inv1  gate1223(.a(s_97), .O(gate165inter4));
  nand2 gate1224(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1225(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1226(.a(G462), .O(gate165inter7));
  inv1  gate1227(.a(G540), .O(gate165inter8));
  nand2 gate1228(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1229(.a(s_97), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1230(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1231(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1232(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1443(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1444(.a(gate168inter0), .b(s_128), .O(gate168inter1));
  and2  gate1445(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1446(.a(s_128), .O(gate168inter3));
  inv1  gate1447(.a(s_129), .O(gate168inter4));
  nand2 gate1448(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1449(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1450(.a(G471), .O(gate168inter7));
  inv1  gate1451(.a(G543), .O(gate168inter8));
  nand2 gate1452(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1453(.a(s_129), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1454(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1455(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1456(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2801(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2802(.a(gate169inter0), .b(s_322), .O(gate169inter1));
  and2  gate2803(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2804(.a(s_322), .O(gate169inter3));
  inv1  gate2805(.a(s_323), .O(gate169inter4));
  nand2 gate2806(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2807(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2808(.a(G474), .O(gate169inter7));
  inv1  gate2809(.a(G546), .O(gate169inter8));
  nand2 gate2810(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2811(.a(s_323), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2812(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2813(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2814(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2031(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2032(.a(gate171inter0), .b(s_212), .O(gate171inter1));
  and2  gate2033(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2034(.a(s_212), .O(gate171inter3));
  inv1  gate2035(.a(s_213), .O(gate171inter4));
  nand2 gate2036(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2037(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2038(.a(G480), .O(gate171inter7));
  inv1  gate2039(.a(G549), .O(gate171inter8));
  nand2 gate2040(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2041(.a(s_213), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2042(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2043(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2044(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate925(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate926(.a(gate173inter0), .b(s_54), .O(gate173inter1));
  and2  gate927(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate928(.a(s_54), .O(gate173inter3));
  inv1  gate929(.a(s_55), .O(gate173inter4));
  nand2 gate930(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate931(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate932(.a(G486), .O(gate173inter7));
  inv1  gate933(.a(G552), .O(gate173inter8));
  nand2 gate934(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate935(.a(s_55), .b(gate173inter3), .O(gate173inter10));
  nor2  gate936(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate937(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate938(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate3193(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate3194(.a(gate175inter0), .b(s_378), .O(gate175inter1));
  and2  gate3195(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate3196(.a(s_378), .O(gate175inter3));
  inv1  gate3197(.a(s_379), .O(gate175inter4));
  nand2 gate3198(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate3199(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate3200(.a(G492), .O(gate175inter7));
  inv1  gate3201(.a(G555), .O(gate175inter8));
  nand2 gate3202(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate3203(.a(s_379), .b(gate175inter3), .O(gate175inter10));
  nor2  gate3204(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate3205(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate3206(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1975(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1976(.a(gate176inter0), .b(s_204), .O(gate176inter1));
  and2  gate1977(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1978(.a(s_204), .O(gate176inter3));
  inv1  gate1979(.a(s_205), .O(gate176inter4));
  nand2 gate1980(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1981(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1982(.a(G495), .O(gate176inter7));
  inv1  gate1983(.a(G555), .O(gate176inter8));
  nand2 gate1984(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1985(.a(s_205), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1986(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1987(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1988(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate1541(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1542(.a(gate177inter0), .b(s_142), .O(gate177inter1));
  and2  gate1543(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1544(.a(s_142), .O(gate177inter3));
  inv1  gate1545(.a(s_143), .O(gate177inter4));
  nand2 gate1546(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1547(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1548(.a(G498), .O(gate177inter7));
  inv1  gate1549(.a(G558), .O(gate177inter8));
  nand2 gate1550(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1551(.a(s_143), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1552(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1553(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1554(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2017(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2018(.a(gate179inter0), .b(s_210), .O(gate179inter1));
  and2  gate2019(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2020(.a(s_210), .O(gate179inter3));
  inv1  gate2021(.a(s_211), .O(gate179inter4));
  nand2 gate2022(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2023(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2024(.a(G504), .O(gate179inter7));
  inv1  gate2025(.a(G561), .O(gate179inter8));
  nand2 gate2026(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2027(.a(s_211), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2028(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2029(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2030(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1415(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1416(.a(gate181inter0), .b(s_124), .O(gate181inter1));
  and2  gate1417(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1418(.a(s_124), .O(gate181inter3));
  inv1  gate1419(.a(s_125), .O(gate181inter4));
  nand2 gate1420(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1421(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1422(.a(G510), .O(gate181inter7));
  inv1  gate1423(.a(G564), .O(gate181inter8));
  nand2 gate1424(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1425(.a(s_125), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1426(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1427(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1428(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate3123(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate3124(.a(gate182inter0), .b(s_368), .O(gate182inter1));
  and2  gate3125(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate3126(.a(s_368), .O(gate182inter3));
  inv1  gate3127(.a(s_369), .O(gate182inter4));
  nand2 gate3128(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate3129(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate3130(.a(G513), .O(gate182inter7));
  inv1  gate3131(.a(G564), .O(gate182inter8));
  nand2 gate3132(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate3133(.a(s_369), .b(gate182inter3), .O(gate182inter10));
  nor2  gate3134(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate3135(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate3136(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1471(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1472(.a(gate184inter0), .b(s_132), .O(gate184inter1));
  and2  gate1473(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1474(.a(s_132), .O(gate184inter3));
  inv1  gate1475(.a(s_133), .O(gate184inter4));
  nand2 gate1476(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1477(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1478(.a(G519), .O(gate184inter7));
  inv1  gate1479(.a(G567), .O(gate184inter8));
  nand2 gate1480(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1481(.a(s_133), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1482(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1483(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1484(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2059(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2060(.a(gate190inter0), .b(s_216), .O(gate190inter1));
  and2  gate2061(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2062(.a(s_216), .O(gate190inter3));
  inv1  gate2063(.a(s_217), .O(gate190inter4));
  nand2 gate2064(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2065(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2066(.a(G580), .O(gate190inter7));
  inv1  gate2067(.a(G581), .O(gate190inter8));
  nand2 gate2068(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2069(.a(s_217), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2070(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2071(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2072(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2913(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2914(.a(gate193inter0), .b(s_338), .O(gate193inter1));
  and2  gate2915(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2916(.a(s_338), .O(gate193inter3));
  inv1  gate2917(.a(s_339), .O(gate193inter4));
  nand2 gate2918(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2919(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2920(.a(G586), .O(gate193inter7));
  inv1  gate2921(.a(G587), .O(gate193inter8));
  nand2 gate2922(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2923(.a(s_339), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2924(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2925(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2926(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1947(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1948(.a(gate194inter0), .b(s_200), .O(gate194inter1));
  and2  gate1949(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1950(.a(s_200), .O(gate194inter3));
  inv1  gate1951(.a(s_201), .O(gate194inter4));
  nand2 gate1952(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1953(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1954(.a(G588), .O(gate194inter7));
  inv1  gate1955(.a(G589), .O(gate194inter8));
  nand2 gate1956(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1957(.a(s_201), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1958(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1959(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1960(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1611(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1612(.a(gate195inter0), .b(s_152), .O(gate195inter1));
  and2  gate1613(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1614(.a(s_152), .O(gate195inter3));
  inv1  gate1615(.a(s_153), .O(gate195inter4));
  nand2 gate1616(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1617(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1618(.a(G590), .O(gate195inter7));
  inv1  gate1619(.a(G591), .O(gate195inter8));
  nand2 gate1620(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1621(.a(s_153), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1622(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1623(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1624(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1835(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1836(.a(gate200inter0), .b(s_184), .O(gate200inter1));
  and2  gate1837(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1838(.a(s_184), .O(gate200inter3));
  inv1  gate1839(.a(s_185), .O(gate200inter4));
  nand2 gate1840(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1841(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1842(.a(G600), .O(gate200inter7));
  inv1  gate1843(.a(G601), .O(gate200inter8));
  nand2 gate1844(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1845(.a(s_185), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1846(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1847(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1848(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1555(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1556(.a(gate201inter0), .b(s_144), .O(gate201inter1));
  and2  gate1557(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1558(.a(s_144), .O(gate201inter3));
  inv1  gate1559(.a(s_145), .O(gate201inter4));
  nand2 gate1560(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1561(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1562(.a(G602), .O(gate201inter7));
  inv1  gate1563(.a(G607), .O(gate201inter8));
  nand2 gate1564(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1565(.a(s_145), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1566(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1567(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1568(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate911(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate912(.a(gate203inter0), .b(s_52), .O(gate203inter1));
  and2  gate913(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate914(.a(s_52), .O(gate203inter3));
  inv1  gate915(.a(s_53), .O(gate203inter4));
  nand2 gate916(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate917(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate918(.a(G602), .O(gate203inter7));
  inv1  gate919(.a(G612), .O(gate203inter8));
  nand2 gate920(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate921(.a(s_53), .b(gate203inter3), .O(gate203inter10));
  nor2  gate922(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate923(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate924(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1513(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1514(.a(gate204inter0), .b(s_138), .O(gate204inter1));
  and2  gate1515(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1516(.a(s_138), .O(gate204inter3));
  inv1  gate1517(.a(s_139), .O(gate204inter4));
  nand2 gate1518(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1519(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1520(.a(G607), .O(gate204inter7));
  inv1  gate1521(.a(G617), .O(gate204inter8));
  nand2 gate1522(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1523(.a(s_139), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1524(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1525(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1526(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate645(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate646(.a(gate206inter0), .b(s_14), .O(gate206inter1));
  and2  gate647(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate648(.a(s_14), .O(gate206inter3));
  inv1  gate649(.a(s_15), .O(gate206inter4));
  nand2 gate650(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate651(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate652(.a(G632), .O(gate206inter7));
  inv1  gate653(.a(G637), .O(gate206inter8));
  nand2 gate654(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate655(.a(s_15), .b(gate206inter3), .O(gate206inter10));
  nor2  gate656(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate657(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate658(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate799(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate800(.a(gate207inter0), .b(s_36), .O(gate207inter1));
  and2  gate801(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate802(.a(s_36), .O(gate207inter3));
  inv1  gate803(.a(s_37), .O(gate207inter4));
  nand2 gate804(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate805(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate806(.a(G622), .O(gate207inter7));
  inv1  gate807(.a(G632), .O(gate207inter8));
  nand2 gate808(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate809(.a(s_37), .b(gate207inter3), .O(gate207inter10));
  nor2  gate810(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate811(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate812(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate3011(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate3012(.a(gate211inter0), .b(s_352), .O(gate211inter1));
  and2  gate3013(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate3014(.a(s_352), .O(gate211inter3));
  inv1  gate3015(.a(s_353), .O(gate211inter4));
  nand2 gate3016(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate3017(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate3018(.a(G612), .O(gate211inter7));
  inv1  gate3019(.a(G669), .O(gate211inter8));
  nand2 gate3020(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate3021(.a(s_353), .b(gate211inter3), .O(gate211inter10));
  nor2  gate3022(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate3023(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate3024(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2731(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2732(.a(gate218inter0), .b(s_312), .O(gate218inter1));
  and2  gate2733(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2734(.a(s_312), .O(gate218inter3));
  inv1  gate2735(.a(s_313), .O(gate218inter4));
  nand2 gate2736(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2737(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2738(.a(G627), .O(gate218inter7));
  inv1  gate2739(.a(G678), .O(gate218inter8));
  nand2 gate2740(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2741(.a(s_313), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2742(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2743(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2744(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2283(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2284(.a(gate219inter0), .b(s_248), .O(gate219inter1));
  and2  gate2285(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2286(.a(s_248), .O(gate219inter3));
  inv1  gate2287(.a(s_249), .O(gate219inter4));
  nand2 gate2288(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2289(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2290(.a(G632), .O(gate219inter7));
  inv1  gate2291(.a(G681), .O(gate219inter8));
  nand2 gate2292(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2293(.a(s_249), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2294(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2295(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2296(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1261(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1262(.a(gate222inter0), .b(s_102), .O(gate222inter1));
  and2  gate1263(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1264(.a(s_102), .O(gate222inter3));
  inv1  gate1265(.a(s_103), .O(gate222inter4));
  nand2 gate1266(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1267(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1268(.a(G632), .O(gate222inter7));
  inv1  gate1269(.a(G684), .O(gate222inter8));
  nand2 gate1270(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1271(.a(s_103), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1272(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1273(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1274(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1387(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1388(.a(gate224inter0), .b(s_120), .O(gate224inter1));
  and2  gate1389(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1390(.a(s_120), .O(gate224inter3));
  inv1  gate1391(.a(s_121), .O(gate224inter4));
  nand2 gate1392(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1393(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1394(.a(G637), .O(gate224inter7));
  inv1  gate1395(.a(G687), .O(gate224inter8));
  nand2 gate1396(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1397(.a(s_121), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1398(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1399(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1400(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2745(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2746(.a(gate227inter0), .b(s_314), .O(gate227inter1));
  and2  gate2747(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2748(.a(s_314), .O(gate227inter3));
  inv1  gate2749(.a(s_315), .O(gate227inter4));
  nand2 gate2750(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2751(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2752(.a(G694), .O(gate227inter7));
  inv1  gate2753(.a(G695), .O(gate227inter8));
  nand2 gate2754(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2755(.a(s_315), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2756(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2757(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2758(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate687(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate688(.a(gate228inter0), .b(s_20), .O(gate228inter1));
  and2  gate689(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate690(.a(s_20), .O(gate228inter3));
  inv1  gate691(.a(s_21), .O(gate228inter4));
  nand2 gate692(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate693(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate694(.a(G696), .O(gate228inter7));
  inv1  gate695(.a(G697), .O(gate228inter8));
  nand2 gate696(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate697(.a(s_21), .b(gate228inter3), .O(gate228inter10));
  nor2  gate698(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate699(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate700(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2717(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2718(.a(gate231inter0), .b(s_310), .O(gate231inter1));
  and2  gate2719(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2720(.a(s_310), .O(gate231inter3));
  inv1  gate2721(.a(s_311), .O(gate231inter4));
  nand2 gate2722(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2723(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2724(.a(G702), .O(gate231inter7));
  inv1  gate2725(.a(G703), .O(gate231inter8));
  nand2 gate2726(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2727(.a(s_311), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2728(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2729(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2730(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2157(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2158(.a(gate233inter0), .b(s_230), .O(gate233inter1));
  and2  gate2159(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2160(.a(s_230), .O(gate233inter3));
  inv1  gate2161(.a(s_231), .O(gate233inter4));
  nand2 gate2162(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2163(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2164(.a(G242), .O(gate233inter7));
  inv1  gate2165(.a(G718), .O(gate233inter8));
  nand2 gate2166(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2167(.a(s_231), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2168(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2169(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2170(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2899(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2900(.a(gate234inter0), .b(s_336), .O(gate234inter1));
  and2  gate2901(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2902(.a(s_336), .O(gate234inter3));
  inv1  gate2903(.a(s_337), .O(gate234inter4));
  nand2 gate2904(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2905(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2906(.a(G245), .O(gate234inter7));
  inv1  gate2907(.a(G721), .O(gate234inter8));
  nand2 gate2908(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2909(.a(s_337), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2910(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2911(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2912(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1037(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1038(.a(gate235inter0), .b(s_70), .O(gate235inter1));
  and2  gate1039(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1040(.a(s_70), .O(gate235inter3));
  inv1  gate1041(.a(s_71), .O(gate235inter4));
  nand2 gate1042(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1043(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1044(.a(G248), .O(gate235inter7));
  inv1  gate1045(.a(G724), .O(gate235inter8));
  nand2 gate1046(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1047(.a(s_71), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1048(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1049(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1050(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate897(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate898(.a(gate236inter0), .b(s_50), .O(gate236inter1));
  and2  gate899(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate900(.a(s_50), .O(gate236inter3));
  inv1  gate901(.a(s_51), .O(gate236inter4));
  nand2 gate902(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate903(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate904(.a(G251), .O(gate236inter7));
  inv1  gate905(.a(G727), .O(gate236inter8));
  nand2 gate906(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate907(.a(s_51), .b(gate236inter3), .O(gate236inter10));
  nor2  gate908(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate909(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate910(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate575(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate576(.a(gate237inter0), .b(s_4), .O(gate237inter1));
  and2  gate577(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate578(.a(s_4), .O(gate237inter3));
  inv1  gate579(.a(s_5), .O(gate237inter4));
  nand2 gate580(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate581(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate582(.a(G254), .O(gate237inter7));
  inv1  gate583(.a(G706), .O(gate237inter8));
  nand2 gate584(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate585(.a(s_5), .b(gate237inter3), .O(gate237inter10));
  nor2  gate586(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate587(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate588(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2815(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2816(.a(gate239inter0), .b(s_324), .O(gate239inter1));
  and2  gate2817(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2818(.a(s_324), .O(gate239inter3));
  inv1  gate2819(.a(s_325), .O(gate239inter4));
  nand2 gate2820(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2821(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2822(.a(G260), .O(gate239inter7));
  inv1  gate2823(.a(G712), .O(gate239inter8));
  nand2 gate2824(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2825(.a(s_325), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2826(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2827(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2828(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate2969(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2970(.a(gate240inter0), .b(s_346), .O(gate240inter1));
  and2  gate2971(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2972(.a(s_346), .O(gate240inter3));
  inv1  gate2973(.a(s_347), .O(gate240inter4));
  nand2 gate2974(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2975(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2976(.a(G263), .O(gate240inter7));
  inv1  gate2977(.a(G715), .O(gate240inter8));
  nand2 gate2978(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2979(.a(s_347), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2980(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2981(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2982(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate2073(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2074(.a(gate241inter0), .b(s_218), .O(gate241inter1));
  and2  gate2075(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2076(.a(s_218), .O(gate241inter3));
  inv1  gate2077(.a(s_219), .O(gate241inter4));
  nand2 gate2078(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2079(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2080(.a(G242), .O(gate241inter7));
  inv1  gate2081(.a(G730), .O(gate241inter8));
  nand2 gate2082(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2083(.a(s_219), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2084(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2085(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2086(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1667(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1668(.a(gate253inter0), .b(s_160), .O(gate253inter1));
  and2  gate1669(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1670(.a(s_160), .O(gate253inter3));
  inv1  gate1671(.a(s_161), .O(gate253inter4));
  nand2 gate1672(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1673(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1674(.a(G260), .O(gate253inter7));
  inv1  gate1675(.a(G748), .O(gate253inter8));
  nand2 gate1676(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1677(.a(s_161), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1678(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1679(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1680(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1499(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1500(.a(gate255inter0), .b(s_136), .O(gate255inter1));
  and2  gate1501(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1502(.a(s_136), .O(gate255inter3));
  inv1  gate1503(.a(s_137), .O(gate255inter4));
  nand2 gate1504(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1505(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1506(.a(G263), .O(gate255inter7));
  inv1  gate1507(.a(G751), .O(gate255inter8));
  nand2 gate1508(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1509(.a(s_137), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1510(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1511(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1512(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1625(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1626(.a(gate256inter0), .b(s_154), .O(gate256inter1));
  and2  gate1627(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1628(.a(s_154), .O(gate256inter3));
  inv1  gate1629(.a(s_155), .O(gate256inter4));
  nand2 gate1630(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1631(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1632(.a(G715), .O(gate256inter7));
  inv1  gate1633(.a(G751), .O(gate256inter8));
  nand2 gate1634(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1635(.a(s_155), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1636(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1637(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1638(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate2577(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2578(.a(gate257inter0), .b(s_290), .O(gate257inter1));
  and2  gate2579(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2580(.a(s_290), .O(gate257inter3));
  inv1  gate2581(.a(s_291), .O(gate257inter4));
  nand2 gate2582(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2583(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2584(.a(G754), .O(gate257inter7));
  inv1  gate2585(.a(G755), .O(gate257inter8));
  nand2 gate2586(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2587(.a(s_291), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2588(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2589(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2590(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate757(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate758(.a(gate258inter0), .b(s_30), .O(gate258inter1));
  and2  gate759(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate760(.a(s_30), .O(gate258inter3));
  inv1  gate761(.a(s_31), .O(gate258inter4));
  nand2 gate762(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate763(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate764(.a(G756), .O(gate258inter7));
  inv1  gate765(.a(G757), .O(gate258inter8));
  nand2 gate766(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate767(.a(s_31), .b(gate258inter3), .O(gate258inter10));
  nor2  gate768(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate769(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate770(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2353(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2354(.a(gate261inter0), .b(s_258), .O(gate261inter1));
  and2  gate2355(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2356(.a(s_258), .O(gate261inter3));
  inv1  gate2357(.a(s_259), .O(gate261inter4));
  nand2 gate2358(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2359(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2360(.a(G762), .O(gate261inter7));
  inv1  gate2361(.a(G763), .O(gate261inter8));
  nand2 gate2362(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2363(.a(s_259), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2364(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2365(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2366(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate3025(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate3026(.a(gate262inter0), .b(s_354), .O(gate262inter1));
  and2  gate3027(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate3028(.a(s_354), .O(gate262inter3));
  inv1  gate3029(.a(s_355), .O(gate262inter4));
  nand2 gate3030(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate3031(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate3032(.a(G764), .O(gate262inter7));
  inv1  gate3033(.a(G765), .O(gate262inter8));
  nand2 gate3034(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate3035(.a(s_355), .b(gate262inter3), .O(gate262inter10));
  nor2  gate3036(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate3037(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate3038(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate841(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate842(.a(gate263inter0), .b(s_42), .O(gate263inter1));
  and2  gate843(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate844(.a(s_42), .O(gate263inter3));
  inv1  gate845(.a(s_43), .O(gate263inter4));
  nand2 gate846(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate847(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate848(.a(G766), .O(gate263inter7));
  inv1  gate849(.a(G767), .O(gate263inter8));
  nand2 gate850(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate851(.a(s_43), .b(gate263inter3), .O(gate263inter10));
  nor2  gate852(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate853(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate854(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2115(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2116(.a(gate264inter0), .b(s_224), .O(gate264inter1));
  and2  gate2117(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2118(.a(s_224), .O(gate264inter3));
  inv1  gate2119(.a(s_225), .O(gate264inter4));
  nand2 gate2120(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2121(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2122(.a(G768), .O(gate264inter7));
  inv1  gate2123(.a(G769), .O(gate264inter8));
  nand2 gate2124(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2125(.a(s_225), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2126(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2127(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2128(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1457(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1458(.a(gate267inter0), .b(s_130), .O(gate267inter1));
  and2  gate1459(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1460(.a(s_130), .O(gate267inter3));
  inv1  gate1461(.a(s_131), .O(gate267inter4));
  nand2 gate1462(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1463(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1464(.a(G648), .O(gate267inter7));
  inv1  gate1465(.a(G776), .O(gate267inter8));
  nand2 gate1466(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1467(.a(s_131), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1468(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1469(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1470(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate967(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate968(.a(gate268inter0), .b(s_60), .O(gate268inter1));
  and2  gate969(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate970(.a(s_60), .O(gate268inter3));
  inv1  gate971(.a(s_61), .O(gate268inter4));
  nand2 gate972(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate973(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate974(.a(G651), .O(gate268inter7));
  inv1  gate975(.a(G779), .O(gate268inter8));
  nand2 gate976(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate977(.a(s_61), .b(gate268inter3), .O(gate268inter10));
  nor2  gate978(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate979(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate980(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2535(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2536(.a(gate270inter0), .b(s_284), .O(gate270inter1));
  and2  gate2537(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2538(.a(s_284), .O(gate270inter3));
  inv1  gate2539(.a(s_285), .O(gate270inter4));
  nand2 gate2540(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2541(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2542(.a(G657), .O(gate270inter7));
  inv1  gate2543(.a(G785), .O(gate270inter8));
  nand2 gate2544(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2545(.a(s_285), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2546(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2547(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2548(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1751(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1752(.a(gate271inter0), .b(s_172), .O(gate271inter1));
  and2  gate1753(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1754(.a(s_172), .O(gate271inter3));
  inv1  gate1755(.a(s_173), .O(gate271inter4));
  nand2 gate1756(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1757(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1758(.a(G660), .O(gate271inter7));
  inv1  gate1759(.a(G788), .O(gate271inter8));
  nand2 gate1760(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1761(.a(s_173), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1762(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1763(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1764(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate869(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate870(.a(gate277inter0), .b(s_46), .O(gate277inter1));
  and2  gate871(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate872(.a(s_46), .O(gate277inter3));
  inv1  gate873(.a(s_47), .O(gate277inter4));
  nand2 gate874(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate875(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate876(.a(G648), .O(gate277inter7));
  inv1  gate877(.a(G800), .O(gate277inter8));
  nand2 gate878(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate879(.a(s_47), .b(gate277inter3), .O(gate277inter10));
  nor2  gate880(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate881(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate882(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1877(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1878(.a(gate278inter0), .b(s_190), .O(gate278inter1));
  and2  gate1879(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1880(.a(s_190), .O(gate278inter3));
  inv1  gate1881(.a(s_191), .O(gate278inter4));
  nand2 gate1882(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1883(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1884(.a(G776), .O(gate278inter7));
  inv1  gate1885(.a(G800), .O(gate278inter8));
  nand2 gate1886(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1887(.a(s_191), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1888(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1889(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1890(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate2647(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2648(.a(gate279inter0), .b(s_300), .O(gate279inter1));
  and2  gate2649(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2650(.a(s_300), .O(gate279inter3));
  inv1  gate2651(.a(s_301), .O(gate279inter4));
  nand2 gate2652(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2653(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2654(.a(G651), .O(gate279inter7));
  inv1  gate2655(.a(G803), .O(gate279inter8));
  nand2 gate2656(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2657(.a(s_301), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2658(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2659(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2660(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate883(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate884(.a(gate280inter0), .b(s_48), .O(gate280inter1));
  and2  gate885(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate886(.a(s_48), .O(gate280inter3));
  inv1  gate887(.a(s_49), .O(gate280inter4));
  nand2 gate888(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate889(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate890(.a(G779), .O(gate280inter7));
  inv1  gate891(.a(G803), .O(gate280inter8));
  nand2 gate892(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate893(.a(s_49), .b(gate280inter3), .O(gate280inter10));
  nor2  gate894(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate895(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate896(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1093(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1094(.a(gate282inter0), .b(s_78), .O(gate282inter1));
  and2  gate1095(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1096(.a(s_78), .O(gate282inter3));
  inv1  gate1097(.a(s_79), .O(gate282inter4));
  nand2 gate1098(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1099(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1100(.a(G782), .O(gate282inter7));
  inv1  gate1101(.a(G806), .O(gate282inter8));
  nand2 gate1102(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1103(.a(s_79), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1104(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1105(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1106(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2885(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2886(.a(gate285inter0), .b(s_334), .O(gate285inter1));
  and2  gate2887(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2888(.a(s_334), .O(gate285inter3));
  inv1  gate2889(.a(s_335), .O(gate285inter4));
  nand2 gate2890(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2891(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2892(.a(G660), .O(gate285inter7));
  inv1  gate2893(.a(G812), .O(gate285inter8));
  nand2 gate2894(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2895(.a(s_335), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2896(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2897(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2898(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2101(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2102(.a(gate287inter0), .b(s_222), .O(gate287inter1));
  and2  gate2103(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2104(.a(s_222), .O(gate287inter3));
  inv1  gate2105(.a(s_223), .O(gate287inter4));
  nand2 gate2106(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2107(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2108(.a(G663), .O(gate287inter7));
  inv1  gate2109(.a(G815), .O(gate287inter8));
  nand2 gate2110(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2111(.a(s_223), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2112(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2113(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2114(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate2871(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2872(.a(gate288inter0), .b(s_332), .O(gate288inter1));
  and2  gate2873(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2874(.a(s_332), .O(gate288inter3));
  inv1  gate2875(.a(s_333), .O(gate288inter4));
  nand2 gate2876(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2877(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2878(.a(G791), .O(gate288inter7));
  inv1  gate2879(.a(G815), .O(gate288inter8));
  nand2 gate2880(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2881(.a(s_333), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2882(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2883(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2884(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate701(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate702(.a(gate292inter0), .b(s_22), .O(gate292inter1));
  and2  gate703(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate704(.a(s_22), .O(gate292inter3));
  inv1  gate705(.a(s_23), .O(gate292inter4));
  nand2 gate706(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate707(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate708(.a(G824), .O(gate292inter7));
  inv1  gate709(.a(G825), .O(gate292inter8));
  nand2 gate710(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate711(.a(s_23), .b(gate292inter3), .O(gate292inter10));
  nor2  gate712(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate713(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate714(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1849(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1850(.a(gate293inter0), .b(s_186), .O(gate293inter1));
  and2  gate1851(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1852(.a(s_186), .O(gate293inter3));
  inv1  gate1853(.a(s_187), .O(gate293inter4));
  nand2 gate1854(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1855(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1856(.a(G828), .O(gate293inter7));
  inv1  gate1857(.a(G829), .O(gate293inter8));
  nand2 gate1858(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1859(.a(s_187), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1860(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1861(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1862(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate547(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate548(.a(gate294inter0), .b(s_0), .O(gate294inter1));
  and2  gate549(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate550(.a(s_0), .O(gate294inter3));
  inv1  gate551(.a(s_1), .O(gate294inter4));
  nand2 gate552(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate553(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate554(.a(G832), .O(gate294inter7));
  inv1  gate555(.a(G833), .O(gate294inter8));
  nand2 gate556(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate557(.a(s_1), .b(gate294inter3), .O(gate294inter10));
  nor2  gate558(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate559(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate560(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1639(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1640(.a(gate296inter0), .b(s_156), .O(gate296inter1));
  and2  gate1641(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1642(.a(s_156), .O(gate296inter3));
  inv1  gate1643(.a(s_157), .O(gate296inter4));
  nand2 gate1644(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1645(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1646(.a(G826), .O(gate296inter7));
  inv1  gate1647(.a(G827), .O(gate296inter8));
  nand2 gate1648(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1649(.a(s_157), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1650(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1651(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1652(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1485(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1486(.a(gate388inter0), .b(s_134), .O(gate388inter1));
  and2  gate1487(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1488(.a(s_134), .O(gate388inter3));
  inv1  gate1489(.a(s_135), .O(gate388inter4));
  nand2 gate1490(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1491(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1492(.a(G2), .O(gate388inter7));
  inv1  gate1493(.a(G1039), .O(gate388inter8));
  nand2 gate1494(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1495(.a(s_135), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1496(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1497(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1498(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2185(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2186(.a(gate389inter0), .b(s_234), .O(gate389inter1));
  and2  gate2187(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2188(.a(s_234), .O(gate389inter3));
  inv1  gate2189(.a(s_235), .O(gate389inter4));
  nand2 gate2190(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2191(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2192(.a(G3), .O(gate389inter7));
  inv1  gate2193(.a(G1042), .O(gate389inter8));
  nand2 gate2194(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2195(.a(s_235), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2196(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2197(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2198(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate995(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate996(.a(gate390inter0), .b(s_64), .O(gate390inter1));
  and2  gate997(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate998(.a(s_64), .O(gate390inter3));
  inv1  gate999(.a(s_65), .O(gate390inter4));
  nand2 gate1000(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1001(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1002(.a(G4), .O(gate390inter7));
  inv1  gate1003(.a(G1045), .O(gate390inter8));
  nand2 gate1004(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1005(.a(s_65), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1006(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1007(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1008(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1191(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1192(.a(gate391inter0), .b(s_92), .O(gate391inter1));
  and2  gate1193(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1194(.a(s_92), .O(gate391inter3));
  inv1  gate1195(.a(s_93), .O(gate391inter4));
  nand2 gate1196(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1197(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1198(.a(G5), .O(gate391inter7));
  inv1  gate1199(.a(G1048), .O(gate391inter8));
  nand2 gate1200(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1201(.a(s_93), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1202(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1203(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1204(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1989(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1990(.a(gate393inter0), .b(s_206), .O(gate393inter1));
  and2  gate1991(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1992(.a(s_206), .O(gate393inter3));
  inv1  gate1993(.a(s_207), .O(gate393inter4));
  nand2 gate1994(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1995(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1996(.a(G7), .O(gate393inter7));
  inv1  gate1997(.a(G1054), .O(gate393inter8));
  nand2 gate1998(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1999(.a(s_207), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2000(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2001(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2002(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1793(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1794(.a(gate396inter0), .b(s_178), .O(gate396inter1));
  and2  gate1795(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1796(.a(s_178), .O(gate396inter3));
  inv1  gate1797(.a(s_179), .O(gate396inter4));
  nand2 gate1798(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1799(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1800(.a(G10), .O(gate396inter7));
  inv1  gate1801(.a(G1063), .O(gate396inter8));
  nand2 gate1802(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1803(.a(s_179), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1804(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1805(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1806(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2661(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2662(.a(gate398inter0), .b(s_302), .O(gate398inter1));
  and2  gate2663(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2664(.a(s_302), .O(gate398inter3));
  inv1  gate2665(.a(s_303), .O(gate398inter4));
  nand2 gate2666(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2667(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2668(.a(G12), .O(gate398inter7));
  inv1  gate2669(.a(G1069), .O(gate398inter8));
  nand2 gate2670(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2671(.a(s_303), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2672(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2673(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2674(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2269(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2270(.a(gate404inter0), .b(s_246), .O(gate404inter1));
  and2  gate2271(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2272(.a(s_246), .O(gate404inter3));
  inv1  gate2273(.a(s_247), .O(gate404inter4));
  nand2 gate2274(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2275(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2276(.a(G18), .O(gate404inter7));
  inv1  gate2277(.a(G1087), .O(gate404inter8));
  nand2 gate2278(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2279(.a(s_247), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2280(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2281(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2282(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate939(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate940(.a(gate406inter0), .b(s_56), .O(gate406inter1));
  and2  gate941(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate942(.a(s_56), .O(gate406inter3));
  inv1  gate943(.a(s_57), .O(gate406inter4));
  nand2 gate944(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate945(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate946(.a(G20), .O(gate406inter7));
  inv1  gate947(.a(G1093), .O(gate406inter8));
  nand2 gate948(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate949(.a(s_57), .b(gate406inter3), .O(gate406inter10));
  nor2  gate950(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate951(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate952(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1527(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1528(.a(gate408inter0), .b(s_140), .O(gate408inter1));
  and2  gate1529(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1530(.a(s_140), .O(gate408inter3));
  inv1  gate1531(.a(s_141), .O(gate408inter4));
  nand2 gate1532(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1533(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1534(.a(G22), .O(gate408inter7));
  inv1  gate1535(.a(G1099), .O(gate408inter8));
  nand2 gate1536(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1537(.a(s_141), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1538(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1539(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1540(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate3053(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate3054(.a(gate409inter0), .b(s_358), .O(gate409inter1));
  and2  gate3055(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate3056(.a(s_358), .O(gate409inter3));
  inv1  gate3057(.a(s_359), .O(gate409inter4));
  nand2 gate3058(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate3059(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate3060(.a(G23), .O(gate409inter7));
  inv1  gate3061(.a(G1102), .O(gate409inter8));
  nand2 gate3062(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate3063(.a(s_359), .b(gate409inter3), .O(gate409inter10));
  nor2  gate3064(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate3065(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate3066(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2591(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2592(.a(gate411inter0), .b(s_292), .O(gate411inter1));
  and2  gate2593(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2594(.a(s_292), .O(gate411inter3));
  inv1  gate2595(.a(s_293), .O(gate411inter4));
  nand2 gate2596(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2597(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2598(.a(G25), .O(gate411inter7));
  inv1  gate2599(.a(G1108), .O(gate411inter8));
  nand2 gate2600(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2601(.a(s_293), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2602(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2603(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2604(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2983(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2984(.a(gate415inter0), .b(s_348), .O(gate415inter1));
  and2  gate2985(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2986(.a(s_348), .O(gate415inter3));
  inv1  gate2987(.a(s_349), .O(gate415inter4));
  nand2 gate2988(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2989(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2990(.a(G29), .O(gate415inter7));
  inv1  gate2991(.a(G1120), .O(gate415inter8));
  nand2 gate2992(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2993(.a(s_349), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2994(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2995(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2996(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate2773(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2774(.a(gate416inter0), .b(s_318), .O(gate416inter1));
  and2  gate2775(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2776(.a(s_318), .O(gate416inter3));
  inv1  gate2777(.a(s_319), .O(gate416inter4));
  nand2 gate2778(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2779(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2780(.a(G30), .O(gate416inter7));
  inv1  gate2781(.a(G1123), .O(gate416inter8));
  nand2 gate2782(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2783(.a(s_319), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2784(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2785(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2786(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1919(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1920(.a(gate417inter0), .b(s_196), .O(gate417inter1));
  and2  gate1921(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1922(.a(s_196), .O(gate417inter3));
  inv1  gate1923(.a(s_197), .O(gate417inter4));
  nand2 gate1924(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1925(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1926(.a(G31), .O(gate417inter7));
  inv1  gate1927(.a(G1126), .O(gate417inter8));
  nand2 gate1928(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1929(.a(s_197), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1930(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1931(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1932(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate589(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate590(.a(gate418inter0), .b(s_6), .O(gate418inter1));
  and2  gate591(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate592(.a(s_6), .O(gate418inter3));
  inv1  gate593(.a(s_7), .O(gate418inter4));
  nand2 gate594(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate595(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate596(.a(G32), .O(gate418inter7));
  inv1  gate597(.a(G1129), .O(gate418inter8));
  nand2 gate598(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate599(.a(s_7), .b(gate418inter3), .O(gate418inter10));
  nor2  gate600(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate601(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate602(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1821(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1822(.a(gate420inter0), .b(s_182), .O(gate420inter1));
  and2  gate1823(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1824(.a(s_182), .O(gate420inter3));
  inv1  gate1825(.a(s_183), .O(gate420inter4));
  nand2 gate1826(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1827(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1828(.a(G1036), .O(gate420inter7));
  inv1  gate1829(.a(G1132), .O(gate420inter8));
  nand2 gate1830(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1831(.a(s_183), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1832(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1833(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1834(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1779(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1780(.a(gate422inter0), .b(s_176), .O(gate422inter1));
  and2  gate1781(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1782(.a(s_176), .O(gate422inter3));
  inv1  gate1783(.a(s_177), .O(gate422inter4));
  nand2 gate1784(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1785(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1786(.a(G1039), .O(gate422inter7));
  inv1  gate1787(.a(G1135), .O(gate422inter8));
  nand2 gate1788(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1789(.a(s_177), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1790(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1791(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1792(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1765(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1766(.a(gate425inter0), .b(s_174), .O(gate425inter1));
  and2  gate1767(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1768(.a(s_174), .O(gate425inter3));
  inv1  gate1769(.a(s_175), .O(gate425inter4));
  nand2 gate1770(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1771(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1772(.a(G4), .O(gate425inter7));
  inv1  gate1773(.a(G1141), .O(gate425inter8));
  nand2 gate1774(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1775(.a(s_175), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1776(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1777(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1778(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate715(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate716(.a(gate428inter0), .b(s_24), .O(gate428inter1));
  and2  gate717(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate718(.a(s_24), .O(gate428inter3));
  inv1  gate719(.a(s_25), .O(gate428inter4));
  nand2 gate720(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate721(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate722(.a(G1048), .O(gate428inter7));
  inv1  gate723(.a(G1144), .O(gate428inter8));
  nand2 gate724(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate725(.a(s_25), .b(gate428inter3), .O(gate428inter10));
  nor2  gate726(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate727(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate728(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate3109(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate3110(.a(gate434inter0), .b(s_366), .O(gate434inter1));
  and2  gate3111(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate3112(.a(s_366), .O(gate434inter3));
  inv1  gate3113(.a(s_367), .O(gate434inter4));
  nand2 gate3114(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate3115(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate3116(.a(G1057), .O(gate434inter7));
  inv1  gate3117(.a(G1153), .O(gate434inter8));
  nand2 gate3118(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate3119(.a(s_367), .b(gate434inter3), .O(gate434inter10));
  nor2  gate3120(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate3121(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate3122(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate3081(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate3082(.a(gate440inter0), .b(s_362), .O(gate440inter1));
  and2  gate3083(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate3084(.a(s_362), .O(gate440inter3));
  inv1  gate3085(.a(s_363), .O(gate440inter4));
  nand2 gate3086(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate3087(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate3088(.a(G1066), .O(gate440inter7));
  inv1  gate3089(.a(G1162), .O(gate440inter8));
  nand2 gate3090(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate3091(.a(s_363), .b(gate440inter3), .O(gate440inter10));
  nor2  gate3092(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate3093(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate3094(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate3207(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate3208(.a(gate441inter0), .b(s_380), .O(gate441inter1));
  and2  gate3209(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate3210(.a(s_380), .O(gate441inter3));
  inv1  gate3211(.a(s_381), .O(gate441inter4));
  nand2 gate3212(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate3213(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate3214(.a(G12), .O(gate441inter7));
  inv1  gate3215(.a(G1165), .O(gate441inter8));
  nand2 gate3216(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate3217(.a(s_381), .b(gate441inter3), .O(gate441inter10));
  nor2  gate3218(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate3219(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate3220(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1373(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1374(.a(gate445inter0), .b(s_118), .O(gate445inter1));
  and2  gate1375(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1376(.a(s_118), .O(gate445inter3));
  inv1  gate1377(.a(s_119), .O(gate445inter4));
  nand2 gate1378(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1379(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1380(.a(G14), .O(gate445inter7));
  inv1  gate1381(.a(G1171), .O(gate445inter8));
  nand2 gate1382(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1383(.a(s_119), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1384(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1385(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1386(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1401(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1402(.a(gate446inter0), .b(s_122), .O(gate446inter1));
  and2  gate1403(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1404(.a(s_122), .O(gate446inter3));
  inv1  gate1405(.a(s_123), .O(gate446inter4));
  nand2 gate1406(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1407(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1408(.a(G1075), .O(gate446inter7));
  inv1  gate1409(.a(G1171), .O(gate446inter8));
  nand2 gate1410(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1411(.a(s_123), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1412(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1413(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1414(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2857(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2858(.a(gate448inter0), .b(s_330), .O(gate448inter1));
  and2  gate2859(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2860(.a(s_330), .O(gate448inter3));
  inv1  gate2861(.a(s_331), .O(gate448inter4));
  nand2 gate2862(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2863(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2864(.a(G1078), .O(gate448inter7));
  inv1  gate2865(.a(G1174), .O(gate448inter8));
  nand2 gate2866(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2867(.a(s_331), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2868(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2869(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2870(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate729(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate730(.a(gate451inter0), .b(s_26), .O(gate451inter1));
  and2  gate731(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate732(.a(s_26), .O(gate451inter3));
  inv1  gate733(.a(s_27), .O(gate451inter4));
  nand2 gate734(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate735(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate736(.a(G17), .O(gate451inter7));
  inv1  gate737(.a(G1180), .O(gate451inter8));
  nand2 gate738(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate739(.a(s_27), .b(gate451inter3), .O(gate451inter10));
  nor2  gate740(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate741(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate742(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1177(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1178(.a(gate453inter0), .b(s_90), .O(gate453inter1));
  and2  gate1179(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1180(.a(s_90), .O(gate453inter3));
  inv1  gate1181(.a(s_91), .O(gate453inter4));
  nand2 gate1182(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1183(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1184(.a(G18), .O(gate453inter7));
  inv1  gate1185(.a(G1183), .O(gate453inter8));
  nand2 gate1186(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1187(.a(s_91), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1188(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1189(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1190(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate631(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate632(.a(gate455inter0), .b(s_12), .O(gate455inter1));
  and2  gate633(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate634(.a(s_12), .O(gate455inter3));
  inv1  gate635(.a(s_13), .O(gate455inter4));
  nand2 gate636(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate637(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate638(.a(G19), .O(gate455inter7));
  inv1  gate639(.a(G1186), .O(gate455inter8));
  nand2 gate640(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate641(.a(s_13), .b(gate455inter3), .O(gate455inter10));
  nor2  gate642(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate643(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate644(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate2143(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2144(.a(gate456inter0), .b(s_228), .O(gate456inter1));
  and2  gate2145(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2146(.a(s_228), .O(gate456inter3));
  inv1  gate2147(.a(s_229), .O(gate456inter4));
  nand2 gate2148(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2149(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2150(.a(G1090), .O(gate456inter7));
  inv1  gate2151(.a(G1186), .O(gate456inter8));
  nand2 gate2152(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2153(.a(s_229), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2154(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2155(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2156(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate3095(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate3096(.a(gate458inter0), .b(s_364), .O(gate458inter1));
  and2  gate3097(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate3098(.a(s_364), .O(gate458inter3));
  inv1  gate3099(.a(s_365), .O(gate458inter4));
  nand2 gate3100(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate3101(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate3102(.a(G1093), .O(gate458inter7));
  inv1  gate3103(.a(G1189), .O(gate458inter8));
  nand2 gate3104(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate3105(.a(s_365), .b(gate458inter3), .O(gate458inter10));
  nor2  gate3106(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate3107(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate3108(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate617(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate618(.a(gate460inter0), .b(s_10), .O(gate460inter1));
  and2  gate619(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate620(.a(s_10), .O(gate460inter3));
  inv1  gate621(.a(s_11), .O(gate460inter4));
  nand2 gate622(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate623(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate624(.a(G1096), .O(gate460inter7));
  inv1  gate625(.a(G1192), .O(gate460inter8));
  nand2 gate626(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate627(.a(s_11), .b(gate460inter3), .O(gate460inter10));
  nor2  gate628(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate629(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate630(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2605(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2606(.a(gate461inter0), .b(s_294), .O(gate461inter1));
  and2  gate2607(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2608(.a(s_294), .O(gate461inter3));
  inv1  gate2609(.a(s_295), .O(gate461inter4));
  nand2 gate2610(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2611(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2612(.a(G22), .O(gate461inter7));
  inv1  gate2613(.a(G1195), .O(gate461inter8));
  nand2 gate2614(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2615(.a(s_295), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2616(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2617(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2618(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate603(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate604(.a(gate468inter0), .b(s_8), .O(gate468inter1));
  and2  gate605(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate606(.a(s_8), .O(gate468inter3));
  inv1  gate607(.a(s_9), .O(gate468inter4));
  nand2 gate608(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate609(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate610(.a(G1108), .O(gate468inter7));
  inv1  gate611(.a(G1204), .O(gate468inter8));
  nand2 gate612(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate613(.a(s_9), .b(gate468inter3), .O(gate468inter10));
  nor2  gate614(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate615(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate616(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate1429(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1430(.a(gate469inter0), .b(s_126), .O(gate469inter1));
  and2  gate1431(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1432(.a(s_126), .O(gate469inter3));
  inv1  gate1433(.a(s_127), .O(gate469inter4));
  nand2 gate1434(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1435(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1436(.a(G26), .O(gate469inter7));
  inv1  gate1437(.a(G1207), .O(gate469inter8));
  nand2 gate1438(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1439(.a(s_127), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1440(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1441(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1442(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1737(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1738(.a(gate471inter0), .b(s_170), .O(gate471inter1));
  and2  gate1739(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1740(.a(s_170), .O(gate471inter3));
  inv1  gate1741(.a(s_171), .O(gate471inter4));
  nand2 gate1742(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1743(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1744(.a(G27), .O(gate471inter7));
  inv1  gate1745(.a(G1210), .O(gate471inter8));
  nand2 gate1746(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1747(.a(s_171), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1748(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1749(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1750(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2325(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2326(.a(gate472inter0), .b(s_254), .O(gate472inter1));
  and2  gate2327(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2328(.a(s_254), .O(gate472inter3));
  inv1  gate2329(.a(s_255), .O(gate472inter4));
  nand2 gate2330(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2331(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2332(.a(G1114), .O(gate472inter7));
  inv1  gate2333(.a(G1210), .O(gate472inter8));
  nand2 gate2334(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2335(.a(s_255), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2336(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2337(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2338(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate771(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate772(.a(gate477inter0), .b(s_32), .O(gate477inter1));
  and2  gate773(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate774(.a(s_32), .O(gate477inter3));
  inv1  gate775(.a(s_33), .O(gate477inter4));
  nand2 gate776(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate777(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate778(.a(G30), .O(gate477inter7));
  inv1  gate779(.a(G1219), .O(gate477inter8));
  nand2 gate780(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate781(.a(s_33), .b(gate477inter3), .O(gate477inter10));
  nor2  gate782(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate783(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate784(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2633(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2634(.a(gate478inter0), .b(s_298), .O(gate478inter1));
  and2  gate2635(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2636(.a(s_298), .O(gate478inter3));
  inv1  gate2637(.a(s_299), .O(gate478inter4));
  nand2 gate2638(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2639(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2640(.a(G1123), .O(gate478inter7));
  inv1  gate2641(.a(G1219), .O(gate478inter8));
  nand2 gate2642(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2643(.a(s_299), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2644(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2645(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2646(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate673(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate674(.a(gate479inter0), .b(s_18), .O(gate479inter1));
  and2  gate675(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate676(.a(s_18), .O(gate479inter3));
  inv1  gate677(.a(s_19), .O(gate479inter4));
  nand2 gate678(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate679(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate680(.a(G31), .O(gate479inter7));
  inv1  gate681(.a(G1222), .O(gate479inter8));
  nand2 gate682(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate683(.a(s_19), .b(gate479inter3), .O(gate479inter10));
  nor2  gate684(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate685(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate686(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1135(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1136(.a(gate481inter0), .b(s_84), .O(gate481inter1));
  and2  gate1137(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1138(.a(s_84), .O(gate481inter3));
  inv1  gate1139(.a(s_85), .O(gate481inter4));
  nand2 gate1140(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1141(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1142(.a(G32), .O(gate481inter7));
  inv1  gate1143(.a(G1225), .O(gate481inter8));
  nand2 gate1144(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1145(.a(s_85), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1146(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1147(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1148(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate981(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate982(.a(gate482inter0), .b(s_62), .O(gate482inter1));
  and2  gate983(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate984(.a(s_62), .O(gate482inter3));
  inv1  gate985(.a(s_63), .O(gate482inter4));
  nand2 gate986(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate987(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate988(.a(G1129), .O(gate482inter7));
  inv1  gate989(.a(G1225), .O(gate482inter8));
  nand2 gate990(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate991(.a(s_63), .b(gate482inter3), .O(gate482inter10));
  nor2  gate992(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate993(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate994(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1065(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1066(.a(gate485inter0), .b(s_74), .O(gate485inter1));
  and2  gate1067(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1068(.a(s_74), .O(gate485inter3));
  inv1  gate1069(.a(s_75), .O(gate485inter4));
  nand2 gate1070(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1071(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1072(.a(G1232), .O(gate485inter7));
  inv1  gate1073(.a(G1233), .O(gate485inter8));
  nand2 gate1074(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1075(.a(s_75), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1076(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1077(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1078(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate3067(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate3068(.a(gate487inter0), .b(s_360), .O(gate487inter1));
  and2  gate3069(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate3070(.a(s_360), .O(gate487inter3));
  inv1  gate3071(.a(s_361), .O(gate487inter4));
  nand2 gate3072(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate3073(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate3074(.a(G1236), .O(gate487inter7));
  inv1  gate3075(.a(G1237), .O(gate487inter8));
  nand2 gate3076(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate3077(.a(s_361), .b(gate487inter3), .O(gate487inter10));
  nor2  gate3078(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate3079(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate3080(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2437(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2438(.a(gate488inter0), .b(s_270), .O(gate488inter1));
  and2  gate2439(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2440(.a(s_270), .O(gate488inter3));
  inv1  gate2441(.a(s_271), .O(gate488inter4));
  nand2 gate2442(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2443(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2444(.a(G1238), .O(gate488inter7));
  inv1  gate2445(.a(G1239), .O(gate488inter8));
  nand2 gate2446(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2447(.a(s_271), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2448(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2449(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2450(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate2213(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2214(.a(gate489inter0), .b(s_238), .O(gate489inter1));
  and2  gate2215(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2216(.a(s_238), .O(gate489inter3));
  inv1  gate2217(.a(s_239), .O(gate489inter4));
  nand2 gate2218(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2219(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2220(.a(G1240), .O(gate489inter7));
  inv1  gate2221(.a(G1241), .O(gate489inter8));
  nand2 gate2222(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2223(.a(s_239), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2224(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2225(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2226(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate3137(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate3138(.a(gate490inter0), .b(s_370), .O(gate490inter1));
  and2  gate3139(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate3140(.a(s_370), .O(gate490inter3));
  inv1  gate3141(.a(s_371), .O(gate490inter4));
  nand2 gate3142(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate3143(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate3144(.a(G1242), .O(gate490inter7));
  inv1  gate3145(.a(G1243), .O(gate490inter8));
  nand2 gate3146(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate3147(.a(s_371), .b(gate490inter3), .O(gate490inter10));
  nor2  gate3148(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate3149(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate3150(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate3179(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate3180(.a(gate493inter0), .b(s_376), .O(gate493inter1));
  and2  gate3181(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate3182(.a(s_376), .O(gate493inter3));
  inv1  gate3183(.a(s_377), .O(gate493inter4));
  nand2 gate3184(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate3185(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate3186(.a(G1248), .O(gate493inter7));
  inv1  gate3187(.a(G1249), .O(gate493inter8));
  nand2 gate3188(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate3189(.a(s_377), .b(gate493inter3), .O(gate493inter10));
  nor2  gate3190(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate3191(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate3192(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate2297(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2298(.a(gate495inter0), .b(s_250), .O(gate495inter1));
  and2  gate2299(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2300(.a(s_250), .O(gate495inter3));
  inv1  gate2301(.a(s_251), .O(gate495inter4));
  nand2 gate2302(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2303(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2304(.a(G1252), .O(gate495inter7));
  inv1  gate2305(.a(G1253), .O(gate495inter8));
  nand2 gate2306(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2307(.a(s_251), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2308(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2309(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2310(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2339(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2340(.a(gate497inter0), .b(s_256), .O(gate497inter1));
  and2  gate2341(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2342(.a(s_256), .O(gate497inter3));
  inv1  gate2343(.a(s_257), .O(gate497inter4));
  nand2 gate2344(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2345(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2346(.a(G1256), .O(gate497inter7));
  inv1  gate2347(.a(G1257), .O(gate497inter8));
  nand2 gate2348(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2349(.a(s_257), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2350(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2351(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2352(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1709(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1710(.a(gate500inter0), .b(s_166), .O(gate500inter1));
  and2  gate1711(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1712(.a(s_166), .O(gate500inter3));
  inv1  gate1713(.a(s_167), .O(gate500inter4));
  nand2 gate1714(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1715(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1716(.a(G1262), .O(gate500inter7));
  inv1  gate1717(.a(G1263), .O(gate500inter8));
  nand2 gate1718(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1719(.a(s_167), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1720(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1721(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1722(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2409(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2410(.a(gate508inter0), .b(s_266), .O(gate508inter1));
  and2  gate2411(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2412(.a(s_266), .O(gate508inter3));
  inv1  gate2413(.a(s_267), .O(gate508inter4));
  nand2 gate2414(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2415(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2416(.a(G1278), .O(gate508inter7));
  inv1  gate2417(.a(G1279), .O(gate508inter8));
  nand2 gate2418(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2419(.a(s_267), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2420(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2421(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2422(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1275(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1276(.a(gate510inter0), .b(s_104), .O(gate510inter1));
  and2  gate1277(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1278(.a(s_104), .O(gate510inter3));
  inv1  gate1279(.a(s_105), .O(gate510inter4));
  nand2 gate1280(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1281(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1282(.a(G1282), .O(gate510inter7));
  inv1  gate1283(.a(G1283), .O(gate510inter8));
  nand2 gate1284(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1285(.a(s_105), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1286(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1287(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1288(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2955(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2956(.a(gate514inter0), .b(s_344), .O(gate514inter1));
  and2  gate2957(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2958(.a(s_344), .O(gate514inter3));
  inv1  gate2959(.a(s_345), .O(gate514inter4));
  nand2 gate2960(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2961(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2962(.a(G1290), .O(gate514inter7));
  inv1  gate2963(.a(G1291), .O(gate514inter8));
  nand2 gate2964(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2965(.a(s_345), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2966(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2967(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2968(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule