module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate729(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate730(.a(gate10inter0), .b(s_26), .O(gate10inter1));
  and2  gate731(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate732(.a(s_26), .O(gate10inter3));
  inv1  gate733(.a(s_27), .O(gate10inter4));
  nand2 gate734(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate735(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate736(.a(G3), .O(gate10inter7));
  inv1  gate737(.a(G4), .O(gate10inter8));
  nand2 gate738(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate739(.a(s_27), .b(gate10inter3), .O(gate10inter10));
  nor2  gate740(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate741(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate742(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate1387(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1388(.a(gate11inter0), .b(s_120), .O(gate11inter1));
  and2  gate1389(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1390(.a(s_120), .O(gate11inter3));
  inv1  gate1391(.a(s_121), .O(gate11inter4));
  nand2 gate1392(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1393(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1394(.a(G5), .O(gate11inter7));
  inv1  gate1395(.a(G6), .O(gate11inter8));
  nand2 gate1396(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1397(.a(s_121), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1398(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1399(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1400(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate659(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate660(.a(gate13inter0), .b(s_16), .O(gate13inter1));
  and2  gate661(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate662(.a(s_16), .O(gate13inter3));
  inv1  gate663(.a(s_17), .O(gate13inter4));
  nand2 gate664(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate665(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate666(.a(G9), .O(gate13inter7));
  inv1  gate667(.a(G10), .O(gate13inter8));
  nand2 gate668(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate669(.a(s_17), .b(gate13inter3), .O(gate13inter10));
  nor2  gate670(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate671(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate672(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate799(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate800(.a(gate14inter0), .b(s_36), .O(gate14inter1));
  and2  gate801(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate802(.a(s_36), .O(gate14inter3));
  inv1  gate803(.a(s_37), .O(gate14inter4));
  nand2 gate804(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate805(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate806(.a(G11), .O(gate14inter7));
  inv1  gate807(.a(G12), .O(gate14inter8));
  nand2 gate808(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate809(.a(s_37), .b(gate14inter3), .O(gate14inter10));
  nor2  gate810(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate811(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate812(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1289(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1290(.a(gate16inter0), .b(s_106), .O(gate16inter1));
  and2  gate1291(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1292(.a(s_106), .O(gate16inter3));
  inv1  gate1293(.a(s_107), .O(gate16inter4));
  nand2 gate1294(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1295(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1296(.a(G15), .O(gate16inter7));
  inv1  gate1297(.a(G16), .O(gate16inter8));
  nand2 gate1298(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1299(.a(s_107), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1300(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1301(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1302(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate673(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate674(.a(gate17inter0), .b(s_18), .O(gate17inter1));
  and2  gate675(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate676(.a(s_18), .O(gate17inter3));
  inv1  gate677(.a(s_19), .O(gate17inter4));
  nand2 gate678(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate679(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate680(.a(G17), .O(gate17inter7));
  inv1  gate681(.a(G18), .O(gate17inter8));
  nand2 gate682(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate683(.a(s_19), .b(gate17inter3), .O(gate17inter10));
  nor2  gate684(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate685(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate686(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate953(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate954(.a(gate20inter0), .b(s_58), .O(gate20inter1));
  and2  gate955(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate956(.a(s_58), .O(gate20inter3));
  inv1  gate957(.a(s_59), .O(gate20inter4));
  nand2 gate958(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate959(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate960(.a(G23), .O(gate20inter7));
  inv1  gate961(.a(G24), .O(gate20inter8));
  nand2 gate962(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate963(.a(s_59), .b(gate20inter3), .O(gate20inter10));
  nor2  gate964(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate965(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate966(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1135(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1136(.a(gate22inter0), .b(s_84), .O(gate22inter1));
  and2  gate1137(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1138(.a(s_84), .O(gate22inter3));
  inv1  gate1139(.a(s_85), .O(gate22inter4));
  nand2 gate1140(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1141(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1142(.a(G27), .O(gate22inter7));
  inv1  gate1143(.a(G28), .O(gate22inter8));
  nand2 gate1144(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1145(.a(s_85), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1146(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1147(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1148(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate939(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate940(.a(gate34inter0), .b(s_56), .O(gate34inter1));
  and2  gate941(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate942(.a(s_56), .O(gate34inter3));
  inv1  gate943(.a(s_57), .O(gate34inter4));
  nand2 gate944(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate945(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate946(.a(G25), .O(gate34inter7));
  inv1  gate947(.a(G29), .O(gate34inter8));
  nand2 gate948(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate949(.a(s_57), .b(gate34inter3), .O(gate34inter10));
  nor2  gate950(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate951(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate952(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate827(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate828(.a(gate43inter0), .b(s_40), .O(gate43inter1));
  and2  gate829(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate830(.a(s_40), .O(gate43inter3));
  inv1  gate831(.a(s_41), .O(gate43inter4));
  nand2 gate832(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate833(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate834(.a(G3), .O(gate43inter7));
  inv1  gate835(.a(G269), .O(gate43inter8));
  nand2 gate836(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate837(.a(s_41), .b(gate43inter3), .O(gate43inter10));
  nor2  gate838(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate839(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate840(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1107(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1108(.a(gate44inter0), .b(s_80), .O(gate44inter1));
  and2  gate1109(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1110(.a(s_80), .O(gate44inter3));
  inv1  gate1111(.a(s_81), .O(gate44inter4));
  nand2 gate1112(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1113(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1114(.a(G4), .O(gate44inter7));
  inv1  gate1115(.a(G269), .O(gate44inter8));
  nand2 gate1116(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1117(.a(s_81), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1118(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1119(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1120(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate715(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate716(.a(gate55inter0), .b(s_24), .O(gate55inter1));
  and2  gate717(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate718(.a(s_24), .O(gate55inter3));
  inv1  gate719(.a(s_25), .O(gate55inter4));
  nand2 gate720(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate721(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate722(.a(G15), .O(gate55inter7));
  inv1  gate723(.a(G287), .O(gate55inter8));
  nand2 gate724(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate725(.a(s_25), .b(gate55inter3), .O(gate55inter10));
  nor2  gate726(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate727(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate728(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate687(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate688(.a(gate66inter0), .b(s_20), .O(gate66inter1));
  and2  gate689(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate690(.a(s_20), .O(gate66inter3));
  inv1  gate691(.a(s_21), .O(gate66inter4));
  nand2 gate692(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate693(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate694(.a(G26), .O(gate66inter7));
  inv1  gate695(.a(G302), .O(gate66inter8));
  nand2 gate696(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate697(.a(s_21), .b(gate66inter3), .O(gate66inter10));
  nor2  gate698(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate699(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate700(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate785(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate786(.a(gate67inter0), .b(s_34), .O(gate67inter1));
  and2  gate787(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate788(.a(s_34), .O(gate67inter3));
  inv1  gate789(.a(s_35), .O(gate67inter4));
  nand2 gate790(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate791(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate792(.a(G27), .O(gate67inter7));
  inv1  gate793(.a(G305), .O(gate67inter8));
  nand2 gate794(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate795(.a(s_35), .b(gate67inter3), .O(gate67inter10));
  nor2  gate796(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate797(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate798(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1317(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1318(.a(gate68inter0), .b(s_110), .O(gate68inter1));
  and2  gate1319(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1320(.a(s_110), .O(gate68inter3));
  inv1  gate1321(.a(s_111), .O(gate68inter4));
  nand2 gate1322(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1323(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1324(.a(G28), .O(gate68inter7));
  inv1  gate1325(.a(G305), .O(gate68inter8));
  nand2 gate1326(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1327(.a(s_111), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1328(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1329(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1330(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate897(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate898(.a(gate69inter0), .b(s_50), .O(gate69inter1));
  and2  gate899(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate900(.a(s_50), .O(gate69inter3));
  inv1  gate901(.a(s_51), .O(gate69inter4));
  nand2 gate902(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate903(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate904(.a(G29), .O(gate69inter7));
  inv1  gate905(.a(G308), .O(gate69inter8));
  nand2 gate906(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate907(.a(s_51), .b(gate69inter3), .O(gate69inter10));
  nor2  gate908(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate909(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate910(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1233(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1234(.a(gate71inter0), .b(s_98), .O(gate71inter1));
  and2  gate1235(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1236(.a(s_98), .O(gate71inter3));
  inv1  gate1237(.a(s_99), .O(gate71inter4));
  nand2 gate1238(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1239(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1240(.a(G31), .O(gate71inter7));
  inv1  gate1241(.a(G311), .O(gate71inter8));
  nand2 gate1242(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1243(.a(s_99), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1244(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1245(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1246(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate561(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate562(.a(gate103inter0), .b(s_2), .O(gate103inter1));
  and2  gate563(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate564(.a(s_2), .O(gate103inter3));
  inv1  gate565(.a(s_3), .O(gate103inter4));
  nand2 gate566(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate567(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate568(.a(G28), .O(gate103inter7));
  inv1  gate569(.a(G359), .O(gate103inter8));
  nand2 gate570(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate571(.a(s_3), .b(gate103inter3), .O(gate103inter10));
  nor2  gate572(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate573(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate574(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate757(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate758(.a(gate119inter0), .b(s_30), .O(gate119inter1));
  and2  gate759(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate760(.a(s_30), .O(gate119inter3));
  inv1  gate761(.a(s_31), .O(gate119inter4));
  nand2 gate762(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate763(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate764(.a(G390), .O(gate119inter7));
  inv1  gate765(.a(G391), .O(gate119inter8));
  nand2 gate766(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate767(.a(s_31), .b(gate119inter3), .O(gate119inter10));
  nor2  gate768(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate769(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate770(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1023(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1024(.a(gate120inter0), .b(s_68), .O(gate120inter1));
  and2  gate1025(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1026(.a(s_68), .O(gate120inter3));
  inv1  gate1027(.a(s_69), .O(gate120inter4));
  nand2 gate1028(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1029(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1030(.a(G392), .O(gate120inter7));
  inv1  gate1031(.a(G393), .O(gate120inter8));
  nand2 gate1032(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1033(.a(s_69), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1034(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1035(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1036(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1261(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1262(.a(gate126inter0), .b(s_102), .O(gate126inter1));
  and2  gate1263(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1264(.a(s_102), .O(gate126inter3));
  inv1  gate1265(.a(s_103), .O(gate126inter4));
  nand2 gate1266(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1267(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1268(.a(G404), .O(gate126inter7));
  inv1  gate1269(.a(G405), .O(gate126inter8));
  nand2 gate1270(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1271(.a(s_103), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1272(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1273(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1274(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1359(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1360(.a(gate132inter0), .b(s_116), .O(gate132inter1));
  and2  gate1361(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1362(.a(s_116), .O(gate132inter3));
  inv1  gate1363(.a(s_117), .O(gate132inter4));
  nand2 gate1364(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1365(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1366(.a(G416), .O(gate132inter7));
  inv1  gate1367(.a(G417), .O(gate132inter8));
  nand2 gate1368(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1369(.a(s_117), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1370(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1371(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1372(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate603(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate604(.a(gate140inter0), .b(s_8), .O(gate140inter1));
  and2  gate605(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate606(.a(s_8), .O(gate140inter3));
  inv1  gate607(.a(s_9), .O(gate140inter4));
  nand2 gate608(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate609(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate610(.a(G444), .O(gate140inter7));
  inv1  gate611(.a(G447), .O(gate140inter8));
  nand2 gate612(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate613(.a(s_9), .b(gate140inter3), .O(gate140inter10));
  nor2  gate614(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate615(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate616(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1205(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1206(.a(gate146inter0), .b(s_94), .O(gate146inter1));
  and2  gate1207(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1208(.a(s_94), .O(gate146inter3));
  inv1  gate1209(.a(s_95), .O(gate146inter4));
  nand2 gate1210(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1211(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1212(.a(G480), .O(gate146inter7));
  inv1  gate1213(.a(G483), .O(gate146inter8));
  nand2 gate1214(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1215(.a(s_95), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1216(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1217(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1218(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1177(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1178(.a(gate157inter0), .b(s_90), .O(gate157inter1));
  and2  gate1179(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1180(.a(s_90), .O(gate157inter3));
  inv1  gate1181(.a(s_91), .O(gate157inter4));
  nand2 gate1182(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1183(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1184(.a(G438), .O(gate157inter7));
  inv1  gate1185(.a(G528), .O(gate157inter8));
  nand2 gate1186(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1187(.a(s_91), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1188(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1189(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1190(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate645(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate646(.a(gate161inter0), .b(s_14), .O(gate161inter1));
  and2  gate647(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate648(.a(s_14), .O(gate161inter3));
  inv1  gate649(.a(s_15), .O(gate161inter4));
  nand2 gate650(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate651(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate652(.a(G450), .O(gate161inter7));
  inv1  gate653(.a(G534), .O(gate161inter8));
  nand2 gate654(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate655(.a(s_15), .b(gate161inter3), .O(gate161inter10));
  nor2  gate656(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate657(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate658(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1331(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1332(.a(gate164inter0), .b(s_112), .O(gate164inter1));
  and2  gate1333(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1334(.a(s_112), .O(gate164inter3));
  inv1  gate1335(.a(s_113), .O(gate164inter4));
  nand2 gate1336(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1337(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1338(.a(G459), .O(gate164inter7));
  inv1  gate1339(.a(G537), .O(gate164inter8));
  nand2 gate1340(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1341(.a(s_113), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1342(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1343(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1344(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate813(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate814(.a(gate165inter0), .b(s_38), .O(gate165inter1));
  and2  gate815(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate816(.a(s_38), .O(gate165inter3));
  inv1  gate817(.a(s_39), .O(gate165inter4));
  nand2 gate818(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate819(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate820(.a(G462), .O(gate165inter7));
  inv1  gate821(.a(G540), .O(gate165inter8));
  nand2 gate822(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate823(.a(s_39), .b(gate165inter3), .O(gate165inter10));
  nor2  gate824(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate825(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate826(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate743(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate744(.a(gate166inter0), .b(s_28), .O(gate166inter1));
  and2  gate745(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate746(.a(s_28), .O(gate166inter3));
  inv1  gate747(.a(s_29), .O(gate166inter4));
  nand2 gate748(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate749(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate750(.a(G465), .O(gate166inter7));
  inv1  gate751(.a(G540), .O(gate166inter8));
  nand2 gate752(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate753(.a(s_29), .b(gate166inter3), .O(gate166inter10));
  nor2  gate754(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate755(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate756(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1163(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1164(.a(gate172inter0), .b(s_88), .O(gate172inter1));
  and2  gate1165(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1166(.a(s_88), .O(gate172inter3));
  inv1  gate1167(.a(s_89), .O(gate172inter4));
  nand2 gate1168(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1169(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1170(.a(G483), .O(gate172inter7));
  inv1  gate1171(.a(G549), .O(gate172inter8));
  nand2 gate1172(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1173(.a(s_89), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1174(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1175(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1176(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1247(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1248(.a(gate185inter0), .b(s_100), .O(gate185inter1));
  and2  gate1249(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1250(.a(s_100), .O(gate185inter3));
  inv1  gate1251(.a(s_101), .O(gate185inter4));
  nand2 gate1252(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1253(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1254(.a(G570), .O(gate185inter7));
  inv1  gate1255(.a(G571), .O(gate185inter8));
  nand2 gate1256(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1257(.a(s_101), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1258(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1259(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1260(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate631(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate632(.a(gate193inter0), .b(s_12), .O(gate193inter1));
  and2  gate633(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate634(.a(s_12), .O(gate193inter3));
  inv1  gate635(.a(s_13), .O(gate193inter4));
  nand2 gate636(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate637(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate638(.a(G586), .O(gate193inter7));
  inv1  gate639(.a(G587), .O(gate193inter8));
  nand2 gate640(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate641(.a(s_13), .b(gate193inter3), .O(gate193inter10));
  nor2  gate642(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate643(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate644(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate701(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate702(.a(gate200inter0), .b(s_22), .O(gate200inter1));
  and2  gate703(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate704(.a(s_22), .O(gate200inter3));
  inv1  gate705(.a(s_23), .O(gate200inter4));
  nand2 gate706(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate707(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate708(.a(G600), .O(gate200inter7));
  inv1  gate709(.a(G601), .O(gate200inter8));
  nand2 gate710(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate711(.a(s_23), .b(gate200inter3), .O(gate200inter10));
  nor2  gate712(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate713(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate714(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1121(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1122(.a(gate205inter0), .b(s_82), .O(gate205inter1));
  and2  gate1123(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1124(.a(s_82), .O(gate205inter3));
  inv1  gate1125(.a(s_83), .O(gate205inter4));
  nand2 gate1126(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1127(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1128(.a(G622), .O(gate205inter7));
  inv1  gate1129(.a(G627), .O(gate205inter8));
  nand2 gate1130(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1131(.a(s_83), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1132(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1133(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1134(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1345(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1346(.a(gate233inter0), .b(s_114), .O(gate233inter1));
  and2  gate1347(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1348(.a(s_114), .O(gate233inter3));
  inv1  gate1349(.a(s_115), .O(gate233inter4));
  nand2 gate1350(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1351(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1352(.a(G242), .O(gate233inter7));
  inv1  gate1353(.a(G718), .O(gate233inter8));
  nand2 gate1354(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1355(.a(s_115), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1356(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1357(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1358(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1373(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1374(.a(gate240inter0), .b(s_118), .O(gate240inter1));
  and2  gate1375(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1376(.a(s_118), .O(gate240inter3));
  inv1  gate1377(.a(s_119), .O(gate240inter4));
  nand2 gate1378(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1379(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1380(.a(G263), .O(gate240inter7));
  inv1  gate1381(.a(G715), .O(gate240inter8));
  nand2 gate1382(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1383(.a(s_119), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1384(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1385(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1386(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate617(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate618(.a(gate241inter0), .b(s_10), .O(gate241inter1));
  and2  gate619(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate620(.a(s_10), .O(gate241inter3));
  inv1  gate621(.a(s_11), .O(gate241inter4));
  nand2 gate622(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate623(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate624(.a(G242), .O(gate241inter7));
  inv1  gate625(.a(G730), .O(gate241inter8));
  nand2 gate626(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate627(.a(s_11), .b(gate241inter3), .O(gate241inter10));
  nor2  gate628(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate629(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate630(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1219(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1220(.a(gate267inter0), .b(s_96), .O(gate267inter1));
  and2  gate1221(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1222(.a(s_96), .O(gate267inter3));
  inv1  gate1223(.a(s_97), .O(gate267inter4));
  nand2 gate1224(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1225(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1226(.a(G648), .O(gate267inter7));
  inv1  gate1227(.a(G776), .O(gate267inter8));
  nand2 gate1228(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1229(.a(s_97), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1230(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1231(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1232(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1149(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1150(.a(gate275inter0), .b(s_86), .O(gate275inter1));
  and2  gate1151(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1152(.a(s_86), .O(gate275inter3));
  inv1  gate1153(.a(s_87), .O(gate275inter4));
  nand2 gate1154(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1155(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1156(.a(G645), .O(gate275inter7));
  inv1  gate1157(.a(G797), .O(gate275inter8));
  nand2 gate1158(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1159(.a(s_87), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1160(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1161(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1162(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate883(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate884(.a(gate286inter0), .b(s_48), .O(gate286inter1));
  and2  gate885(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate886(.a(s_48), .O(gate286inter3));
  inv1  gate887(.a(s_49), .O(gate286inter4));
  nand2 gate888(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate889(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate890(.a(G788), .O(gate286inter7));
  inv1  gate891(.a(G812), .O(gate286inter8));
  nand2 gate892(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate893(.a(s_49), .b(gate286inter3), .O(gate286inter10));
  nor2  gate894(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate895(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate896(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate841(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate842(.a(gate296inter0), .b(s_42), .O(gate296inter1));
  and2  gate843(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate844(.a(s_42), .O(gate296inter3));
  inv1  gate845(.a(s_43), .O(gate296inter4));
  nand2 gate846(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate847(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate848(.a(G826), .O(gate296inter7));
  inv1  gate849(.a(G827), .O(gate296inter8));
  nand2 gate850(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate851(.a(s_43), .b(gate296inter3), .O(gate296inter10));
  nor2  gate852(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate853(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate854(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate855(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate856(.a(gate395inter0), .b(s_44), .O(gate395inter1));
  and2  gate857(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate858(.a(s_44), .O(gate395inter3));
  inv1  gate859(.a(s_45), .O(gate395inter4));
  nand2 gate860(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate861(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate862(.a(G9), .O(gate395inter7));
  inv1  gate863(.a(G1060), .O(gate395inter8));
  nand2 gate864(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate865(.a(s_45), .b(gate395inter3), .O(gate395inter10));
  nor2  gate866(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate867(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate868(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1037(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1038(.a(gate396inter0), .b(s_70), .O(gate396inter1));
  and2  gate1039(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1040(.a(s_70), .O(gate396inter3));
  inv1  gate1041(.a(s_71), .O(gate396inter4));
  nand2 gate1042(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1043(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1044(.a(G10), .O(gate396inter7));
  inv1  gate1045(.a(G1063), .O(gate396inter8));
  nand2 gate1046(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1047(.a(s_71), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1048(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1049(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1050(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate925(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate926(.a(gate409inter0), .b(s_54), .O(gate409inter1));
  and2  gate927(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate928(.a(s_54), .O(gate409inter3));
  inv1  gate929(.a(s_55), .O(gate409inter4));
  nand2 gate930(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate931(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate932(.a(G23), .O(gate409inter7));
  inv1  gate933(.a(G1102), .O(gate409inter8));
  nand2 gate934(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate935(.a(s_55), .b(gate409inter3), .O(gate409inter10));
  nor2  gate936(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate937(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate938(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate995(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate996(.a(gate411inter0), .b(s_64), .O(gate411inter1));
  and2  gate997(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate998(.a(s_64), .O(gate411inter3));
  inv1  gate999(.a(s_65), .O(gate411inter4));
  nand2 gate1000(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1001(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1002(.a(G25), .O(gate411inter7));
  inv1  gate1003(.a(G1108), .O(gate411inter8));
  nand2 gate1004(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1005(.a(s_65), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1006(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1007(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1008(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1051(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1052(.a(gate415inter0), .b(s_72), .O(gate415inter1));
  and2  gate1053(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1054(.a(s_72), .O(gate415inter3));
  inv1  gate1055(.a(s_73), .O(gate415inter4));
  nand2 gate1056(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1057(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1058(.a(G29), .O(gate415inter7));
  inv1  gate1059(.a(G1120), .O(gate415inter8));
  nand2 gate1060(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1061(.a(s_73), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1062(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1063(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1064(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1079(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1080(.a(gate419inter0), .b(s_76), .O(gate419inter1));
  and2  gate1081(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1082(.a(s_76), .O(gate419inter3));
  inv1  gate1083(.a(s_77), .O(gate419inter4));
  nand2 gate1084(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1085(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1086(.a(G1), .O(gate419inter7));
  inv1  gate1087(.a(G1132), .O(gate419inter8));
  nand2 gate1088(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1089(.a(s_77), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1090(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1091(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1092(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate589(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate590(.a(gate422inter0), .b(s_6), .O(gate422inter1));
  and2  gate591(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate592(.a(s_6), .O(gate422inter3));
  inv1  gate593(.a(s_7), .O(gate422inter4));
  nand2 gate594(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate595(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate596(.a(G1039), .O(gate422inter7));
  inv1  gate597(.a(G1135), .O(gate422inter8));
  nand2 gate598(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate599(.a(s_7), .b(gate422inter3), .O(gate422inter10));
  nor2  gate600(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate601(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate602(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate981(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate982(.a(gate433inter0), .b(s_62), .O(gate433inter1));
  and2  gate983(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate984(.a(s_62), .O(gate433inter3));
  inv1  gate985(.a(s_63), .O(gate433inter4));
  nand2 gate986(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate987(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate988(.a(G8), .O(gate433inter7));
  inv1  gate989(.a(G1153), .O(gate433inter8));
  nand2 gate990(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate991(.a(s_63), .b(gate433inter3), .O(gate433inter10));
  nor2  gate992(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate993(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate994(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1065(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1066(.a(gate438inter0), .b(s_74), .O(gate438inter1));
  and2  gate1067(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1068(.a(s_74), .O(gate438inter3));
  inv1  gate1069(.a(s_75), .O(gate438inter4));
  nand2 gate1070(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1071(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1072(.a(G1063), .O(gate438inter7));
  inv1  gate1073(.a(G1159), .O(gate438inter8));
  nand2 gate1074(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1075(.a(s_75), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1076(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1077(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1078(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1093(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1094(.a(gate446inter0), .b(s_78), .O(gate446inter1));
  and2  gate1095(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1096(.a(s_78), .O(gate446inter3));
  inv1  gate1097(.a(s_79), .O(gate446inter4));
  nand2 gate1098(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1099(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1100(.a(G1075), .O(gate446inter7));
  inv1  gate1101(.a(G1171), .O(gate446inter8));
  nand2 gate1102(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1103(.a(s_79), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1104(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1105(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1106(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate771(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate772(.a(gate459inter0), .b(s_32), .O(gate459inter1));
  and2  gate773(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate774(.a(s_32), .O(gate459inter3));
  inv1  gate775(.a(s_33), .O(gate459inter4));
  nand2 gate776(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate777(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate778(.a(G21), .O(gate459inter7));
  inv1  gate779(.a(G1192), .O(gate459inter8));
  nand2 gate780(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate781(.a(s_33), .b(gate459inter3), .O(gate459inter10));
  nor2  gate782(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate783(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate784(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate967(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate968(.a(gate464inter0), .b(s_60), .O(gate464inter1));
  and2  gate969(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate970(.a(s_60), .O(gate464inter3));
  inv1  gate971(.a(s_61), .O(gate464inter4));
  nand2 gate972(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate973(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate974(.a(G1102), .O(gate464inter7));
  inv1  gate975(.a(G1198), .O(gate464inter8));
  nand2 gate976(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate977(.a(s_61), .b(gate464inter3), .O(gate464inter10));
  nor2  gate978(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate979(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate980(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1303(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1304(.a(gate469inter0), .b(s_108), .O(gate469inter1));
  and2  gate1305(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1306(.a(s_108), .O(gate469inter3));
  inv1  gate1307(.a(s_109), .O(gate469inter4));
  nand2 gate1308(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1309(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1310(.a(G26), .O(gate469inter7));
  inv1  gate1311(.a(G1207), .O(gate469inter8));
  nand2 gate1312(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1313(.a(s_109), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1314(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1315(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1316(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1275(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1276(.a(gate477inter0), .b(s_104), .O(gate477inter1));
  and2  gate1277(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1278(.a(s_104), .O(gate477inter3));
  inv1  gate1279(.a(s_105), .O(gate477inter4));
  nand2 gate1280(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1281(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1282(.a(G30), .O(gate477inter7));
  inv1  gate1283(.a(G1219), .O(gate477inter8));
  nand2 gate1284(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1285(.a(s_105), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1286(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1287(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1288(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate575(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate576(.a(gate480inter0), .b(s_4), .O(gate480inter1));
  and2  gate577(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate578(.a(s_4), .O(gate480inter3));
  inv1  gate579(.a(s_5), .O(gate480inter4));
  nand2 gate580(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate581(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate582(.a(G1126), .O(gate480inter7));
  inv1  gate583(.a(G1222), .O(gate480inter8));
  nand2 gate584(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate585(.a(s_5), .b(gate480inter3), .O(gate480inter10));
  nor2  gate586(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate587(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate588(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate547(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate548(.a(gate487inter0), .b(s_0), .O(gate487inter1));
  and2  gate549(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate550(.a(s_0), .O(gate487inter3));
  inv1  gate551(.a(s_1), .O(gate487inter4));
  nand2 gate552(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate553(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate554(.a(G1236), .O(gate487inter7));
  inv1  gate555(.a(G1237), .O(gate487inter8));
  nand2 gate556(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate557(.a(s_1), .b(gate487inter3), .O(gate487inter10));
  nor2  gate558(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate559(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate560(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate869(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate870(.a(gate494inter0), .b(s_46), .O(gate494inter1));
  and2  gate871(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate872(.a(s_46), .O(gate494inter3));
  inv1  gate873(.a(s_47), .O(gate494inter4));
  nand2 gate874(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate875(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate876(.a(G1250), .O(gate494inter7));
  inv1  gate877(.a(G1251), .O(gate494inter8));
  nand2 gate878(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate879(.a(s_47), .b(gate494inter3), .O(gate494inter10));
  nor2  gate880(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate881(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate882(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1191(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1192(.a(gate495inter0), .b(s_92), .O(gate495inter1));
  and2  gate1193(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1194(.a(s_92), .O(gate495inter3));
  inv1  gate1195(.a(s_93), .O(gate495inter4));
  nand2 gate1196(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1197(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1198(.a(G1252), .O(gate495inter7));
  inv1  gate1199(.a(G1253), .O(gate495inter8));
  nand2 gate1200(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1201(.a(s_93), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1202(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1203(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1204(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1009(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1010(.a(gate505inter0), .b(s_66), .O(gate505inter1));
  and2  gate1011(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1012(.a(s_66), .O(gate505inter3));
  inv1  gate1013(.a(s_67), .O(gate505inter4));
  nand2 gate1014(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1015(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1016(.a(G1272), .O(gate505inter7));
  inv1  gate1017(.a(G1273), .O(gate505inter8));
  nand2 gate1018(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1019(.a(s_67), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1020(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1021(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1022(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate911(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate912(.a(gate513inter0), .b(s_52), .O(gate513inter1));
  and2  gate913(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate914(.a(s_52), .O(gate513inter3));
  inv1  gate915(.a(s_53), .O(gate513inter4));
  nand2 gate916(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate917(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate918(.a(G1288), .O(gate513inter7));
  inv1  gate919(.a(G1289), .O(gate513inter8));
  nand2 gate920(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate921(.a(s_53), .b(gate513inter3), .O(gate513inter10));
  nor2  gate922(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate923(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate924(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule