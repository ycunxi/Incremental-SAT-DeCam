module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2479(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2480(.a(gate9inter0), .b(s_276), .O(gate9inter1));
  and2  gate2481(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2482(.a(s_276), .O(gate9inter3));
  inv1  gate2483(.a(s_277), .O(gate9inter4));
  nand2 gate2484(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2485(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2486(.a(G1), .O(gate9inter7));
  inv1  gate2487(.a(G2), .O(gate9inter8));
  nand2 gate2488(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2489(.a(s_277), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2490(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2491(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2492(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1205(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1206(.a(gate10inter0), .b(s_94), .O(gate10inter1));
  and2  gate1207(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1208(.a(s_94), .O(gate10inter3));
  inv1  gate1209(.a(s_95), .O(gate10inter4));
  nand2 gate1210(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1211(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1212(.a(G3), .O(gate10inter7));
  inv1  gate1213(.a(G4), .O(gate10inter8));
  nand2 gate1214(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1215(.a(s_95), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1216(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1217(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1218(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2143(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2144(.a(gate12inter0), .b(s_228), .O(gate12inter1));
  and2  gate2145(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2146(.a(s_228), .O(gate12inter3));
  inv1  gate2147(.a(s_229), .O(gate12inter4));
  nand2 gate2148(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2149(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2150(.a(G7), .O(gate12inter7));
  inv1  gate2151(.a(G8), .O(gate12inter8));
  nand2 gate2152(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2153(.a(s_229), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2154(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2155(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2156(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1163(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1164(.a(gate15inter0), .b(s_88), .O(gate15inter1));
  and2  gate1165(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1166(.a(s_88), .O(gate15inter3));
  inv1  gate1167(.a(s_89), .O(gate15inter4));
  nand2 gate1168(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1169(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1170(.a(G13), .O(gate15inter7));
  inv1  gate1171(.a(G14), .O(gate15inter8));
  nand2 gate1172(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1173(.a(s_89), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1174(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1175(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1176(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2381(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2382(.a(gate18inter0), .b(s_262), .O(gate18inter1));
  and2  gate2383(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2384(.a(s_262), .O(gate18inter3));
  inv1  gate2385(.a(s_263), .O(gate18inter4));
  nand2 gate2386(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2387(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2388(.a(G19), .O(gate18inter7));
  inv1  gate2389(.a(G20), .O(gate18inter8));
  nand2 gate2390(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2391(.a(s_263), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2392(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2393(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2394(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1905(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1906(.a(gate19inter0), .b(s_194), .O(gate19inter1));
  and2  gate1907(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1908(.a(s_194), .O(gate19inter3));
  inv1  gate1909(.a(s_195), .O(gate19inter4));
  nand2 gate1910(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1911(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1912(.a(G21), .O(gate19inter7));
  inv1  gate1913(.a(G22), .O(gate19inter8));
  nand2 gate1914(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1915(.a(s_195), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1916(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1917(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1918(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2367(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2368(.a(gate20inter0), .b(s_260), .O(gate20inter1));
  and2  gate2369(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2370(.a(s_260), .O(gate20inter3));
  inv1  gate2371(.a(s_261), .O(gate20inter4));
  nand2 gate2372(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2373(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2374(.a(G23), .O(gate20inter7));
  inv1  gate2375(.a(G24), .O(gate20inter8));
  nand2 gate2376(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2377(.a(s_261), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2378(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2379(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2380(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1821(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1822(.a(gate21inter0), .b(s_182), .O(gate21inter1));
  and2  gate1823(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1824(.a(s_182), .O(gate21inter3));
  inv1  gate1825(.a(s_183), .O(gate21inter4));
  nand2 gate1826(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1827(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1828(.a(G25), .O(gate21inter7));
  inv1  gate1829(.a(G26), .O(gate21inter8));
  nand2 gate1830(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1831(.a(s_183), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1832(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1833(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1834(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1121(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1122(.a(gate22inter0), .b(s_82), .O(gate22inter1));
  and2  gate1123(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1124(.a(s_82), .O(gate22inter3));
  inv1  gate1125(.a(s_83), .O(gate22inter4));
  nand2 gate1126(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1127(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1128(.a(G27), .O(gate22inter7));
  inv1  gate1129(.a(G28), .O(gate22inter8));
  nand2 gate1130(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1131(.a(s_83), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1132(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1133(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1134(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1807(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1808(.a(gate23inter0), .b(s_180), .O(gate23inter1));
  and2  gate1809(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1810(.a(s_180), .O(gate23inter3));
  inv1  gate1811(.a(s_181), .O(gate23inter4));
  nand2 gate1812(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1813(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1814(.a(G29), .O(gate23inter7));
  inv1  gate1815(.a(G30), .O(gate23inter8));
  nand2 gate1816(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1817(.a(s_181), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1818(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1819(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1820(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2857(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2858(.a(gate28inter0), .b(s_330), .O(gate28inter1));
  and2  gate2859(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2860(.a(s_330), .O(gate28inter3));
  inv1  gate2861(.a(s_331), .O(gate28inter4));
  nand2 gate2862(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2863(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2864(.a(G10), .O(gate28inter7));
  inv1  gate2865(.a(G14), .O(gate28inter8));
  nand2 gate2866(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2867(.a(s_331), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2868(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2869(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2870(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2703(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2704(.a(gate31inter0), .b(s_308), .O(gate31inter1));
  and2  gate2705(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2706(.a(s_308), .O(gate31inter3));
  inv1  gate2707(.a(s_309), .O(gate31inter4));
  nand2 gate2708(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2709(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2710(.a(G4), .O(gate31inter7));
  inv1  gate2711(.a(G8), .O(gate31inter8));
  nand2 gate2712(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2713(.a(s_309), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2714(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2715(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2716(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1107(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1108(.a(gate32inter0), .b(s_80), .O(gate32inter1));
  and2  gate1109(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1110(.a(s_80), .O(gate32inter3));
  inv1  gate1111(.a(s_81), .O(gate32inter4));
  nand2 gate1112(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1113(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1114(.a(G12), .O(gate32inter7));
  inv1  gate1115(.a(G16), .O(gate32inter8));
  nand2 gate1116(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1117(.a(s_81), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1118(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1119(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1120(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1135(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1136(.a(gate33inter0), .b(s_84), .O(gate33inter1));
  and2  gate1137(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1138(.a(s_84), .O(gate33inter3));
  inv1  gate1139(.a(s_85), .O(gate33inter4));
  nand2 gate1140(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1141(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1142(.a(G17), .O(gate33inter7));
  inv1  gate1143(.a(G21), .O(gate33inter8));
  nand2 gate1144(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1145(.a(s_85), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1146(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1147(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1148(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate547(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate548(.a(gate34inter0), .b(s_0), .O(gate34inter1));
  and2  gate549(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate550(.a(s_0), .O(gate34inter3));
  inv1  gate551(.a(s_1), .O(gate34inter4));
  nand2 gate552(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate553(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate554(.a(G25), .O(gate34inter7));
  inv1  gate555(.a(G29), .O(gate34inter8));
  nand2 gate556(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate557(.a(s_1), .b(gate34inter3), .O(gate34inter10));
  nor2  gate558(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate559(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate560(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1989(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1990(.a(gate35inter0), .b(s_206), .O(gate35inter1));
  and2  gate1991(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1992(.a(s_206), .O(gate35inter3));
  inv1  gate1993(.a(s_207), .O(gate35inter4));
  nand2 gate1994(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1995(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1996(.a(G18), .O(gate35inter7));
  inv1  gate1997(.a(G22), .O(gate35inter8));
  nand2 gate1998(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1999(.a(s_207), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2000(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2001(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2002(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1933(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1934(.a(gate43inter0), .b(s_198), .O(gate43inter1));
  and2  gate1935(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1936(.a(s_198), .O(gate43inter3));
  inv1  gate1937(.a(s_199), .O(gate43inter4));
  nand2 gate1938(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1939(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1940(.a(G3), .O(gate43inter7));
  inv1  gate1941(.a(G269), .O(gate43inter8));
  nand2 gate1942(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1943(.a(s_199), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1944(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1945(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1946(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2451(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2452(.a(gate44inter0), .b(s_272), .O(gate44inter1));
  and2  gate2453(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2454(.a(s_272), .O(gate44inter3));
  inv1  gate2455(.a(s_273), .O(gate44inter4));
  nand2 gate2456(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2457(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2458(.a(G4), .O(gate44inter7));
  inv1  gate2459(.a(G269), .O(gate44inter8));
  nand2 gate2460(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2461(.a(s_273), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2462(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2463(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2464(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate939(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate940(.a(gate46inter0), .b(s_56), .O(gate46inter1));
  and2  gate941(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate942(.a(s_56), .O(gate46inter3));
  inv1  gate943(.a(s_57), .O(gate46inter4));
  nand2 gate944(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate945(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate946(.a(G6), .O(gate46inter7));
  inv1  gate947(.a(G272), .O(gate46inter8));
  nand2 gate948(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate949(.a(s_57), .b(gate46inter3), .O(gate46inter10));
  nor2  gate950(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate951(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate952(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2843(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2844(.a(gate48inter0), .b(s_328), .O(gate48inter1));
  and2  gate2845(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2846(.a(s_328), .O(gate48inter3));
  inv1  gate2847(.a(s_329), .O(gate48inter4));
  nand2 gate2848(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2849(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2850(.a(G8), .O(gate48inter7));
  inv1  gate2851(.a(G275), .O(gate48inter8));
  nand2 gate2852(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2853(.a(s_329), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2854(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2855(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2856(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate715(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate716(.a(gate49inter0), .b(s_24), .O(gate49inter1));
  and2  gate717(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate718(.a(s_24), .O(gate49inter3));
  inv1  gate719(.a(s_25), .O(gate49inter4));
  nand2 gate720(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate721(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate722(.a(G9), .O(gate49inter7));
  inv1  gate723(.a(G278), .O(gate49inter8));
  nand2 gate724(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate725(.a(s_25), .b(gate49inter3), .O(gate49inter10));
  nor2  gate726(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate727(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate728(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1443(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1444(.a(gate57inter0), .b(s_128), .O(gate57inter1));
  and2  gate1445(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1446(.a(s_128), .O(gate57inter3));
  inv1  gate1447(.a(s_129), .O(gate57inter4));
  nand2 gate1448(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1449(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1450(.a(G17), .O(gate57inter7));
  inv1  gate1451(.a(G290), .O(gate57inter8));
  nand2 gate1452(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1453(.a(s_129), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1454(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1455(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1456(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2185(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2186(.a(gate59inter0), .b(s_234), .O(gate59inter1));
  and2  gate2187(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2188(.a(s_234), .O(gate59inter3));
  inv1  gate2189(.a(s_235), .O(gate59inter4));
  nand2 gate2190(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2191(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2192(.a(G19), .O(gate59inter7));
  inv1  gate2193(.a(G293), .O(gate59inter8));
  nand2 gate2194(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2195(.a(s_235), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2196(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2197(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2198(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate603(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate604(.a(gate60inter0), .b(s_8), .O(gate60inter1));
  and2  gate605(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate606(.a(s_8), .O(gate60inter3));
  inv1  gate607(.a(s_9), .O(gate60inter4));
  nand2 gate608(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate609(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate610(.a(G20), .O(gate60inter7));
  inv1  gate611(.a(G293), .O(gate60inter8));
  nand2 gate612(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate613(.a(s_9), .b(gate60inter3), .O(gate60inter10));
  nor2  gate614(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate615(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate616(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1359(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1360(.a(gate62inter0), .b(s_116), .O(gate62inter1));
  and2  gate1361(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1362(.a(s_116), .O(gate62inter3));
  inv1  gate1363(.a(s_117), .O(gate62inter4));
  nand2 gate1364(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1365(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1366(.a(G22), .O(gate62inter7));
  inv1  gate1367(.a(G296), .O(gate62inter8));
  nand2 gate1368(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1369(.a(s_117), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1370(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1371(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1372(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate855(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate856(.a(gate63inter0), .b(s_44), .O(gate63inter1));
  and2  gate857(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate858(.a(s_44), .O(gate63inter3));
  inv1  gate859(.a(s_45), .O(gate63inter4));
  nand2 gate860(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate861(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate862(.a(G23), .O(gate63inter7));
  inv1  gate863(.a(G299), .O(gate63inter8));
  nand2 gate864(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate865(.a(s_45), .b(gate63inter3), .O(gate63inter10));
  nor2  gate866(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate867(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate868(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2717(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2718(.a(gate66inter0), .b(s_310), .O(gate66inter1));
  and2  gate2719(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2720(.a(s_310), .O(gate66inter3));
  inv1  gate2721(.a(s_311), .O(gate66inter4));
  nand2 gate2722(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2723(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2724(.a(G26), .O(gate66inter7));
  inv1  gate2725(.a(G302), .O(gate66inter8));
  nand2 gate2726(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2727(.a(s_311), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2728(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2729(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2730(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1891(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1892(.a(gate67inter0), .b(s_192), .O(gate67inter1));
  and2  gate1893(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1894(.a(s_192), .O(gate67inter3));
  inv1  gate1895(.a(s_193), .O(gate67inter4));
  nand2 gate1896(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1897(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1898(.a(G27), .O(gate67inter7));
  inv1  gate1899(.a(G305), .O(gate67inter8));
  nand2 gate1900(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1901(.a(s_193), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1902(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1903(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1904(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate2675(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2676(.a(gate68inter0), .b(s_304), .O(gate68inter1));
  and2  gate2677(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2678(.a(s_304), .O(gate68inter3));
  inv1  gate2679(.a(s_305), .O(gate68inter4));
  nand2 gate2680(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2681(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2682(.a(G28), .O(gate68inter7));
  inv1  gate2683(.a(G305), .O(gate68inter8));
  nand2 gate2684(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2685(.a(s_305), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2686(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2687(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2688(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate1499(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1500(.a(gate69inter0), .b(s_136), .O(gate69inter1));
  and2  gate1501(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1502(.a(s_136), .O(gate69inter3));
  inv1  gate1503(.a(s_137), .O(gate69inter4));
  nand2 gate1504(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1505(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1506(.a(G29), .O(gate69inter7));
  inv1  gate1507(.a(G308), .O(gate69inter8));
  nand2 gate1508(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1509(.a(s_137), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1510(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1511(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1512(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate673(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate674(.a(gate76inter0), .b(s_18), .O(gate76inter1));
  and2  gate675(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate676(.a(s_18), .O(gate76inter3));
  inv1  gate677(.a(s_19), .O(gate76inter4));
  nand2 gate678(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate679(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate680(.a(G13), .O(gate76inter7));
  inv1  gate681(.a(G317), .O(gate76inter8));
  nand2 gate682(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate683(.a(s_19), .b(gate76inter3), .O(gate76inter10));
  nor2  gate684(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate685(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate686(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate757(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate758(.a(gate77inter0), .b(s_30), .O(gate77inter1));
  and2  gate759(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate760(.a(s_30), .O(gate77inter3));
  inv1  gate761(.a(s_31), .O(gate77inter4));
  nand2 gate762(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate763(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate764(.a(G2), .O(gate77inter7));
  inv1  gate765(.a(G320), .O(gate77inter8));
  nand2 gate766(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate767(.a(s_31), .b(gate77inter3), .O(gate77inter10));
  nor2  gate768(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate769(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate770(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2311(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2312(.a(gate80inter0), .b(s_252), .O(gate80inter1));
  and2  gate2313(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2314(.a(s_252), .O(gate80inter3));
  inv1  gate2315(.a(s_253), .O(gate80inter4));
  nand2 gate2316(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2317(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2318(.a(G14), .O(gate80inter7));
  inv1  gate2319(.a(G323), .O(gate80inter8));
  nand2 gate2320(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2321(.a(s_253), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2322(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2323(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2324(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate911(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate912(.a(gate81inter0), .b(s_52), .O(gate81inter1));
  and2  gate913(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate914(.a(s_52), .O(gate81inter3));
  inv1  gate915(.a(s_53), .O(gate81inter4));
  nand2 gate916(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate917(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate918(.a(G3), .O(gate81inter7));
  inv1  gate919(.a(G326), .O(gate81inter8));
  nand2 gate920(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate921(.a(s_53), .b(gate81inter3), .O(gate81inter10));
  nor2  gate922(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate923(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate924(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1429(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1430(.a(gate87inter0), .b(s_126), .O(gate87inter1));
  and2  gate1431(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1432(.a(s_126), .O(gate87inter3));
  inv1  gate1433(.a(s_127), .O(gate87inter4));
  nand2 gate1434(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1435(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1436(.a(G12), .O(gate87inter7));
  inv1  gate1437(.a(G335), .O(gate87inter8));
  nand2 gate1438(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1439(.a(s_127), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1440(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1441(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1442(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate897(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate898(.a(gate88inter0), .b(s_50), .O(gate88inter1));
  and2  gate899(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate900(.a(s_50), .O(gate88inter3));
  inv1  gate901(.a(s_51), .O(gate88inter4));
  nand2 gate902(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate903(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate904(.a(G16), .O(gate88inter7));
  inv1  gate905(.a(G335), .O(gate88inter8));
  nand2 gate906(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate907(.a(s_51), .b(gate88inter3), .O(gate88inter10));
  nor2  gate908(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate909(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate910(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2577(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2578(.a(gate92inter0), .b(s_290), .O(gate92inter1));
  and2  gate2579(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2580(.a(s_290), .O(gate92inter3));
  inv1  gate2581(.a(s_291), .O(gate92inter4));
  nand2 gate2582(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2583(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2584(.a(G29), .O(gate92inter7));
  inv1  gate2585(.a(G341), .O(gate92inter8));
  nand2 gate2586(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2587(.a(s_291), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2588(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2589(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2590(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1555(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1556(.a(gate93inter0), .b(s_144), .O(gate93inter1));
  and2  gate1557(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1558(.a(s_144), .O(gate93inter3));
  inv1  gate1559(.a(s_145), .O(gate93inter4));
  nand2 gate1560(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1561(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1562(.a(G18), .O(gate93inter7));
  inv1  gate1563(.a(G344), .O(gate93inter8));
  nand2 gate1564(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1565(.a(s_145), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1566(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1567(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1568(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate883(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate884(.a(gate98inter0), .b(s_48), .O(gate98inter1));
  and2  gate885(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate886(.a(s_48), .O(gate98inter3));
  inv1  gate887(.a(s_49), .O(gate98inter4));
  nand2 gate888(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate889(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate890(.a(G23), .O(gate98inter7));
  inv1  gate891(.a(G350), .O(gate98inter8));
  nand2 gate892(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate893(.a(s_49), .b(gate98inter3), .O(gate98inter10));
  nor2  gate894(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate895(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate896(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1387(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1388(.a(gate99inter0), .b(s_120), .O(gate99inter1));
  and2  gate1389(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1390(.a(s_120), .O(gate99inter3));
  inv1  gate1391(.a(s_121), .O(gate99inter4));
  nand2 gate1392(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1393(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1394(.a(G27), .O(gate99inter7));
  inv1  gate1395(.a(G353), .O(gate99inter8));
  nand2 gate1396(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1397(.a(s_121), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1398(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1399(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1400(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1401(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1402(.a(gate101inter0), .b(s_122), .O(gate101inter1));
  and2  gate1403(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1404(.a(s_122), .O(gate101inter3));
  inv1  gate1405(.a(s_123), .O(gate101inter4));
  nand2 gate1406(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1407(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1408(.a(G20), .O(gate101inter7));
  inv1  gate1409(.a(G356), .O(gate101inter8));
  nand2 gate1410(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1411(.a(s_123), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1412(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1413(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1414(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2353(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2354(.a(gate105inter0), .b(s_258), .O(gate105inter1));
  and2  gate2355(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2356(.a(s_258), .O(gate105inter3));
  inv1  gate2357(.a(s_259), .O(gate105inter4));
  nand2 gate2358(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2359(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2360(.a(G362), .O(gate105inter7));
  inv1  gate2361(.a(G363), .O(gate105inter8));
  nand2 gate2362(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2363(.a(s_259), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2364(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2365(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2366(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate631(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate632(.a(gate109inter0), .b(s_12), .O(gate109inter1));
  and2  gate633(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate634(.a(s_12), .O(gate109inter3));
  inv1  gate635(.a(s_13), .O(gate109inter4));
  nand2 gate636(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate637(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate638(.a(G370), .O(gate109inter7));
  inv1  gate639(.a(G371), .O(gate109inter8));
  nand2 gate640(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate641(.a(s_13), .b(gate109inter3), .O(gate109inter10));
  nor2  gate642(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate643(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate644(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1527(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1528(.a(gate110inter0), .b(s_140), .O(gate110inter1));
  and2  gate1529(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1530(.a(s_140), .O(gate110inter3));
  inv1  gate1531(.a(s_141), .O(gate110inter4));
  nand2 gate1532(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1533(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1534(.a(G372), .O(gate110inter7));
  inv1  gate1535(.a(G373), .O(gate110inter8));
  nand2 gate1536(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1537(.a(s_141), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1538(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1539(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1540(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1569(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1570(.a(gate113inter0), .b(s_146), .O(gate113inter1));
  and2  gate1571(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1572(.a(s_146), .O(gate113inter3));
  inv1  gate1573(.a(s_147), .O(gate113inter4));
  nand2 gate1574(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1575(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1576(.a(G378), .O(gate113inter7));
  inv1  gate1577(.a(G379), .O(gate113inter8));
  nand2 gate1578(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1579(.a(s_147), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1580(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1581(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1582(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1233(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1234(.a(gate115inter0), .b(s_98), .O(gate115inter1));
  and2  gate1235(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1236(.a(s_98), .O(gate115inter3));
  inv1  gate1237(.a(s_99), .O(gate115inter4));
  nand2 gate1238(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1239(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1240(.a(G382), .O(gate115inter7));
  inv1  gate1241(.a(G383), .O(gate115inter8));
  nand2 gate1242(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1243(.a(s_99), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1244(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1245(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1246(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1723(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1724(.a(gate116inter0), .b(s_168), .O(gate116inter1));
  and2  gate1725(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1726(.a(s_168), .O(gate116inter3));
  inv1  gate1727(.a(s_169), .O(gate116inter4));
  nand2 gate1728(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1729(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1730(.a(G384), .O(gate116inter7));
  inv1  gate1731(.a(G385), .O(gate116inter8));
  nand2 gate1732(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1733(.a(s_169), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1734(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1735(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1736(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1541(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1542(.a(gate118inter0), .b(s_142), .O(gate118inter1));
  and2  gate1543(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1544(.a(s_142), .O(gate118inter3));
  inv1  gate1545(.a(s_143), .O(gate118inter4));
  nand2 gate1546(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1547(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1548(.a(G388), .O(gate118inter7));
  inv1  gate1549(.a(G389), .O(gate118inter8));
  nand2 gate1550(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1551(.a(s_143), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1552(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1553(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1554(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2801(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2802(.a(gate119inter0), .b(s_322), .O(gate119inter1));
  and2  gate2803(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2804(.a(s_322), .O(gate119inter3));
  inv1  gate2805(.a(s_323), .O(gate119inter4));
  nand2 gate2806(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2807(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2808(.a(G390), .O(gate119inter7));
  inv1  gate2809(.a(G391), .O(gate119inter8));
  nand2 gate2810(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2811(.a(s_323), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2812(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2813(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2814(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate645(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate646(.a(gate123inter0), .b(s_14), .O(gate123inter1));
  and2  gate647(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate648(.a(s_14), .O(gate123inter3));
  inv1  gate649(.a(s_15), .O(gate123inter4));
  nand2 gate650(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate651(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate652(.a(G398), .O(gate123inter7));
  inv1  gate653(.a(G399), .O(gate123inter8));
  nand2 gate654(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate655(.a(s_15), .b(gate123inter3), .O(gate123inter10));
  nor2  gate656(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate657(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate658(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2829(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2830(.a(gate125inter0), .b(s_326), .O(gate125inter1));
  and2  gate2831(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2832(.a(s_326), .O(gate125inter3));
  inv1  gate2833(.a(s_327), .O(gate125inter4));
  nand2 gate2834(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2835(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2836(.a(G402), .O(gate125inter7));
  inv1  gate2837(.a(G403), .O(gate125inter8));
  nand2 gate2838(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2839(.a(s_327), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2840(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2841(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2842(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1303(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1304(.a(gate130inter0), .b(s_108), .O(gate130inter1));
  and2  gate1305(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1306(.a(s_108), .O(gate130inter3));
  inv1  gate1307(.a(s_109), .O(gate130inter4));
  nand2 gate1308(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1309(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1310(.a(G412), .O(gate130inter7));
  inv1  gate1311(.a(G413), .O(gate130inter8));
  nand2 gate1312(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1313(.a(s_109), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1314(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1315(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1316(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2507(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2508(.a(gate131inter0), .b(s_280), .O(gate131inter1));
  and2  gate2509(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2510(.a(s_280), .O(gate131inter3));
  inv1  gate2511(.a(s_281), .O(gate131inter4));
  nand2 gate2512(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2513(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2514(.a(G414), .O(gate131inter7));
  inv1  gate2515(.a(G415), .O(gate131inter8));
  nand2 gate2516(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2517(.a(s_281), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2518(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2519(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2520(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate2731(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2732(.a(gate132inter0), .b(s_312), .O(gate132inter1));
  and2  gate2733(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2734(.a(s_312), .O(gate132inter3));
  inv1  gate2735(.a(s_313), .O(gate132inter4));
  nand2 gate2736(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2737(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2738(.a(G416), .O(gate132inter7));
  inv1  gate2739(.a(G417), .O(gate132inter8));
  nand2 gate2740(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2741(.a(s_313), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2742(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2743(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2744(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2325(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2326(.a(gate136inter0), .b(s_254), .O(gate136inter1));
  and2  gate2327(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2328(.a(s_254), .O(gate136inter3));
  inv1  gate2329(.a(s_255), .O(gate136inter4));
  nand2 gate2330(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2331(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2332(.a(G424), .O(gate136inter7));
  inv1  gate2333(.a(G425), .O(gate136inter8));
  nand2 gate2334(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2335(.a(s_255), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2336(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2337(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2338(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1653(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1654(.a(gate137inter0), .b(s_158), .O(gate137inter1));
  and2  gate1655(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1656(.a(s_158), .O(gate137inter3));
  inv1  gate1657(.a(s_159), .O(gate137inter4));
  nand2 gate1658(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1659(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1660(.a(G426), .O(gate137inter7));
  inv1  gate1661(.a(G429), .O(gate137inter8));
  nand2 gate1662(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1663(.a(s_159), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1664(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1665(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1666(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1373(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1374(.a(gate138inter0), .b(s_118), .O(gate138inter1));
  and2  gate1375(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1376(.a(s_118), .O(gate138inter3));
  inv1  gate1377(.a(s_119), .O(gate138inter4));
  nand2 gate1378(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1379(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1380(.a(G432), .O(gate138inter7));
  inv1  gate1381(.a(G435), .O(gate138inter8));
  nand2 gate1382(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1383(.a(s_119), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1384(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1385(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1386(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2563(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2564(.a(gate139inter0), .b(s_288), .O(gate139inter1));
  and2  gate2565(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2566(.a(s_288), .O(gate139inter3));
  inv1  gate2567(.a(s_289), .O(gate139inter4));
  nand2 gate2568(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2569(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2570(.a(G438), .O(gate139inter7));
  inv1  gate2571(.a(G441), .O(gate139inter8));
  nand2 gate2572(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2573(.a(s_289), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2574(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2575(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2576(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2815(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2816(.a(gate140inter0), .b(s_324), .O(gate140inter1));
  and2  gate2817(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2818(.a(s_324), .O(gate140inter3));
  inv1  gate2819(.a(s_325), .O(gate140inter4));
  nand2 gate2820(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2821(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2822(.a(G444), .O(gate140inter7));
  inv1  gate2823(.a(G447), .O(gate140inter8));
  nand2 gate2824(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2825(.a(s_325), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2826(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2827(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2828(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate2003(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2004(.a(gate141inter0), .b(s_208), .O(gate141inter1));
  and2  gate2005(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2006(.a(s_208), .O(gate141inter3));
  inv1  gate2007(.a(s_209), .O(gate141inter4));
  nand2 gate2008(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2009(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2010(.a(G450), .O(gate141inter7));
  inv1  gate2011(.a(G453), .O(gate141inter8));
  nand2 gate2012(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2013(.a(s_209), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2014(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2015(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2016(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate617(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate618(.a(gate144inter0), .b(s_10), .O(gate144inter1));
  and2  gate619(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate620(.a(s_10), .O(gate144inter3));
  inv1  gate621(.a(s_11), .O(gate144inter4));
  nand2 gate622(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate623(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate624(.a(G468), .O(gate144inter7));
  inv1  gate625(.a(G471), .O(gate144inter8));
  nand2 gate626(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate627(.a(s_11), .b(gate144inter3), .O(gate144inter10));
  nor2  gate628(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate629(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate630(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate925(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate926(.a(gate147inter0), .b(s_54), .O(gate147inter1));
  and2  gate927(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate928(.a(s_54), .O(gate147inter3));
  inv1  gate929(.a(s_55), .O(gate147inter4));
  nand2 gate930(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate931(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate932(.a(G486), .O(gate147inter7));
  inv1  gate933(.a(G489), .O(gate147inter8));
  nand2 gate934(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate935(.a(s_55), .b(gate147inter3), .O(gate147inter10));
  nor2  gate936(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate937(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate938(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate2073(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2074(.a(gate148inter0), .b(s_218), .O(gate148inter1));
  and2  gate2075(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2076(.a(s_218), .O(gate148inter3));
  inv1  gate2077(.a(s_219), .O(gate148inter4));
  nand2 gate2078(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2079(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2080(.a(G492), .O(gate148inter7));
  inv1  gate2081(.a(G495), .O(gate148inter8));
  nand2 gate2082(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2083(.a(s_219), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2084(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2085(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2086(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2199(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2200(.a(gate150inter0), .b(s_236), .O(gate150inter1));
  and2  gate2201(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2202(.a(s_236), .O(gate150inter3));
  inv1  gate2203(.a(s_237), .O(gate150inter4));
  nand2 gate2204(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2205(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2206(.a(G504), .O(gate150inter7));
  inv1  gate2207(.a(G507), .O(gate150inter8));
  nand2 gate2208(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2209(.a(s_237), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2210(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2211(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2212(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1863(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1864(.a(gate152inter0), .b(s_188), .O(gate152inter1));
  and2  gate1865(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1866(.a(s_188), .O(gate152inter3));
  inv1  gate1867(.a(s_189), .O(gate152inter4));
  nand2 gate1868(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1869(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1870(.a(G516), .O(gate152inter7));
  inv1  gate1871(.a(G519), .O(gate152inter8));
  nand2 gate1872(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1873(.a(s_189), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1874(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1875(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1876(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate1037(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1038(.a(gate153inter0), .b(s_70), .O(gate153inter1));
  and2  gate1039(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1040(.a(s_70), .O(gate153inter3));
  inv1  gate1041(.a(s_71), .O(gate153inter4));
  nand2 gate1042(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1043(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1044(.a(G426), .O(gate153inter7));
  inv1  gate1045(.a(G522), .O(gate153inter8));
  nand2 gate1046(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1047(.a(s_71), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1048(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1049(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1050(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1779(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1780(.a(gate154inter0), .b(s_176), .O(gate154inter1));
  and2  gate1781(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1782(.a(s_176), .O(gate154inter3));
  inv1  gate1783(.a(s_177), .O(gate154inter4));
  nand2 gate1784(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1785(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1786(.a(G429), .O(gate154inter7));
  inv1  gate1787(.a(G522), .O(gate154inter8));
  nand2 gate1788(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1789(.a(s_177), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1790(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1791(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1792(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1681(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1682(.a(gate158inter0), .b(s_162), .O(gate158inter1));
  and2  gate1683(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1684(.a(s_162), .O(gate158inter3));
  inv1  gate1685(.a(s_163), .O(gate158inter4));
  nand2 gate1686(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1687(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1688(.a(G441), .O(gate158inter7));
  inv1  gate1689(.a(G528), .O(gate158inter8));
  nand2 gate1690(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1691(.a(s_163), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1692(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1693(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1694(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1611(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1612(.a(gate163inter0), .b(s_152), .O(gate163inter1));
  and2  gate1613(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1614(.a(s_152), .O(gate163inter3));
  inv1  gate1615(.a(s_153), .O(gate163inter4));
  nand2 gate1616(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1617(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1618(.a(G456), .O(gate163inter7));
  inv1  gate1619(.a(G537), .O(gate163inter8));
  nand2 gate1620(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1621(.a(s_153), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1622(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1623(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1624(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2661(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2662(.a(gate164inter0), .b(s_302), .O(gate164inter1));
  and2  gate2663(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2664(.a(s_302), .O(gate164inter3));
  inv1  gate2665(.a(s_303), .O(gate164inter4));
  nand2 gate2666(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2667(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2668(.a(G459), .O(gate164inter7));
  inv1  gate2669(.a(G537), .O(gate164inter8));
  nand2 gate2670(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2671(.a(s_303), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2672(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2673(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2674(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate659(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate660(.a(gate169inter0), .b(s_16), .O(gate169inter1));
  and2  gate661(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate662(.a(s_16), .O(gate169inter3));
  inv1  gate663(.a(s_17), .O(gate169inter4));
  nand2 gate664(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate665(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate666(.a(G474), .O(gate169inter7));
  inv1  gate667(.a(G546), .O(gate169inter8));
  nand2 gate668(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate669(.a(s_17), .b(gate169inter3), .O(gate169inter10));
  nor2  gate670(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate671(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate672(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2549(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2550(.a(gate171inter0), .b(s_286), .O(gate171inter1));
  and2  gate2551(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2552(.a(s_286), .O(gate171inter3));
  inv1  gate2553(.a(s_287), .O(gate171inter4));
  nand2 gate2554(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2555(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2556(.a(G480), .O(gate171inter7));
  inv1  gate2557(.a(G549), .O(gate171inter8));
  nand2 gate2558(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2559(.a(s_287), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2560(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2561(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2562(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2619(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2620(.a(gate176inter0), .b(s_296), .O(gate176inter1));
  and2  gate2621(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2622(.a(s_296), .O(gate176inter3));
  inv1  gate2623(.a(s_297), .O(gate176inter4));
  nand2 gate2624(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2625(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2626(.a(G495), .O(gate176inter7));
  inv1  gate2627(.a(G555), .O(gate176inter8));
  nand2 gate2628(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2629(.a(s_297), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2630(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2631(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2632(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2283(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2284(.a(gate184inter0), .b(s_248), .O(gate184inter1));
  and2  gate2285(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2286(.a(s_248), .O(gate184inter3));
  inv1  gate2287(.a(s_249), .O(gate184inter4));
  nand2 gate2288(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2289(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2290(.a(G519), .O(gate184inter7));
  inv1  gate2291(.a(G567), .O(gate184inter8));
  nand2 gate2292(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2293(.a(s_249), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2294(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2295(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2296(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate743(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate744(.a(gate185inter0), .b(s_28), .O(gate185inter1));
  and2  gate745(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate746(.a(s_28), .O(gate185inter3));
  inv1  gate747(.a(s_29), .O(gate185inter4));
  nand2 gate748(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate749(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate750(.a(G570), .O(gate185inter7));
  inv1  gate751(.a(G571), .O(gate185inter8));
  nand2 gate752(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate753(.a(s_29), .b(gate185inter3), .O(gate185inter10));
  nor2  gate754(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate755(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate756(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2591(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2592(.a(gate186inter0), .b(s_292), .O(gate186inter1));
  and2  gate2593(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2594(.a(s_292), .O(gate186inter3));
  inv1  gate2595(.a(s_293), .O(gate186inter4));
  nand2 gate2596(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2597(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2598(.a(G572), .O(gate186inter7));
  inv1  gate2599(.a(G573), .O(gate186inter8));
  nand2 gate2600(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2601(.a(s_293), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2602(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2603(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2604(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1751(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1752(.a(gate191inter0), .b(s_172), .O(gate191inter1));
  and2  gate1753(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1754(.a(s_172), .O(gate191inter3));
  inv1  gate1755(.a(s_173), .O(gate191inter4));
  nand2 gate1756(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1757(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1758(.a(G582), .O(gate191inter7));
  inv1  gate1759(.a(G583), .O(gate191inter8));
  nand2 gate1760(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1761(.a(s_173), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1762(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1763(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1764(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1317(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1318(.a(gate192inter0), .b(s_110), .O(gate192inter1));
  and2  gate1319(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1320(.a(s_110), .O(gate192inter3));
  inv1  gate1321(.a(s_111), .O(gate192inter4));
  nand2 gate1322(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1323(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1324(.a(G584), .O(gate192inter7));
  inv1  gate1325(.a(G585), .O(gate192inter8));
  nand2 gate1326(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1327(.a(s_111), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1328(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1329(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1330(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1709(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1710(.a(gate197inter0), .b(s_166), .O(gate197inter1));
  and2  gate1711(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1712(.a(s_166), .O(gate197inter3));
  inv1  gate1713(.a(s_167), .O(gate197inter4));
  nand2 gate1714(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1715(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1716(.a(G594), .O(gate197inter7));
  inv1  gate1717(.a(G595), .O(gate197inter8));
  nand2 gate1718(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1719(.a(s_167), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1720(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1721(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1722(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2213(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2214(.a(gate205inter0), .b(s_238), .O(gate205inter1));
  and2  gate2215(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2216(.a(s_238), .O(gate205inter3));
  inv1  gate2217(.a(s_239), .O(gate205inter4));
  nand2 gate2218(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2219(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2220(.a(G622), .O(gate205inter7));
  inv1  gate2221(.a(G627), .O(gate205inter8));
  nand2 gate2222(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2223(.a(s_239), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2224(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2225(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2226(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1597(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1598(.a(gate206inter0), .b(s_150), .O(gate206inter1));
  and2  gate1599(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1600(.a(s_150), .O(gate206inter3));
  inv1  gate1601(.a(s_151), .O(gate206inter4));
  nand2 gate1602(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1603(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1604(.a(G632), .O(gate206inter7));
  inv1  gate1605(.a(G637), .O(gate206inter8));
  nand2 gate1606(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1607(.a(s_151), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1608(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1609(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1610(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2521(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2522(.a(gate207inter0), .b(s_282), .O(gate207inter1));
  and2  gate2523(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2524(.a(s_282), .O(gate207inter3));
  inv1  gate2525(.a(s_283), .O(gate207inter4));
  nand2 gate2526(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2527(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2528(.a(G622), .O(gate207inter7));
  inv1  gate2529(.a(G632), .O(gate207inter8));
  nand2 gate2530(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2531(.a(s_283), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2532(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2533(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2534(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2017(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2018(.a(gate209inter0), .b(s_210), .O(gate209inter1));
  and2  gate2019(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2020(.a(s_210), .O(gate209inter3));
  inv1  gate2021(.a(s_211), .O(gate209inter4));
  nand2 gate2022(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2023(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2024(.a(G602), .O(gate209inter7));
  inv1  gate2025(.a(G666), .O(gate209inter8));
  nand2 gate2026(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2027(.a(s_211), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2028(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2029(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2030(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate729(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate730(.a(gate210inter0), .b(s_26), .O(gate210inter1));
  and2  gate731(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate732(.a(s_26), .O(gate210inter3));
  inv1  gate733(.a(s_27), .O(gate210inter4));
  nand2 gate734(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate735(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate736(.a(G607), .O(gate210inter7));
  inv1  gate737(.a(G666), .O(gate210inter8));
  nand2 gate738(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate739(.a(s_27), .b(gate210inter3), .O(gate210inter10));
  nor2  gate740(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate741(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate742(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1275(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1276(.a(gate213inter0), .b(s_104), .O(gate213inter1));
  and2  gate1277(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1278(.a(s_104), .O(gate213inter3));
  inv1  gate1279(.a(s_105), .O(gate213inter4));
  nand2 gate1280(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1281(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1282(.a(G602), .O(gate213inter7));
  inv1  gate1283(.a(G672), .O(gate213inter8));
  nand2 gate1284(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1285(.a(s_105), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1286(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1287(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1288(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1079(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1080(.a(gate214inter0), .b(s_76), .O(gate214inter1));
  and2  gate1081(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1082(.a(s_76), .O(gate214inter3));
  inv1  gate1083(.a(s_77), .O(gate214inter4));
  nand2 gate1084(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1085(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1086(.a(G612), .O(gate214inter7));
  inv1  gate1087(.a(G672), .O(gate214inter8));
  nand2 gate1088(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1089(.a(s_77), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1090(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1091(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1092(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate575(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate576(.a(gate216inter0), .b(s_4), .O(gate216inter1));
  and2  gate577(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate578(.a(s_4), .O(gate216inter3));
  inv1  gate579(.a(s_5), .O(gate216inter4));
  nand2 gate580(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate581(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate582(.a(G617), .O(gate216inter7));
  inv1  gate583(.a(G675), .O(gate216inter8));
  nand2 gate584(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate585(.a(s_5), .b(gate216inter3), .O(gate216inter10));
  nor2  gate586(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate587(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate588(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2927(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2928(.a(gate219inter0), .b(s_340), .O(gate219inter1));
  and2  gate2929(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2930(.a(s_340), .O(gate219inter3));
  inv1  gate2931(.a(s_341), .O(gate219inter4));
  nand2 gate2932(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2933(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2934(.a(G632), .O(gate219inter7));
  inv1  gate2935(.a(G681), .O(gate219inter8));
  nand2 gate2936(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2937(.a(s_341), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2938(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2939(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2940(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1877(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1878(.a(gate223inter0), .b(s_190), .O(gate223inter1));
  and2  gate1879(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1880(.a(s_190), .O(gate223inter3));
  inv1  gate1881(.a(s_191), .O(gate223inter4));
  nand2 gate1882(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1883(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1884(.a(G627), .O(gate223inter7));
  inv1  gate1885(.a(G687), .O(gate223inter8));
  nand2 gate1886(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1887(.a(s_191), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1888(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1889(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1890(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1457(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1458(.a(gate224inter0), .b(s_130), .O(gate224inter1));
  and2  gate1459(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1460(.a(s_130), .O(gate224inter3));
  inv1  gate1461(.a(s_131), .O(gate224inter4));
  nand2 gate1462(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1463(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1464(.a(G637), .O(gate224inter7));
  inv1  gate1465(.a(G687), .O(gate224inter8));
  nand2 gate1466(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1467(.a(s_131), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1468(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1469(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1470(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2787(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2788(.a(gate230inter0), .b(s_320), .O(gate230inter1));
  and2  gate2789(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2790(.a(s_320), .O(gate230inter3));
  inv1  gate2791(.a(s_321), .O(gate230inter4));
  nand2 gate2792(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2793(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2794(.a(G700), .O(gate230inter7));
  inv1  gate2795(.a(G701), .O(gate230inter8));
  nand2 gate2796(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2797(.a(s_321), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2798(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2799(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2800(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2255(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2256(.a(gate231inter0), .b(s_244), .O(gate231inter1));
  and2  gate2257(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2258(.a(s_244), .O(gate231inter3));
  inv1  gate2259(.a(s_245), .O(gate231inter4));
  nand2 gate2260(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2261(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2262(.a(G702), .O(gate231inter7));
  inv1  gate2263(.a(G703), .O(gate231inter8));
  nand2 gate2264(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2265(.a(s_245), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2266(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2267(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2268(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2129(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2130(.a(gate234inter0), .b(s_226), .O(gate234inter1));
  and2  gate2131(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2132(.a(s_226), .O(gate234inter3));
  inv1  gate2133(.a(s_227), .O(gate234inter4));
  nand2 gate2134(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2135(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2136(.a(G245), .O(gate234inter7));
  inv1  gate2137(.a(G721), .O(gate234inter8));
  nand2 gate2138(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2139(.a(s_227), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2140(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2141(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2142(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2465(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2466(.a(gate235inter0), .b(s_274), .O(gate235inter1));
  and2  gate2467(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2468(.a(s_274), .O(gate235inter3));
  inv1  gate2469(.a(s_275), .O(gate235inter4));
  nand2 gate2470(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2471(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2472(.a(G248), .O(gate235inter7));
  inv1  gate2473(.a(G724), .O(gate235inter8));
  nand2 gate2474(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2475(.a(s_275), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2476(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2477(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2478(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate813(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate814(.a(gate239inter0), .b(s_38), .O(gate239inter1));
  and2  gate815(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate816(.a(s_38), .O(gate239inter3));
  inv1  gate817(.a(s_39), .O(gate239inter4));
  nand2 gate818(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate819(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate820(.a(G260), .O(gate239inter7));
  inv1  gate821(.a(G712), .O(gate239inter8));
  nand2 gate822(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate823(.a(s_39), .b(gate239inter3), .O(gate239inter10));
  nor2  gate824(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate825(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate826(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1485(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1486(.a(gate241inter0), .b(s_134), .O(gate241inter1));
  and2  gate1487(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1488(.a(s_134), .O(gate241inter3));
  inv1  gate1489(.a(s_135), .O(gate241inter4));
  nand2 gate1490(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1491(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1492(.a(G242), .O(gate241inter7));
  inv1  gate1493(.a(G730), .O(gate241inter8));
  nand2 gate1494(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1495(.a(s_135), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1496(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1497(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1498(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate2157(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2158(.a(gate242inter0), .b(s_230), .O(gate242inter1));
  and2  gate2159(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2160(.a(s_230), .O(gate242inter3));
  inv1  gate2161(.a(s_231), .O(gate242inter4));
  nand2 gate2162(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2163(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2164(.a(G718), .O(gate242inter7));
  inv1  gate2165(.a(G730), .O(gate242inter8));
  nand2 gate2166(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2167(.a(s_231), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2168(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2169(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2170(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate561(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate562(.a(gate243inter0), .b(s_2), .O(gate243inter1));
  and2  gate563(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate564(.a(s_2), .O(gate243inter3));
  inv1  gate565(.a(s_3), .O(gate243inter4));
  nand2 gate566(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate567(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate568(.a(G245), .O(gate243inter7));
  inv1  gate569(.a(G733), .O(gate243inter8));
  nand2 gate570(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate571(.a(s_3), .b(gate243inter3), .O(gate243inter10));
  nor2  gate572(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate573(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate574(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2339(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2340(.a(gate246inter0), .b(s_256), .O(gate246inter1));
  and2  gate2341(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2342(.a(s_256), .O(gate246inter3));
  inv1  gate2343(.a(s_257), .O(gate246inter4));
  nand2 gate2344(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2345(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2346(.a(G724), .O(gate246inter7));
  inv1  gate2347(.a(G736), .O(gate246inter8));
  nand2 gate2348(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2349(.a(s_257), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2350(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2351(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2352(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate771(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate772(.a(gate247inter0), .b(s_32), .O(gate247inter1));
  and2  gate773(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate774(.a(s_32), .O(gate247inter3));
  inv1  gate775(.a(s_33), .O(gate247inter4));
  nand2 gate776(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate777(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate778(.a(G251), .O(gate247inter7));
  inv1  gate779(.a(G739), .O(gate247inter8));
  nand2 gate780(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate781(.a(s_33), .b(gate247inter3), .O(gate247inter10));
  nor2  gate782(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate783(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate784(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1667(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1668(.a(gate250inter0), .b(s_160), .O(gate250inter1));
  and2  gate1669(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1670(.a(s_160), .O(gate250inter3));
  inv1  gate1671(.a(s_161), .O(gate250inter4));
  nand2 gate1672(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1673(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1674(.a(G706), .O(gate250inter7));
  inv1  gate1675(.a(G742), .O(gate250inter8));
  nand2 gate1676(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1677(.a(s_161), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1678(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1679(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1680(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1219(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1220(.a(gate254inter0), .b(s_96), .O(gate254inter1));
  and2  gate1221(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1222(.a(s_96), .O(gate254inter3));
  inv1  gate1223(.a(s_97), .O(gate254inter4));
  nand2 gate1224(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1225(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1226(.a(G712), .O(gate254inter7));
  inv1  gate1227(.a(G748), .O(gate254inter8));
  nand2 gate1228(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1229(.a(s_97), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1230(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1231(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1232(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate2493(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2494(.a(gate255inter0), .b(s_278), .O(gate255inter1));
  and2  gate2495(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2496(.a(s_278), .O(gate255inter3));
  inv1  gate2497(.a(s_279), .O(gate255inter4));
  nand2 gate2498(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2499(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2500(.a(G263), .O(gate255inter7));
  inv1  gate2501(.a(G751), .O(gate255inter8));
  nand2 gate2502(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2503(.a(s_279), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2504(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2505(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2506(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1975(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1976(.a(gate258inter0), .b(s_204), .O(gate258inter1));
  and2  gate1977(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1978(.a(s_204), .O(gate258inter3));
  inv1  gate1979(.a(s_205), .O(gate258inter4));
  nand2 gate1980(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1981(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1982(.a(G756), .O(gate258inter7));
  inv1  gate1983(.a(G757), .O(gate258inter8));
  nand2 gate1984(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1985(.a(s_205), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1986(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1987(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1988(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate2437(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2438(.a(gate259inter0), .b(s_270), .O(gate259inter1));
  and2  gate2439(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2440(.a(s_270), .O(gate259inter3));
  inv1  gate2441(.a(s_271), .O(gate259inter4));
  nand2 gate2442(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2443(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2444(.a(G758), .O(gate259inter7));
  inv1  gate2445(.a(G759), .O(gate259inter8));
  nand2 gate2446(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2447(.a(s_271), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2448(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2449(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2450(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1191(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1192(.a(gate260inter0), .b(s_92), .O(gate260inter1));
  and2  gate1193(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1194(.a(s_92), .O(gate260inter3));
  inv1  gate1195(.a(s_93), .O(gate260inter4));
  nand2 gate1196(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1197(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1198(.a(G760), .O(gate260inter7));
  inv1  gate1199(.a(G761), .O(gate260inter8));
  nand2 gate1200(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1201(.a(s_93), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1202(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1203(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1204(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2899(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2900(.a(gate261inter0), .b(s_336), .O(gate261inter1));
  and2  gate2901(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2902(.a(s_336), .O(gate261inter3));
  inv1  gate2903(.a(s_337), .O(gate261inter4));
  nand2 gate2904(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2905(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2906(.a(G762), .O(gate261inter7));
  inv1  gate2907(.a(G763), .O(gate261inter8));
  nand2 gate2908(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2909(.a(s_337), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2910(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2911(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2912(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1849(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1850(.a(gate262inter0), .b(s_186), .O(gate262inter1));
  and2  gate1851(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1852(.a(s_186), .O(gate262inter3));
  inv1  gate1853(.a(s_187), .O(gate262inter4));
  nand2 gate1854(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1855(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1856(.a(G764), .O(gate262inter7));
  inv1  gate1857(.a(G765), .O(gate262inter8));
  nand2 gate1858(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1859(.a(s_187), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1860(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1861(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1862(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1261(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1262(.a(gate263inter0), .b(s_102), .O(gate263inter1));
  and2  gate1263(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1264(.a(s_102), .O(gate263inter3));
  inv1  gate1265(.a(s_103), .O(gate263inter4));
  nand2 gate1266(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1267(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1268(.a(G766), .O(gate263inter7));
  inv1  gate1269(.a(G767), .O(gate263inter8));
  nand2 gate1270(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1271(.a(s_103), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1272(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1273(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1274(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2605(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2606(.a(gate265inter0), .b(s_294), .O(gate265inter1));
  and2  gate2607(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2608(.a(s_294), .O(gate265inter3));
  inv1  gate2609(.a(s_295), .O(gate265inter4));
  nand2 gate2610(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2611(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2612(.a(G642), .O(gate265inter7));
  inv1  gate2613(.a(G770), .O(gate265inter8));
  nand2 gate2614(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2615(.a(s_295), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2616(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2617(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2618(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate981(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate982(.a(gate271inter0), .b(s_62), .O(gate271inter1));
  and2  gate983(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate984(.a(s_62), .O(gate271inter3));
  inv1  gate985(.a(s_63), .O(gate271inter4));
  nand2 gate986(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate987(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate988(.a(G660), .O(gate271inter7));
  inv1  gate989(.a(G788), .O(gate271inter8));
  nand2 gate990(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate991(.a(s_63), .b(gate271inter3), .O(gate271inter10));
  nor2  gate992(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate993(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate994(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2423(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2424(.a(gate273inter0), .b(s_268), .O(gate273inter1));
  and2  gate2425(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2426(.a(s_268), .O(gate273inter3));
  inv1  gate2427(.a(s_269), .O(gate273inter4));
  nand2 gate2428(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2429(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2430(.a(G642), .O(gate273inter7));
  inv1  gate2431(.a(G794), .O(gate273inter8));
  nand2 gate2432(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2433(.a(s_269), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2434(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2435(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2436(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2115(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2116(.a(gate275inter0), .b(s_224), .O(gate275inter1));
  and2  gate2117(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2118(.a(s_224), .O(gate275inter3));
  inv1  gate2119(.a(s_225), .O(gate275inter4));
  nand2 gate2120(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2121(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2122(.a(G645), .O(gate275inter7));
  inv1  gate2123(.a(G797), .O(gate275inter8));
  nand2 gate2124(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2125(.a(s_225), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2126(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2127(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2128(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate2087(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2088(.a(gate276inter0), .b(s_220), .O(gate276inter1));
  and2  gate2089(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2090(.a(s_220), .O(gate276inter3));
  inv1  gate2091(.a(s_221), .O(gate276inter4));
  nand2 gate2092(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2093(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2094(.a(G773), .O(gate276inter7));
  inv1  gate2095(.a(G797), .O(gate276inter8));
  nand2 gate2096(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2097(.a(s_221), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2098(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2099(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2100(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1961(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1962(.a(gate278inter0), .b(s_202), .O(gate278inter1));
  and2  gate1963(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1964(.a(s_202), .O(gate278inter3));
  inv1  gate1965(.a(s_203), .O(gate278inter4));
  nand2 gate1966(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1967(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1968(.a(G776), .O(gate278inter7));
  inv1  gate1969(.a(G800), .O(gate278inter8));
  nand2 gate1970(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1971(.a(s_203), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1972(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1973(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1974(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate827(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate828(.a(gate279inter0), .b(s_40), .O(gate279inter1));
  and2  gate829(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate830(.a(s_40), .O(gate279inter3));
  inv1  gate831(.a(s_41), .O(gate279inter4));
  nand2 gate832(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate833(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate834(.a(G651), .O(gate279inter7));
  inv1  gate835(.a(G803), .O(gate279inter8));
  nand2 gate836(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate837(.a(s_41), .b(gate279inter3), .O(gate279inter10));
  nor2  gate838(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate839(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate840(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2395(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2396(.a(gate282inter0), .b(s_264), .O(gate282inter1));
  and2  gate2397(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2398(.a(s_264), .O(gate282inter3));
  inv1  gate2399(.a(s_265), .O(gate282inter4));
  nand2 gate2400(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2401(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2402(.a(G782), .O(gate282inter7));
  inv1  gate2403(.a(G806), .O(gate282inter8));
  nand2 gate2404(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2405(.a(s_265), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2406(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2407(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2408(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2689(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2690(.a(gate285inter0), .b(s_306), .O(gate285inter1));
  and2  gate2691(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2692(.a(s_306), .O(gate285inter3));
  inv1  gate2693(.a(s_307), .O(gate285inter4));
  nand2 gate2694(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2695(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2696(.a(G660), .O(gate285inter7));
  inv1  gate2697(.a(G812), .O(gate285inter8));
  nand2 gate2698(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2699(.a(s_307), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2700(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2701(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2702(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2913(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2914(.a(gate287inter0), .b(s_338), .O(gate287inter1));
  and2  gate2915(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2916(.a(s_338), .O(gate287inter3));
  inv1  gate2917(.a(s_339), .O(gate287inter4));
  nand2 gate2918(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2919(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2920(.a(G663), .O(gate287inter7));
  inv1  gate2921(.a(G815), .O(gate287inter8));
  nand2 gate2922(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2923(.a(s_339), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2924(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2925(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2926(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate2773(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2774(.a(gate288inter0), .b(s_318), .O(gate288inter1));
  and2  gate2775(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2776(.a(s_318), .O(gate288inter3));
  inv1  gate2777(.a(s_319), .O(gate288inter4));
  nand2 gate2778(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2779(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2780(.a(G791), .O(gate288inter7));
  inv1  gate2781(.a(G815), .O(gate288inter8));
  nand2 gate2782(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2783(.a(s_319), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2784(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2785(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2786(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate2297(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2298(.a(gate289inter0), .b(s_250), .O(gate289inter1));
  and2  gate2299(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2300(.a(s_250), .O(gate289inter3));
  inv1  gate2301(.a(s_251), .O(gate289inter4));
  nand2 gate2302(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2303(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2304(.a(G818), .O(gate289inter7));
  inv1  gate2305(.a(G819), .O(gate289inter8));
  nand2 gate2306(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2307(.a(s_251), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2308(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2309(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2310(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2269(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2270(.a(gate291inter0), .b(s_246), .O(gate291inter1));
  and2  gate2271(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2272(.a(s_246), .O(gate291inter3));
  inv1  gate2273(.a(s_247), .O(gate291inter4));
  nand2 gate2274(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2275(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2276(.a(G822), .O(gate291inter7));
  inv1  gate2277(.a(G823), .O(gate291inter8));
  nand2 gate2278(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2279(.a(s_247), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2280(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2281(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2282(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1793(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1794(.a(gate294inter0), .b(s_178), .O(gate294inter1));
  and2  gate1795(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1796(.a(s_178), .O(gate294inter3));
  inv1  gate1797(.a(s_179), .O(gate294inter4));
  nand2 gate1798(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1799(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1800(.a(G832), .O(gate294inter7));
  inv1  gate1801(.a(G833), .O(gate294inter8));
  nand2 gate1802(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1803(.a(s_179), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1804(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1805(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1806(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1177(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1178(.a(gate387inter0), .b(s_90), .O(gate387inter1));
  and2  gate1179(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1180(.a(s_90), .O(gate387inter3));
  inv1  gate1181(.a(s_91), .O(gate387inter4));
  nand2 gate1182(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1183(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1184(.a(G1), .O(gate387inter7));
  inv1  gate1185(.a(G1036), .O(gate387inter8));
  nand2 gate1186(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1187(.a(s_91), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1188(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1189(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1190(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1009(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1010(.a(gate388inter0), .b(s_66), .O(gate388inter1));
  and2  gate1011(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1012(.a(s_66), .O(gate388inter3));
  inv1  gate1013(.a(s_67), .O(gate388inter4));
  nand2 gate1014(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1015(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1016(.a(G2), .O(gate388inter7));
  inv1  gate1017(.a(G1039), .O(gate388inter8));
  nand2 gate1018(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1019(.a(s_67), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1020(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1021(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1022(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate785(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate786(.a(gate389inter0), .b(s_34), .O(gate389inter1));
  and2  gate787(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate788(.a(s_34), .O(gate389inter3));
  inv1  gate789(.a(s_35), .O(gate389inter4));
  nand2 gate790(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate791(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate792(.a(G3), .O(gate389inter7));
  inv1  gate793(.a(G1042), .O(gate389inter8));
  nand2 gate794(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate795(.a(s_35), .b(gate389inter3), .O(gate389inter10));
  nor2  gate796(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate797(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate798(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1919(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1920(.a(gate393inter0), .b(s_196), .O(gate393inter1));
  and2  gate1921(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1922(.a(s_196), .O(gate393inter3));
  inv1  gate1923(.a(s_197), .O(gate393inter4));
  nand2 gate1924(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1925(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1926(.a(G7), .O(gate393inter7));
  inv1  gate1927(.a(G1054), .O(gate393inter8));
  nand2 gate1928(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1929(.a(s_197), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1930(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1931(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1932(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2171(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2172(.a(gate409inter0), .b(s_232), .O(gate409inter1));
  and2  gate2173(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2174(.a(s_232), .O(gate409inter3));
  inv1  gate2175(.a(s_233), .O(gate409inter4));
  nand2 gate2176(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2177(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2178(.a(G23), .O(gate409inter7));
  inv1  gate2179(.a(G1102), .O(gate409inter8));
  nand2 gate2180(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2181(.a(s_233), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2182(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2183(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2184(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1639(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1640(.a(gate412inter0), .b(s_156), .O(gate412inter1));
  and2  gate1641(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1642(.a(s_156), .O(gate412inter3));
  inv1  gate1643(.a(s_157), .O(gate412inter4));
  nand2 gate1644(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1645(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1646(.a(G26), .O(gate412inter7));
  inv1  gate1647(.a(G1111), .O(gate412inter8));
  nand2 gate1648(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1649(.a(s_157), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1650(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1651(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1652(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate2633(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2634(.a(gate413inter0), .b(s_298), .O(gate413inter1));
  and2  gate2635(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2636(.a(s_298), .O(gate413inter3));
  inv1  gate2637(.a(s_299), .O(gate413inter4));
  nand2 gate2638(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2639(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2640(.a(G27), .O(gate413inter7));
  inv1  gate2641(.a(G1114), .O(gate413inter8));
  nand2 gate2642(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2643(.a(s_299), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2644(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2645(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2646(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1625(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1626(.a(gate414inter0), .b(s_154), .O(gate414inter1));
  and2  gate1627(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1628(.a(s_154), .O(gate414inter3));
  inv1  gate1629(.a(s_155), .O(gate414inter4));
  nand2 gate1630(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1631(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1632(.a(G28), .O(gate414inter7));
  inv1  gate1633(.a(G1117), .O(gate414inter8));
  nand2 gate1634(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1635(.a(s_155), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1636(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1637(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1638(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1737(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1738(.a(gate415inter0), .b(s_170), .O(gate415inter1));
  and2  gate1739(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1740(.a(s_170), .O(gate415inter3));
  inv1  gate1741(.a(s_171), .O(gate415inter4));
  nand2 gate1742(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1743(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1744(.a(G29), .O(gate415inter7));
  inv1  gate1745(.a(G1120), .O(gate415inter8));
  nand2 gate1746(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1747(.a(s_171), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1748(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1749(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1750(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1947(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1948(.a(gate417inter0), .b(s_200), .O(gate417inter1));
  and2  gate1949(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1950(.a(s_200), .O(gate417inter3));
  inv1  gate1951(.a(s_201), .O(gate417inter4));
  nand2 gate1952(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1953(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1954(.a(G31), .O(gate417inter7));
  inv1  gate1955(.a(G1126), .O(gate417inter8));
  nand2 gate1956(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1957(.a(s_201), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1958(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1959(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1960(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2535(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2536(.a(gate419inter0), .b(s_284), .O(gate419inter1));
  and2  gate2537(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2538(.a(s_284), .O(gate419inter3));
  inv1  gate2539(.a(s_285), .O(gate419inter4));
  nand2 gate2540(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2541(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2542(.a(G1), .O(gate419inter7));
  inv1  gate2543(.a(G1132), .O(gate419inter8));
  nand2 gate2544(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2545(.a(s_285), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2546(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2547(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2548(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1513(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1514(.a(gate421inter0), .b(s_138), .O(gate421inter1));
  and2  gate1515(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1516(.a(s_138), .O(gate421inter3));
  inv1  gate1517(.a(s_139), .O(gate421inter4));
  nand2 gate1518(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1519(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1520(.a(G2), .O(gate421inter7));
  inv1  gate1521(.a(G1135), .O(gate421inter8));
  nand2 gate1522(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1523(.a(s_139), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1524(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1525(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1526(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2871(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2872(.a(gate424inter0), .b(s_332), .O(gate424inter1));
  and2  gate2873(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2874(.a(s_332), .O(gate424inter3));
  inv1  gate2875(.a(s_333), .O(gate424inter4));
  nand2 gate2876(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2877(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2878(.a(G1042), .O(gate424inter7));
  inv1  gate2879(.a(G1138), .O(gate424inter8));
  nand2 gate2880(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2881(.a(s_333), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2882(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2883(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2884(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1583(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1584(.a(gate425inter0), .b(s_148), .O(gate425inter1));
  and2  gate1585(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1586(.a(s_148), .O(gate425inter3));
  inv1  gate1587(.a(s_149), .O(gate425inter4));
  nand2 gate1588(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1589(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1590(.a(G4), .O(gate425inter7));
  inv1  gate1591(.a(G1141), .O(gate425inter8));
  nand2 gate1592(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1593(.a(s_149), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1594(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1595(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1596(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2045(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2046(.a(gate426inter0), .b(s_214), .O(gate426inter1));
  and2  gate2047(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2048(.a(s_214), .O(gate426inter3));
  inv1  gate2049(.a(s_215), .O(gate426inter4));
  nand2 gate2050(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2051(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2052(.a(G1045), .O(gate426inter7));
  inv1  gate2053(.a(G1141), .O(gate426inter8));
  nand2 gate2054(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2055(.a(s_215), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2056(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2057(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2058(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1695(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1696(.a(gate432inter0), .b(s_164), .O(gate432inter1));
  and2  gate1697(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1698(.a(s_164), .O(gate432inter3));
  inv1  gate1699(.a(s_165), .O(gate432inter4));
  nand2 gate1700(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1701(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1702(.a(G1054), .O(gate432inter7));
  inv1  gate1703(.a(G1150), .O(gate432inter8));
  nand2 gate1704(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1705(.a(s_165), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1706(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1707(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1708(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2059(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2060(.a(gate433inter0), .b(s_216), .O(gate433inter1));
  and2  gate2061(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2062(.a(s_216), .O(gate433inter3));
  inv1  gate2063(.a(s_217), .O(gate433inter4));
  nand2 gate2064(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2065(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2066(.a(G8), .O(gate433inter7));
  inv1  gate2067(.a(G1153), .O(gate433inter8));
  nand2 gate2068(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2069(.a(s_217), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2070(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2071(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2072(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate841(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate842(.a(gate435inter0), .b(s_42), .O(gate435inter1));
  and2  gate843(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate844(.a(s_42), .O(gate435inter3));
  inv1  gate845(.a(s_43), .O(gate435inter4));
  nand2 gate846(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate847(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate848(.a(G9), .O(gate435inter7));
  inv1  gate849(.a(G1156), .O(gate435inter8));
  nand2 gate850(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate851(.a(s_43), .b(gate435inter3), .O(gate435inter10));
  nor2  gate852(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate853(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate854(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1247(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1248(.a(gate436inter0), .b(s_100), .O(gate436inter1));
  and2  gate1249(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1250(.a(s_100), .O(gate436inter3));
  inv1  gate1251(.a(s_101), .O(gate436inter4));
  nand2 gate1252(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1253(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1254(.a(G1060), .O(gate436inter7));
  inv1  gate1255(.a(G1156), .O(gate436inter8));
  nand2 gate1256(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1257(.a(s_101), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1258(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1259(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1260(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate701(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate702(.a(gate438inter0), .b(s_22), .O(gate438inter1));
  and2  gate703(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate704(.a(s_22), .O(gate438inter3));
  inv1  gate705(.a(s_23), .O(gate438inter4));
  nand2 gate706(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate707(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate708(.a(G1063), .O(gate438inter7));
  inv1  gate709(.a(G1159), .O(gate438inter8));
  nand2 gate710(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate711(.a(s_23), .b(gate438inter3), .O(gate438inter10));
  nor2  gate712(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate713(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate714(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1765(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1766(.a(gate443inter0), .b(s_174), .O(gate443inter1));
  and2  gate1767(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1768(.a(s_174), .O(gate443inter3));
  inv1  gate1769(.a(s_175), .O(gate443inter4));
  nand2 gate1770(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1771(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1772(.a(G13), .O(gate443inter7));
  inv1  gate1773(.a(G1168), .O(gate443inter8));
  nand2 gate1774(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1775(.a(s_175), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1776(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1777(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1778(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2409(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2410(.a(gate444inter0), .b(s_266), .O(gate444inter1));
  and2  gate2411(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2412(.a(s_266), .O(gate444inter3));
  inv1  gate2413(.a(s_267), .O(gate444inter4));
  nand2 gate2414(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2415(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2416(.a(G1072), .O(gate444inter7));
  inv1  gate2417(.a(G1168), .O(gate444inter8));
  nand2 gate2418(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2419(.a(s_267), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2420(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2421(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2422(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate2241(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2242(.a(gate445inter0), .b(s_242), .O(gate445inter1));
  and2  gate2243(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2244(.a(s_242), .O(gate445inter3));
  inv1  gate2245(.a(s_243), .O(gate445inter4));
  nand2 gate2246(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2247(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2248(.a(G14), .O(gate445inter7));
  inv1  gate2249(.a(G1171), .O(gate445inter8));
  nand2 gate2250(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2251(.a(s_243), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2252(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2253(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2254(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate2885(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2886(.a(gate449inter0), .b(s_334), .O(gate449inter1));
  and2  gate2887(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2888(.a(s_334), .O(gate449inter3));
  inv1  gate2889(.a(s_335), .O(gate449inter4));
  nand2 gate2890(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2891(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2892(.a(G16), .O(gate449inter7));
  inv1  gate2893(.a(G1177), .O(gate449inter8));
  nand2 gate2894(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2895(.a(s_335), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2896(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2897(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2898(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2031(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2032(.a(gate451inter0), .b(s_212), .O(gate451inter1));
  and2  gate2033(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2034(.a(s_212), .O(gate451inter3));
  inv1  gate2035(.a(s_213), .O(gate451inter4));
  nand2 gate2036(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2037(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2038(.a(G17), .O(gate451inter7));
  inv1  gate2039(.a(G1180), .O(gate451inter8));
  nand2 gate2040(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2041(.a(s_213), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2042(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2043(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2044(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1331(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1332(.a(gate452inter0), .b(s_112), .O(gate452inter1));
  and2  gate1333(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1334(.a(s_112), .O(gate452inter3));
  inv1  gate1335(.a(s_113), .O(gate452inter4));
  nand2 gate1336(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1337(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1338(.a(G1084), .O(gate452inter7));
  inv1  gate1339(.a(G1180), .O(gate452inter8));
  nand2 gate1340(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1341(.a(s_113), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1342(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1343(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1344(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1023(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1024(.a(gate456inter0), .b(s_68), .O(gate456inter1));
  and2  gate1025(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1026(.a(s_68), .O(gate456inter3));
  inv1  gate1027(.a(s_69), .O(gate456inter4));
  nand2 gate1028(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1029(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1030(.a(G1090), .O(gate456inter7));
  inv1  gate1031(.a(G1186), .O(gate456inter8));
  nand2 gate1032(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1033(.a(s_69), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1034(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1035(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1036(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate953(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate954(.a(gate457inter0), .b(s_58), .O(gate457inter1));
  and2  gate955(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate956(.a(s_58), .O(gate457inter3));
  inv1  gate957(.a(s_59), .O(gate457inter4));
  nand2 gate958(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate959(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate960(.a(G20), .O(gate457inter7));
  inv1  gate961(.a(G1189), .O(gate457inter8));
  nand2 gate962(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate963(.a(s_59), .b(gate457inter3), .O(gate457inter10));
  nor2  gate964(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate965(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate966(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2745(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2746(.a(gate460inter0), .b(s_314), .O(gate460inter1));
  and2  gate2747(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2748(.a(s_314), .O(gate460inter3));
  inv1  gate2749(.a(s_315), .O(gate460inter4));
  nand2 gate2750(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2751(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2752(.a(G1096), .O(gate460inter7));
  inv1  gate2753(.a(G1192), .O(gate460inter8));
  nand2 gate2754(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2755(.a(s_315), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2756(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2757(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2758(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1415(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1416(.a(gate464inter0), .b(s_124), .O(gate464inter1));
  and2  gate1417(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1418(.a(s_124), .O(gate464inter3));
  inv1  gate1419(.a(s_125), .O(gate464inter4));
  nand2 gate1420(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1421(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1422(.a(G1102), .O(gate464inter7));
  inv1  gate1423(.a(G1198), .O(gate464inter8));
  nand2 gate1424(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1425(.a(s_125), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1426(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1427(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1428(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate967(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate968(.a(gate465inter0), .b(s_60), .O(gate465inter1));
  and2  gate969(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate970(.a(s_60), .O(gate465inter3));
  inv1  gate971(.a(s_61), .O(gate465inter4));
  nand2 gate972(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate973(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate974(.a(G24), .O(gate465inter7));
  inv1  gate975(.a(G1201), .O(gate465inter8));
  nand2 gate976(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate977(.a(s_61), .b(gate465inter3), .O(gate465inter10));
  nor2  gate978(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate979(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate980(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate589(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate590(.a(gate469inter0), .b(s_6), .O(gate469inter1));
  and2  gate591(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate592(.a(s_6), .O(gate469inter3));
  inv1  gate593(.a(s_7), .O(gate469inter4));
  nand2 gate594(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate595(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate596(.a(G26), .O(gate469inter7));
  inv1  gate597(.a(G1207), .O(gate469inter8));
  nand2 gate598(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate599(.a(s_7), .b(gate469inter3), .O(gate469inter10));
  nor2  gate600(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate601(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate602(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2101(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2102(.a(gate470inter0), .b(s_222), .O(gate470inter1));
  and2  gate2103(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2104(.a(s_222), .O(gate470inter3));
  inv1  gate2105(.a(s_223), .O(gate470inter4));
  nand2 gate2106(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2107(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2108(.a(G1111), .O(gate470inter7));
  inv1  gate2109(.a(G1207), .O(gate470inter8));
  nand2 gate2110(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2111(.a(s_223), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2112(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2113(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2114(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1835(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1836(.a(gate471inter0), .b(s_184), .O(gate471inter1));
  and2  gate1837(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1838(.a(s_184), .O(gate471inter3));
  inv1  gate1839(.a(s_185), .O(gate471inter4));
  nand2 gate1840(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1841(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1842(.a(G27), .O(gate471inter7));
  inv1  gate1843(.a(G1210), .O(gate471inter8));
  nand2 gate1844(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1845(.a(s_185), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1846(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1847(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1848(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2647(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2648(.a(gate475inter0), .b(s_300), .O(gate475inter1));
  and2  gate2649(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2650(.a(s_300), .O(gate475inter3));
  inv1  gate2651(.a(s_301), .O(gate475inter4));
  nand2 gate2652(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2653(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2654(.a(G29), .O(gate475inter7));
  inv1  gate2655(.a(G1216), .O(gate475inter8));
  nand2 gate2656(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2657(.a(s_301), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2658(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2659(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2660(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1065(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1066(.a(gate477inter0), .b(s_74), .O(gate477inter1));
  and2  gate1067(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1068(.a(s_74), .O(gate477inter3));
  inv1  gate1069(.a(s_75), .O(gate477inter4));
  nand2 gate1070(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1071(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1072(.a(G30), .O(gate477inter7));
  inv1  gate1073(.a(G1219), .O(gate477inter8));
  nand2 gate1074(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1075(.a(s_75), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1076(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1077(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1078(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate687(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate688(.a(gate478inter0), .b(s_20), .O(gate478inter1));
  and2  gate689(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate690(.a(s_20), .O(gate478inter3));
  inv1  gate691(.a(s_21), .O(gate478inter4));
  nand2 gate692(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate693(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate694(.a(G1123), .O(gate478inter7));
  inv1  gate695(.a(G1219), .O(gate478inter8));
  nand2 gate696(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate697(.a(s_21), .b(gate478inter3), .O(gate478inter10));
  nor2  gate698(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate699(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate700(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate995(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate996(.a(gate481inter0), .b(s_64), .O(gate481inter1));
  and2  gate997(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate998(.a(s_64), .O(gate481inter3));
  inv1  gate999(.a(s_65), .O(gate481inter4));
  nand2 gate1000(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1001(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1002(.a(G32), .O(gate481inter7));
  inv1  gate1003(.a(G1225), .O(gate481inter8));
  nand2 gate1004(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1005(.a(s_65), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1006(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1007(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1008(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate2227(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2228(.a(gate484inter0), .b(s_240), .O(gate484inter1));
  and2  gate2229(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2230(.a(s_240), .O(gate484inter3));
  inv1  gate2231(.a(s_241), .O(gate484inter4));
  nand2 gate2232(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2233(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2234(.a(G1230), .O(gate484inter7));
  inv1  gate2235(.a(G1231), .O(gate484inter8));
  nand2 gate2236(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2237(.a(s_241), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2238(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2239(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2240(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate799(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate800(.a(gate491inter0), .b(s_36), .O(gate491inter1));
  and2  gate801(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate802(.a(s_36), .O(gate491inter3));
  inv1  gate803(.a(s_37), .O(gate491inter4));
  nand2 gate804(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate805(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate806(.a(G1244), .O(gate491inter7));
  inv1  gate807(.a(G1245), .O(gate491inter8));
  nand2 gate808(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate809(.a(s_37), .b(gate491inter3), .O(gate491inter10));
  nor2  gate810(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate811(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate812(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1289(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1290(.a(gate492inter0), .b(s_106), .O(gate492inter1));
  and2  gate1291(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1292(.a(s_106), .O(gate492inter3));
  inv1  gate1293(.a(s_107), .O(gate492inter4));
  nand2 gate1294(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1295(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1296(.a(G1246), .O(gate492inter7));
  inv1  gate1297(.a(G1247), .O(gate492inter8));
  nand2 gate1298(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1299(.a(s_107), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1300(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1301(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1302(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2759(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2760(.a(gate493inter0), .b(s_316), .O(gate493inter1));
  and2  gate2761(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2762(.a(s_316), .O(gate493inter3));
  inv1  gate2763(.a(s_317), .O(gate493inter4));
  nand2 gate2764(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2765(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2766(.a(G1248), .O(gate493inter7));
  inv1  gate2767(.a(G1249), .O(gate493inter8));
  nand2 gate2768(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2769(.a(s_317), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2770(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2771(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2772(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1345(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1346(.a(gate496inter0), .b(s_114), .O(gate496inter1));
  and2  gate1347(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1348(.a(s_114), .O(gate496inter3));
  inv1  gate1349(.a(s_115), .O(gate496inter4));
  nand2 gate1350(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1351(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1352(.a(G1254), .O(gate496inter7));
  inv1  gate1353(.a(G1255), .O(gate496inter8));
  nand2 gate1354(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1355(.a(s_115), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1356(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1357(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1358(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate869(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate870(.a(gate498inter0), .b(s_46), .O(gate498inter1));
  and2  gate871(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate872(.a(s_46), .O(gate498inter3));
  inv1  gate873(.a(s_47), .O(gate498inter4));
  nand2 gate874(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate875(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate876(.a(G1258), .O(gate498inter7));
  inv1  gate877(.a(G1259), .O(gate498inter8));
  nand2 gate878(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate879(.a(s_47), .b(gate498inter3), .O(gate498inter10));
  nor2  gate880(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate881(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate882(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1149(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1150(.a(gate501inter0), .b(s_86), .O(gate501inter1));
  and2  gate1151(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1152(.a(s_86), .O(gate501inter3));
  inv1  gate1153(.a(s_87), .O(gate501inter4));
  nand2 gate1154(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1155(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1156(.a(G1264), .O(gate501inter7));
  inv1  gate1157(.a(G1265), .O(gate501inter8));
  nand2 gate1158(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1159(.a(s_87), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1160(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1161(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1162(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1051(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1052(.a(gate502inter0), .b(s_72), .O(gate502inter1));
  and2  gate1053(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1054(.a(s_72), .O(gate502inter3));
  inv1  gate1055(.a(s_73), .O(gate502inter4));
  nand2 gate1056(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1057(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1058(.a(G1266), .O(gate502inter7));
  inv1  gate1059(.a(G1267), .O(gate502inter8));
  nand2 gate1060(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1061(.a(s_73), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1062(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1063(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1064(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1471(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1472(.a(gate506inter0), .b(s_132), .O(gate506inter1));
  and2  gate1473(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1474(.a(s_132), .O(gate506inter3));
  inv1  gate1475(.a(s_133), .O(gate506inter4));
  nand2 gate1476(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1477(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1478(.a(G1274), .O(gate506inter7));
  inv1  gate1479(.a(G1275), .O(gate506inter8));
  nand2 gate1480(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1481(.a(s_133), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1482(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1483(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1484(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1093(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1094(.a(gate512inter0), .b(s_78), .O(gate512inter1));
  and2  gate1095(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1096(.a(s_78), .O(gate512inter3));
  inv1  gate1097(.a(s_79), .O(gate512inter4));
  nand2 gate1098(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1099(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1100(.a(G1286), .O(gate512inter7));
  inv1  gate1101(.a(G1287), .O(gate512inter8));
  nand2 gate1102(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1103(.a(s_79), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1104(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1105(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1106(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule