module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate824inter0, gate824inter1, gate824inter2, gate824inter3, gate824inter4, gate824inter5, gate824inter6, gate824inter7, gate824inter8, gate824inter9, gate824inter10, gate824inter11, gate824inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate876inter0, gate876inter1, gate876inter2, gate876inter3, gate876inter4, gate876inter5, gate876inter6, gate876inter7, gate876inter8, gate876inter9, gate876inter10, gate876inter11, gate876inter12, gate673inter0, gate673inter1, gate673inter2, gate673inter3, gate673inter4, gate673inter5, gate673inter6, gate673inter7, gate673inter8, gate673inter9, gate673inter10, gate673inter11, gate673inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate801inter0, gate801inter1, gate801inter2, gate801inter3, gate801inter4, gate801inter5, gate801inter6, gate801inter7, gate801inter8, gate801inter9, gate801inter10, gate801inter11, gate801inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate805inter0, gate805inter1, gate805inter2, gate805inter3, gate805inter4, gate805inter5, gate805inter6, gate805inter7, gate805inter8, gate805inter9, gate805inter10, gate805inter11, gate805inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate593inter0, gate593inter1, gate593inter2, gate593inter3, gate593inter4, gate593inter5, gate593inter6, gate593inter7, gate593inter8, gate593inter9, gate593inter10, gate593inter11, gate593inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate607inter0, gate607inter1, gate607inter2, gate607inter3, gate607inter4, gate607inter5, gate607inter6, gate607inter7, gate607inter8, gate607inter9, gate607inter10, gate607inter11, gate607inter12, gate765inter0, gate765inter1, gate765inter2, gate765inter3, gate765inter4, gate765inter5, gate765inter6, gate765inter7, gate765inter8, gate765inter9, gate765inter10, gate765inter11, gate765inter12, gate320inter0, gate320inter1, gate320inter2, gate320inter3, gate320inter4, gate320inter5, gate320inter6, gate320inter7, gate320inter8, gate320inter9, gate320inter10, gate320inter11, gate320inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate794inter0, gate794inter1, gate794inter2, gate794inter3, gate794inter4, gate794inter5, gate794inter6, gate794inter7, gate794inter8, gate794inter9, gate794inter10, gate794inter11, gate794inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate767inter0, gate767inter1, gate767inter2, gate767inter3, gate767inter4, gate767inter5, gate767inter6, gate767inter7, gate767inter8, gate767inter9, gate767inter10, gate767inter11, gate767inter12, gate527inter0, gate527inter1, gate527inter2, gate527inter3, gate527inter4, gate527inter5, gate527inter6, gate527inter7, gate527inter8, gate527inter9, gate527inter10, gate527inter11, gate527inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate370inter0, gate370inter1, gate370inter2, gate370inter3, gate370inter4, gate370inter5, gate370inter6, gate370inter7, gate370inter8, gate370inter9, gate370inter10, gate370inter11, gate370inter12, gate374inter0, gate374inter1, gate374inter2, gate374inter3, gate374inter4, gate374inter5, gate374inter6, gate374inter7, gate374inter8, gate374inter9, gate374inter10, gate374inter11, gate374inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate863inter0, gate863inter1, gate863inter2, gate863inter3, gate863inter4, gate863inter5, gate863inter6, gate863inter7, gate863inter8, gate863inter9, gate863inter10, gate863inter11, gate863inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate523inter0, gate523inter1, gate523inter2, gate523inter3, gate523inter4, gate523inter5, gate523inter6, gate523inter7, gate523inter8, gate523inter9, gate523inter10, gate523inter11, gate523inter12, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate663inter0, gate663inter1, gate663inter2, gate663inter3, gate663inter4, gate663inter5, gate663inter6, gate663inter7, gate663inter8, gate663inter9, gate663inter10, gate663inter11, gate663inter12, gate797inter0, gate797inter1, gate797inter2, gate797inter3, gate797inter4, gate797inter5, gate797inter6, gate797inter7, gate797inter8, gate797inter9, gate797inter10, gate797inter11, gate797inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate539inter0, gate539inter1, gate539inter2, gate539inter3, gate539inter4, gate539inter5, gate539inter6, gate539inter7, gate539inter8, gate539inter9, gate539inter10, gate539inter11, gate539inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate862inter0, gate862inter1, gate862inter2, gate862inter3, gate862inter4, gate862inter5, gate862inter6, gate862inter7, gate862inter8, gate862inter9, gate862inter10, gate862inter11, gate862inter12, gate686inter0, gate686inter1, gate686inter2, gate686inter3, gate686inter4, gate686inter5, gate686inter6, gate686inter7, gate686inter8, gate686inter9, gate686inter10, gate686inter11, gate686inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate851inter0, gate851inter1, gate851inter2, gate851inter3, gate851inter4, gate851inter5, gate851inter6, gate851inter7, gate851inter8, gate851inter9, gate851inter10, gate851inter11, gate851inter12, gate632inter0, gate632inter1, gate632inter2, gate632inter3, gate632inter4, gate632inter5, gate632inter6, gate632inter7, gate632inter8, gate632inter9, gate632inter10, gate632inter11, gate632inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate625inter0, gate625inter1, gate625inter2, gate625inter3, gate625inter4, gate625inter5, gate625inter6, gate625inter7, gate625inter8, gate625inter9, gate625inter10, gate625inter11, gate625inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate780inter0, gate780inter1, gate780inter2, gate780inter3, gate780inter4, gate780inter5, gate780inter6, gate780inter7, gate780inter8, gate780inter9, gate780inter10, gate780inter11, gate780inter12, gate631inter0, gate631inter1, gate631inter2, gate631inter3, gate631inter4, gate631inter5, gate631inter6, gate631inter7, gate631inter8, gate631inter9, gate631inter10, gate631inter11, gate631inter12, gate758inter0, gate758inter1, gate758inter2, gate758inter3, gate758inter4, gate758inter5, gate758inter6, gate758inter7, gate758inter8, gate758inter9, gate758inter10, gate758inter11, gate758inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate543inter0, gate543inter1, gate543inter2, gate543inter3, gate543inter4, gate543inter5, gate543inter6, gate543inter7, gate543inter8, gate543inter9, gate543inter10, gate543inter11, gate543inter12, gate866inter0, gate866inter1, gate866inter2, gate866inter3, gate866inter4, gate866inter5, gate866inter6, gate866inter7, gate866inter8, gate866inter9, gate866inter10, gate866inter11, gate866inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate355inter0, gate355inter1, gate355inter2, gate355inter3, gate355inter4, gate355inter5, gate355inter6, gate355inter7, gate355inter8, gate355inter9, gate355inter10, gate355inter11, gate355inter12, gate669inter0, gate669inter1, gate669inter2, gate669inter3, gate669inter4, gate669inter5, gate669inter6, gate669inter7, gate669inter8, gate669inter9, gate669inter10, gate669inter11, gate669inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate516inter0, gate516inter1, gate516inter2, gate516inter3, gate516inter4, gate516inter5, gate516inter6, gate516inter7, gate516inter8, gate516inter9, gate516inter10, gate516inter11, gate516inter12, gate368inter0, gate368inter1, gate368inter2, gate368inter3, gate368inter4, gate368inter5, gate368inter6, gate368inter7, gate368inter8, gate368inter9, gate368inter10, gate368inter11, gate368inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate775inter0, gate775inter1, gate775inter2, gate775inter3, gate775inter4, gate775inter5, gate775inter6, gate775inter7, gate775inter8, gate775inter9, gate775inter10, gate775inter11, gate775inter12, gate875inter0, gate875inter1, gate875inter2, gate875inter3, gate875inter4, gate875inter5, gate875inter6, gate875inter7, gate875inter8, gate875inter9, gate875inter10, gate875inter11, gate875inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate807inter0, gate807inter1, gate807inter2, gate807inter3, gate807inter4, gate807inter5, gate807inter6, gate807inter7, gate807inter8, gate807inter9, gate807inter10, gate807inter11, gate807inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate338inter0, gate338inter1, gate338inter2, gate338inter3, gate338inter4, gate338inter5, gate338inter6, gate338inter7, gate338inter8, gate338inter9, gate338inter10, gate338inter11, gate338inter12, gate771inter0, gate771inter1, gate771inter2, gate771inter3, gate771inter4, gate771inter5, gate771inter6, gate771inter7, gate771inter8, gate771inter9, gate771inter10, gate771inter11, gate771inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate818inter0, gate818inter1, gate818inter2, gate818inter3, gate818inter4, gate818inter5, gate818inter6, gate818inter7, gate818inter8, gate818inter9, gate818inter10, gate818inter11, gate818inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate675inter0, gate675inter1, gate675inter2, gate675inter3, gate675inter4, gate675inter5, gate675inter6, gate675inter7, gate675inter8, gate675inter9, gate675inter10, gate675inter11, gate675inter12, gate366inter0, gate366inter1, gate366inter2, gate366inter3, gate366inter4, gate366inter5, gate366inter6, gate366inter7, gate366inter8, gate366inter9, gate366inter10, gate366inter11, gate366inter12, gate676inter0, gate676inter1, gate676inter2, gate676inter3, gate676inter4, gate676inter5, gate676inter6, gate676inter7, gate676inter8, gate676inter9, gate676inter10, gate676inter11, gate676inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate642inter0, gate642inter1, gate642inter2, gate642inter3, gate642inter4, gate642inter5, gate642inter6, gate642inter7, gate642inter8, gate642inter9, gate642inter10, gate642inter11, gate642inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate325inter0, gate325inter1, gate325inter2, gate325inter3, gate325inter4, gate325inter5, gate325inter6, gate325inter7, gate325inter8, gate325inter9, gate325inter10, gate325inter11, gate325inter12, gate623inter0, gate623inter1, gate623inter2, gate623inter3, gate623inter4, gate623inter5, gate623inter6, gate623inter7, gate623inter8, gate623inter9, gate623inter10, gate623inter11, gate623inter12, gate528inter0, gate528inter1, gate528inter2, gate528inter3, gate528inter4, gate528inter5, gate528inter6, gate528inter7, gate528inter8, gate528inter9, gate528inter10, gate528inter11, gate528inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate817inter0, gate817inter1, gate817inter2, gate817inter3, gate817inter4, gate817inter5, gate817inter6, gate817inter7, gate817inter8, gate817inter9, gate817inter10, gate817inter11, gate817inter12, gate802inter0, gate802inter1, gate802inter2, gate802inter3, gate802inter4, gate802inter5, gate802inter6, gate802inter7, gate802inter8, gate802inter9, gate802inter10, gate802inter11, gate802inter12, gate798inter0, gate798inter1, gate798inter2, gate798inter3, gate798inter4, gate798inter5, gate798inter6, gate798inter7, gate798inter8, gate798inter9, gate798inter10, gate798inter11, gate798inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate795inter0, gate795inter1, gate795inter2, gate795inter3, gate795inter4, gate795inter5, gate795inter6, gate795inter7, gate795inter8, gate795inter9, gate795inter10, gate795inter11, gate795inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate879inter0, gate879inter1, gate879inter2, gate879inter3, gate879inter4, gate879inter5, gate879inter6, gate879inter7, gate879inter8, gate879inter9, gate879inter10, gate879inter11, gate879inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate608inter0, gate608inter1, gate608inter2, gate608inter3, gate608inter4, gate608inter5, gate608inter6, gate608inter7, gate608inter8, gate608inter9, gate608inter10, gate608inter11, gate608inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate812inter0, gate812inter1, gate812inter2, gate812inter3, gate812inter4, gate812inter5, gate812inter6, gate812inter7, gate812inter8, gate812inter9, gate812inter10, gate812inter11, gate812inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate637inter0, gate637inter1, gate637inter2, gate637inter3, gate637inter4, gate637inter5, gate637inter6, gate637inter7, gate637inter8, gate637inter9, gate637inter10, gate637inter11, gate637inter12, gate345inter0, gate345inter1, gate345inter2, gate345inter3, gate345inter4, gate345inter5, gate345inter6, gate345inter7, gate345inter8, gate345inter9, gate345inter10, gate345inter11, gate345inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate561inter0, gate561inter1, gate561inter2, gate561inter3, gate561inter4, gate561inter5, gate561inter6, gate561inter7, gate561inter8, gate561inter9, gate561inter10, gate561inter11, gate561inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );

  xor2  gate2659(.a(N331), .b(N306), .O(gate78inter0));
  nand2 gate2660(.a(gate78inter0), .b(s_254), .O(gate78inter1));
  and2  gate2661(.a(N331), .b(N306), .O(gate78inter2));
  inv1  gate2662(.a(s_254), .O(gate78inter3));
  inv1  gate2663(.a(s_255), .O(gate78inter4));
  nand2 gate2664(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2665(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2666(.a(N306), .O(gate78inter7));
  inv1  gate2667(.a(N331), .O(gate78inter8));
  nand2 gate2668(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2669(.a(s_255), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2670(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2671(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2672(.a(gate78inter12), .b(gate78inter1), .O(N553));
nand2 gate79( .a(N306), .b(N331), .O(N554) );

  xor2  gate1441(.a(N331), .b(N306), .O(gate80inter0));
  nand2 gate1442(.a(gate80inter0), .b(s_80), .O(gate80inter1));
  and2  gate1443(.a(N331), .b(N306), .O(gate80inter2));
  inv1  gate1444(.a(s_80), .O(gate80inter3));
  inv1  gate1445(.a(s_81), .O(gate80inter4));
  nand2 gate1446(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1447(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1448(.a(N306), .O(gate80inter7));
  inv1  gate1449(.a(N331), .O(gate80inter8));
  nand2 gate1450(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1451(.a(s_81), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1452(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1453(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1454(.a(gate80inter12), .b(gate80inter1), .O(N555));
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate1231(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate1232(.a(gate96inter0), .b(s_50), .O(gate96inter1));
  and2  gate1233(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate1234(.a(s_50), .O(gate96inter3));
  inv1  gate1235(.a(s_51), .O(gate96inter4));
  nand2 gate1236(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1237(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1238(.a(N326), .O(gate96inter7));
  inv1  gate1239(.a(N277), .O(gate96inter8));
  nand2 gate1240(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1241(.a(s_51), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1242(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1243(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1244(.a(gate96inter12), .b(gate96inter1), .O(N601));
nand2 gate97( .a(N326), .b(N280), .O(N602) );

  xor2  gate2463(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate2464(.a(gate98inter0), .b(s_226), .O(gate98inter1));
  and2  gate2465(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate2466(.a(s_226), .O(gate98inter3));
  inv1  gate2467(.a(s_227), .O(gate98inter4));
  nand2 gate2468(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2469(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2470(.a(N260), .O(gate98inter7));
  inv1  gate2471(.a(N72), .O(gate98inter8));
  nand2 gate2472(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2473(.a(s_227), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2474(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2475(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2476(.a(gate98inter12), .b(gate98inter1), .O(N603));

  xor2  gate2407(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate2408(.a(gate99inter0), .b(s_218), .O(gate99inter1));
  and2  gate2409(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate2410(.a(s_218), .O(gate99inter3));
  inv1  gate2411(.a(s_219), .O(gate99inter4));
  nand2 gate2412(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2413(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2414(.a(N260), .O(gate99inter7));
  inv1  gate2415(.a(N300), .O(gate99inter8));
  nand2 gate2416(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2417(.a(s_219), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2418(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2419(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2420(.a(gate99inter12), .b(gate99inter1), .O(N608));
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );

  xor2  gate2281(.a(N612), .b(N49), .O(gate162inter0));
  nand2 gate2282(.a(gate162inter0), .b(s_200), .O(gate162inter1));
  and2  gate2283(.a(N612), .b(N49), .O(gate162inter2));
  inv1  gate2284(.a(s_200), .O(gate162inter3));
  inv1  gate2285(.a(s_201), .O(gate162inter4));
  nand2 gate2286(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2287(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2288(.a(N49), .O(gate162inter7));
  inv1  gate2289(.a(N612), .O(gate162inter8));
  nand2 gate2290(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2291(.a(s_201), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2292(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2293(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2294(.a(gate162inter12), .b(gate162inter1), .O(N907));
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );

  xor2  gate2295(.a(N888), .b(N619), .O(gate233inter0));
  nand2 gate2296(.a(gate233inter0), .b(s_202), .O(gate233inter1));
  and2  gate2297(.a(N888), .b(N619), .O(gate233inter2));
  inv1  gate2298(.a(s_202), .O(gate233inter3));
  inv1  gate2299(.a(s_203), .O(gate233inter4));
  nand2 gate2300(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2301(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2302(.a(N619), .O(gate233inter7));
  inv1  gate2303(.a(N888), .O(gate233inter8));
  nand2 gate2304(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2305(.a(s_203), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2306(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2307(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2308(.a(gate233inter12), .b(gate233inter1), .O(N1054));
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );

  xor2  gate1511(.a(N989), .b(N718), .O(gate240inter0));
  nand2 gate1512(.a(gate240inter0), .b(s_90), .O(gate240inter1));
  and2  gate1513(.a(N989), .b(N718), .O(gate240inter2));
  inv1  gate1514(.a(s_90), .O(gate240inter3));
  inv1  gate1515(.a(s_91), .O(gate240inter4));
  nand2 gate1516(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1517(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1518(.a(N718), .O(gate240inter7));
  inv1  gate1519(.a(N989), .O(gate240inter8));
  nand2 gate1520(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1521(.a(s_91), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1522(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1523(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1524(.a(gate240inter12), .b(gate240inter1), .O(N1120));

  xor2  gate1189(.a(N991), .b(N727), .O(gate241inter0));
  nand2 gate1190(.a(gate241inter0), .b(s_44), .O(gate241inter1));
  and2  gate1191(.a(N991), .b(N727), .O(gate241inter2));
  inv1  gate1192(.a(s_44), .O(gate241inter3));
  inv1  gate1193(.a(s_45), .O(gate241inter4));
  nand2 gate1194(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1195(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1196(.a(N727), .O(gate241inter7));
  inv1  gate1197(.a(N991), .O(gate241inter8));
  nand2 gate1198(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1199(.a(s_45), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1200(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1201(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1202(.a(gate241inter12), .b(gate241inter1), .O(N1121));

  xor2  gate1609(.a(N992), .b(N724), .O(gate242inter0));
  nand2 gate1610(.a(gate242inter0), .b(s_104), .O(gate242inter1));
  and2  gate1611(.a(N992), .b(N724), .O(gate242inter2));
  inv1  gate1612(.a(s_104), .O(gate242inter3));
  inv1  gate1613(.a(s_105), .O(gate242inter4));
  nand2 gate1614(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1615(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1616(.a(N724), .O(gate242inter7));
  inv1  gate1617(.a(N992), .O(gate242inter8));
  nand2 gate1618(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1619(.a(s_105), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1620(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1621(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1622(.a(gate242inter12), .b(gate242inter1), .O(N1122));

  xor2  gate937(.a(N1002), .b(N739), .O(gate243inter0));
  nand2 gate938(.a(gate243inter0), .b(s_8), .O(gate243inter1));
  and2  gate939(.a(N1002), .b(N739), .O(gate243inter2));
  inv1  gate940(.a(s_8), .O(gate243inter3));
  inv1  gate941(.a(s_9), .O(gate243inter4));
  nand2 gate942(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate943(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate944(.a(N739), .O(gate243inter7));
  inv1  gate945(.a(N1002), .O(gate243inter8));
  nand2 gate946(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate947(.a(s_9), .b(gate243inter3), .O(gate243inter10));
  nor2  gate948(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate949(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate950(.a(gate243inter12), .b(gate243inter1), .O(N1128));
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );

  xor2  gate1525(.a(N1008), .b(N751), .O(gate247inter0));
  nand2 gate1526(.a(gate247inter0), .b(s_92), .O(gate247inter1));
  and2  gate1527(.a(N1008), .b(N751), .O(gate247inter2));
  inv1  gate1528(.a(s_92), .O(gate247inter3));
  inv1  gate1529(.a(s_93), .O(gate247inter4));
  nand2 gate1530(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1531(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1532(.a(N751), .O(gate247inter7));
  inv1  gate1533(.a(N1008), .O(gate247inter8));
  nand2 gate1534(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1535(.a(s_93), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1536(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1537(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1538(.a(gate247inter12), .b(gate247inter1), .O(N1132));
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );

  xor2  gate2267(.a(N892), .b(N985), .O(gate261inter0));
  nand2 gate2268(.a(gate261inter0), .b(s_198), .O(gate261inter1));
  and2  gate2269(.a(N892), .b(N985), .O(gate261inter2));
  inv1  gate2270(.a(s_198), .O(gate261inter3));
  inv1  gate2271(.a(s_199), .O(gate261inter4));
  nand2 gate2272(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2273(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2274(.a(N985), .O(gate261inter7));
  inv1  gate2275(.a(N892), .O(gate261inter8));
  nand2 gate2276(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2277(.a(s_199), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2278(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2279(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2280(.a(gate261inter12), .b(gate261inter1), .O(N1160));
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate1273(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate1274(.a(gate268inter0), .b(s_56), .O(gate268inter1));
  and2  gate1275(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate1276(.a(s_56), .O(gate268inter3));
  inv1  gate1277(.a(s_57), .O(gate268inter4));
  nand2 gate1278(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1279(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1280(.a(N921), .O(gate268inter7));
  inv1  gate1281(.a(N923), .O(gate268inter8));
  nand2 gate1282(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1283(.a(s_57), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1284(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1285(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1286(.a(gate268inter12), .b(gate268inter1), .O(N1171));
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate1749(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate1750(.a(gate277inter0), .b(s_124), .O(gate277inter1));
  and2  gate1751(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate1752(.a(s_124), .O(gate277inter3));
  inv1  gate1753(.a(s_125), .O(gate277inter4));
  nand2 gate1754(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1755(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1756(.a(N1019), .O(gate277inter7));
  inv1  gate1757(.a(N950), .O(gate277inter8));
  nand2 gate1758(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1759(.a(s_125), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1760(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1761(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1762(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );

  xor2  gate1595(.a(N976), .b(N1040), .O(gate291inter0));
  nand2 gate1596(.a(gate291inter0), .b(s_102), .O(gate291inter1));
  and2  gate1597(.a(N976), .b(N1040), .O(gate291inter2));
  inv1  gate1598(.a(s_102), .O(gate291inter3));
  inv1  gate1599(.a(s_103), .O(gate291inter4));
  nand2 gate1600(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1601(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1602(.a(N1040), .O(gate291inter7));
  inv1  gate1603(.a(N976), .O(gate291inter8));
  nand2 gate1604(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1605(.a(s_103), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1606(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1607(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1608(.a(gate291inter12), .b(gate291inter1), .O(N1226));
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );

  xor2  gate895(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate896(.a(gate297inter0), .b(s_2), .O(gate297inter1));
  and2  gate897(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate898(.a(s_2), .O(gate297inter3));
  inv1  gate899(.a(s_3), .O(gate297inter4));
  nand2 gate900(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate901(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate902(.a(N1119), .O(gate297inter7));
  inv1  gate903(.a(N1120), .O(gate297inter8));
  nand2 gate904(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate905(.a(s_3), .b(gate297inter3), .O(gate297inter10));
  nor2  gate906(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate907(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate908(.a(gate297inter12), .b(gate297inter1), .O(N1232));

  xor2  gate993(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate994(.a(gate298inter0), .b(s_16), .O(gate298inter1));
  and2  gate995(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate996(.a(s_16), .O(gate298inter3));
  inv1  gate997(.a(s_17), .O(gate298inter4));
  nand2 gate998(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate999(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate1000(.a(N1121), .O(gate298inter7));
  inv1  gate1001(.a(N1122), .O(gate298inter8));
  nand2 gate1002(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate1003(.a(s_17), .b(gate298inter3), .O(gate298inter10));
  nor2  gate1004(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate1005(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate1006(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate2589(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate2590(.a(gate312inter0), .b(s_244), .O(gate312inter1));
  and2  gate2591(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate2592(.a(s_244), .O(gate312inter3));
  inv1  gate2593(.a(s_245), .O(gate312inter4));
  nand2 gate2594(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate2595(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate2596(.a(N631), .O(gate312inter7));
  inv1  gate2597(.a(N1159), .O(gate312inter8));
  nand2 gate2598(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate2599(.a(s_245), .b(gate312inter3), .O(gate312inter10));
  nor2  gate2600(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate2601(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate2602(.a(gate312inter12), .b(gate312inter1), .O(N1267));
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );

  xor2  gate1133(.a(N1223), .b(N709), .O(gate320inter0));
  nand2 gate1134(.a(gate320inter0), .b(s_36), .O(gate320inter1));
  and2  gate1135(.a(N1223), .b(N709), .O(gate320inter2));
  inv1  gate1136(.a(s_36), .O(gate320inter3));
  inv1  gate1137(.a(s_37), .O(gate320inter4));
  nand2 gate1138(.a(gate320inter4), .b(gate320inter3), .O(gate320inter5));
  nor2  gate1139(.a(gate320inter5), .b(gate320inter2), .O(gate320inter6));
  inv1  gate1140(.a(N709), .O(gate320inter7));
  inv1  gate1141(.a(N1223), .O(gate320inter8));
  nand2 gate1142(.a(gate320inter8), .b(gate320inter7), .O(gate320inter9));
  nand2 gate1143(.a(s_37), .b(gate320inter3), .O(gate320inter10));
  nor2  gate1144(.a(gate320inter10), .b(gate320inter9), .O(gate320inter11));
  nor2  gate1145(.a(gate320inter11), .b(gate320inter6), .O(gate320inter12));
  nand2 gate1146(.a(gate320inter12), .b(gate320inter1), .O(N1316));
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );

  xor2  gate2225(.a(N1238), .b(N730), .O(gate325inter0));
  nand2 gate2226(.a(gate325inter0), .b(s_192), .O(gate325inter1));
  and2  gate2227(.a(N1238), .b(N730), .O(gate325inter2));
  inv1  gate2228(.a(s_192), .O(gate325inter3));
  inv1  gate2229(.a(s_193), .O(gate325inter4));
  nand2 gate2230(.a(gate325inter4), .b(gate325inter3), .O(gate325inter5));
  nor2  gate2231(.a(gate325inter5), .b(gate325inter2), .O(gate325inter6));
  inv1  gate2232(.a(N730), .O(gate325inter7));
  inv1  gate2233(.a(N1238), .O(gate325inter8));
  nand2 gate2234(.a(gate325inter8), .b(gate325inter7), .O(gate325inter9));
  nand2 gate2235(.a(s_193), .b(gate325inter3), .O(gate325inter10));
  nor2  gate2236(.a(gate325inter10), .b(gate325inter9), .O(gate325inter11));
  nor2  gate2237(.a(gate325inter11), .b(gate325inter6), .O(gate325inter12));
  nand2 gate2238(.a(gate325inter12), .b(gate325inter1), .O(N1327));
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );

  xor2  gate2575(.a(N1210), .b(N1311), .O(gate337inter0));
  nand2 gate2576(.a(gate337inter0), .b(s_242), .O(gate337inter1));
  and2  gate2577(.a(N1210), .b(N1311), .O(gate337inter2));
  inv1  gate2578(.a(s_242), .O(gate337inter3));
  inv1  gate2579(.a(s_243), .O(gate337inter4));
  nand2 gate2580(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate2581(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate2582(.a(N1311), .O(gate337inter7));
  inv1  gate2583(.a(N1210), .O(gate337inter8));
  nand2 gate2584(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate2585(.a(s_243), .b(gate337inter3), .O(gate337inter10));
  nor2  gate2586(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate2587(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate2588(.a(gate337inter12), .b(gate337inter1), .O(N1358));

  xor2  gate2015(.a(N1212), .b(N1312), .O(gate338inter0));
  nand2 gate2016(.a(gate338inter0), .b(s_162), .O(gate338inter1));
  and2  gate2017(.a(N1212), .b(N1312), .O(gate338inter2));
  inv1  gate2018(.a(s_162), .O(gate338inter3));
  inv1  gate2019(.a(s_163), .O(gate338inter4));
  nand2 gate2020(.a(gate338inter4), .b(gate338inter3), .O(gate338inter5));
  nor2  gate2021(.a(gate338inter5), .b(gate338inter2), .O(gate338inter6));
  inv1  gate2022(.a(N1312), .O(gate338inter7));
  inv1  gate2023(.a(N1212), .O(gate338inter8));
  nand2 gate2024(.a(gate338inter8), .b(gate338inter7), .O(gate338inter9));
  nand2 gate2025(.a(s_163), .b(gate338inter3), .O(gate338inter10));
  nor2  gate2026(.a(gate338inter10), .b(gate338inter9), .O(gate338inter11));
  nor2  gate2027(.a(gate338inter11), .b(gate338inter6), .O(gate338inter12));
  nand2 gate2028(.a(gate338inter12), .b(gate338inter1), .O(N1361));
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );

  xor2  gate2645(.a(N1231), .b(N1322), .O(gate345inter0));
  nand2 gate2646(.a(gate345inter0), .b(s_252), .O(gate345inter1));
  and2  gate2647(.a(N1231), .b(N1322), .O(gate345inter2));
  inv1  gate2648(.a(s_252), .O(gate345inter3));
  inv1  gate2649(.a(s_253), .O(gate345inter4));
  nand2 gate2650(.a(gate345inter4), .b(gate345inter3), .O(gate345inter5));
  nor2  gate2651(.a(gate345inter5), .b(gate345inter2), .O(gate345inter6));
  inv1  gate2652(.a(N1322), .O(gate345inter7));
  inv1  gate2653(.a(N1231), .O(gate345inter8));
  nand2 gate2654(.a(gate345inter8), .b(gate345inter7), .O(gate345inter9));
  nand2 gate2655(.a(s_253), .b(gate345inter3), .O(gate345inter10));
  nor2  gate2656(.a(gate345inter10), .b(gate345inter9), .O(gate345inter11));
  nor2  gate2657(.a(gate345inter11), .b(gate345inter6), .O(gate345inter12));
  nand2 gate2658(.a(gate345inter12), .b(gate345inter1), .O(N1383));
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );

  xor2  gate1819(.a(N1007), .b(N1246), .O(gate355inter0));
  nand2 gate1820(.a(gate355inter0), .b(s_134), .O(gate355inter1));
  and2  gate1821(.a(N1007), .b(N1246), .O(gate355inter2));
  inv1  gate1822(.a(s_134), .O(gate355inter3));
  inv1  gate1823(.a(s_135), .O(gate355inter4));
  nand2 gate1824(.a(gate355inter4), .b(gate355inter3), .O(gate355inter5));
  nor2  gate1825(.a(gate355inter5), .b(gate355inter2), .O(gate355inter6));
  inv1  gate1826(.a(N1246), .O(gate355inter7));
  inv1  gate1827(.a(N1007), .O(gate355inter8));
  nand2 gate1828(.a(gate355inter8), .b(gate355inter7), .O(gate355inter9));
  nand2 gate1829(.a(s_135), .b(gate355inter3), .O(gate355inter10));
  nor2  gate1830(.a(gate355inter10), .b(gate355inter9), .O(gate355inter11));
  nor2  gate1831(.a(gate355inter11), .b(gate355inter6), .O(gate355inter12));
  nand2 gate1832(.a(gate355inter12), .b(gate355inter1), .O(N1399));
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );

  xor2  gate1063(.a(N1388), .b(N637), .O(gate362inter0));
  nand2 gate1064(.a(gate362inter0), .b(s_26), .O(gate362inter1));
  and2  gate1065(.a(N1388), .b(N637), .O(gate362inter2));
  inv1  gate1066(.a(s_26), .O(gate362inter3));
  inv1  gate1067(.a(s_27), .O(gate362inter4));
  nand2 gate1068(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate1069(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate1070(.a(N637), .O(gate362inter7));
  inv1  gate1071(.a(N1388), .O(gate362inter8));
  nand2 gate1072(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate1073(.a(s_27), .b(gate362inter3), .O(gate362inter10));
  nor2  gate1074(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate1075(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate1076(.a(gate362inter12), .b(gate362inter1), .O(N1434));
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );

  xor2  gate1413(.a(N1398), .b(N646), .O(gate364inter0));
  nand2 gate1414(.a(gate364inter0), .b(s_76), .O(gate364inter1));
  and2  gate1415(.a(N1398), .b(N646), .O(gate364inter2));
  inv1  gate1416(.a(s_76), .O(gate364inter3));
  inv1  gate1417(.a(s_77), .O(gate364inter4));
  nand2 gate1418(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate1419(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate1420(.a(N646), .O(gate364inter7));
  inv1  gate1421(.a(N1398), .O(gate364inter8));
  nand2 gate1422(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate1423(.a(s_77), .b(gate364inter3), .O(gate364inter10));
  nor2  gate1424(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate1425(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate1426(.a(gate364inter12), .b(gate364inter1), .O(N1439));
inv1 gate365( .a(N1344), .O(N1440) );

  xor2  gate2155(.a(N1148), .b(N1355), .O(gate366inter0));
  nand2 gate2156(.a(gate366inter0), .b(s_182), .O(gate366inter1));
  and2  gate2157(.a(N1148), .b(N1355), .O(gate366inter2));
  inv1  gate2158(.a(s_182), .O(gate366inter3));
  inv1  gate2159(.a(s_183), .O(gate366inter4));
  nand2 gate2160(.a(gate366inter4), .b(gate366inter3), .O(gate366inter5));
  nor2  gate2161(.a(gate366inter5), .b(gate366inter2), .O(gate366inter6));
  inv1  gate2162(.a(N1355), .O(gate366inter7));
  inv1  gate2163(.a(N1148), .O(gate366inter8));
  nand2 gate2164(.a(gate366inter8), .b(gate366inter7), .O(gate366inter9));
  nand2 gate2165(.a(s_183), .b(gate366inter3), .O(gate366inter10));
  nor2  gate2166(.a(gate366inter10), .b(gate366inter9), .O(gate366inter11));
  nor2  gate2167(.a(gate366inter11), .b(gate366inter6), .O(gate366inter12));
  nand2 gate2168(.a(gate366inter12), .b(gate366inter1), .O(N1443));
inv1 gate367( .a(N1355), .O(N1444) );

  xor2  gate1889(.a(N1149), .b(N1352), .O(gate368inter0));
  nand2 gate1890(.a(gate368inter0), .b(s_144), .O(gate368inter1));
  and2  gate1891(.a(N1149), .b(N1352), .O(gate368inter2));
  inv1  gate1892(.a(s_144), .O(gate368inter3));
  inv1  gate1893(.a(s_145), .O(gate368inter4));
  nand2 gate1894(.a(gate368inter4), .b(gate368inter3), .O(gate368inter5));
  nor2  gate1895(.a(gate368inter5), .b(gate368inter2), .O(gate368inter6));
  inv1  gate1896(.a(N1352), .O(gate368inter7));
  inv1  gate1897(.a(N1149), .O(gate368inter8));
  nand2 gate1898(.a(gate368inter8), .b(gate368inter7), .O(gate368inter9));
  nand2 gate1899(.a(s_145), .b(gate368inter3), .O(gate368inter10));
  nor2  gate1900(.a(gate368inter10), .b(gate368inter9), .O(gate368inter11));
  nor2  gate1901(.a(gate368inter11), .b(gate368inter6), .O(gate368inter12));
  nand2 gate1902(.a(gate368inter12), .b(gate368inter1), .O(N1445));
inv1 gate369( .a(N1352), .O(N1446) );

  xor2  gate1245(.a(N1151), .b(N1358), .O(gate370inter0));
  nand2 gate1246(.a(gate370inter0), .b(s_52), .O(gate370inter1));
  and2  gate1247(.a(N1151), .b(N1358), .O(gate370inter2));
  inv1  gate1248(.a(s_52), .O(gate370inter3));
  inv1  gate1249(.a(s_53), .O(gate370inter4));
  nand2 gate1250(.a(gate370inter4), .b(gate370inter3), .O(gate370inter5));
  nor2  gate1251(.a(gate370inter5), .b(gate370inter2), .O(gate370inter6));
  inv1  gate1252(.a(N1358), .O(gate370inter7));
  inv1  gate1253(.a(N1151), .O(gate370inter8));
  nand2 gate1254(.a(gate370inter8), .b(gate370inter7), .O(gate370inter9));
  nand2 gate1255(.a(s_53), .b(gate370inter3), .O(gate370inter10));
  nor2  gate1256(.a(gate370inter10), .b(gate370inter9), .O(gate370inter11));
  nor2  gate1257(.a(gate370inter11), .b(gate370inter6), .O(gate370inter12));
  nand2 gate1258(.a(gate370inter12), .b(gate370inter1), .O(N1447));
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );

  xor2  gate1259(.a(N1153), .b(N1367), .O(gate374inter0));
  nand2 gate1260(.a(gate374inter0), .b(s_54), .O(gate374inter1));
  and2  gate1261(.a(N1153), .b(N1367), .O(gate374inter2));
  inv1  gate1262(.a(s_54), .O(gate374inter3));
  inv1  gate1263(.a(s_55), .O(gate374inter4));
  nand2 gate1264(.a(gate374inter4), .b(gate374inter3), .O(gate374inter5));
  nor2  gate1265(.a(gate374inter5), .b(gate374inter2), .O(gate374inter6));
  inv1  gate1266(.a(N1367), .O(gate374inter7));
  inv1  gate1267(.a(N1153), .O(gate374inter8));
  nand2 gate1268(.a(gate374inter8), .b(gate374inter7), .O(gate374inter9));
  nand2 gate1269(.a(s_55), .b(gate374inter3), .O(gate374inter10));
  nor2  gate1270(.a(gate374inter10), .b(gate374inter9), .O(gate374inter11));
  nor2  gate1271(.a(gate374inter11), .b(gate374inter6), .O(gate374inter12));
  nand2 gate1272(.a(gate374inter12), .b(gate374inter1), .O(N1453));
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate1987(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate1988(.a(gate376inter0), .b(s_158), .O(gate376inter1));
  and2  gate1989(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate1990(.a(s_158), .O(gate376inter3));
  inv1  gate1991(.a(s_159), .O(gate376inter4));
  nand2 gate1992(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate1993(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate1994(.a(N1364), .O(gate376inter7));
  inv1  gate1995(.a(N1154), .O(gate376inter8));
  nand2 gate1996(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate1997(.a(s_159), .b(gate376inter3), .O(gate376inter10));
  nor2  gate1998(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate1999(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate2000(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate2673(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate2674(.a(gate383inter0), .b(s_256), .O(gate383inter1));
  and2  gate2675(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate2676(.a(s_256), .O(gate383inter3));
  inv1  gate2677(.a(s_257), .O(gate383inter4));
  nand2 gate2678(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate2679(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate2680(.a(N1393), .O(gate383inter7));
  inv1  gate2681(.a(N1161), .O(gate383inter8));
  nand2 gate2682(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate2683(.a(s_257), .b(gate383inter3), .O(gate383inter10));
  nor2  gate2684(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate2685(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate2686(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );

  xor2  gate1707(.a(N1222), .b(N1370), .O(gate387inter0));
  nand2 gate1708(.a(gate387inter0), .b(s_118), .O(gate387inter1));
  and2  gate1709(.a(N1222), .b(N1370), .O(gate387inter2));
  inv1  gate1710(.a(s_118), .O(gate387inter3));
  inv1  gate1711(.a(s_119), .O(gate387inter4));
  nand2 gate1712(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1713(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1714(.a(N1370), .O(gate387inter7));
  inv1  gate1715(.a(N1222), .O(gate387inter8));
  nand2 gate1716(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1717(.a(s_119), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1718(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1719(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1720(.a(gate387inter12), .b(gate387inter1), .O(N1469));
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );

  xor2  gate2099(.a(N1433), .b(N1387), .O(gate390inter0));
  nand2 gate2100(.a(gate390inter0), .b(s_174), .O(gate390inter1));
  and2  gate2101(.a(N1433), .b(N1387), .O(gate390inter2));
  inv1  gate2102(.a(s_174), .O(gate390inter3));
  inv1  gate2103(.a(s_175), .O(gate390inter4));
  nand2 gate2104(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2105(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2106(.a(N1387), .O(gate390inter7));
  inv1  gate2107(.a(N1433), .O(gate390inter8));
  nand2 gate2108(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2109(.a(s_175), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2110(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2111(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2112(.a(gate390inter12), .b(gate390inter1), .O(N1472));
inv1 gate391( .a(N1390), .O(N1475) );

  xor2  gate1847(.a(N1240), .b(N1390), .O(gate392inter0));
  nand2 gate1848(.a(gate392inter0), .b(s_138), .O(gate392inter1));
  and2  gate1849(.a(N1240), .b(N1390), .O(gate392inter2));
  inv1  gate1850(.a(s_138), .O(gate392inter3));
  inv1  gate1851(.a(s_139), .O(gate392inter4));
  nand2 gate1852(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1853(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1854(.a(N1390), .O(gate392inter7));
  inv1  gate1855(.a(N1240), .O(gate392inter8));
  nand2 gate1856(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1857(.a(s_139), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1858(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1859(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1860(.a(gate392inter12), .b(gate392inter1), .O(N1476));

  xor2  gate2547(.a(N1434), .b(N1389), .O(gate393inter0));
  nand2 gate2548(.a(gate393inter0), .b(s_238), .O(gate393inter1));
  and2  gate2549(.a(N1434), .b(N1389), .O(gate393inter2));
  inv1  gate2550(.a(s_238), .O(gate393inter3));
  inv1  gate2551(.a(s_239), .O(gate393inter4));
  nand2 gate2552(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2553(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2554(.a(N1389), .O(gate393inter7));
  inv1  gate2555(.a(N1434), .O(gate393inter8));
  nand2 gate2556(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2557(.a(s_239), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2558(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2559(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2560(.a(gate393inter12), .b(gate393inter1), .O(N1478));
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );

  xor2  gate2379(.a(N1444), .b(N939), .O(gate396inter0));
  nand2 gate2380(.a(gate396inter0), .b(s_214), .O(gate396inter1));
  and2  gate2381(.a(N1444), .b(N939), .O(gate396inter2));
  inv1  gate2382(.a(s_214), .O(gate396inter3));
  inv1  gate2383(.a(s_215), .O(gate396inter4));
  nand2 gate2384(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2385(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2386(.a(N939), .O(gate396inter7));
  inv1  gate2387(.a(N1444), .O(gate396inter8));
  nand2 gate2388(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2389(.a(s_215), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2390(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2391(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2392(.a(gate396inter12), .b(gate396inter1), .O(N1487));
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );

  xor2  gate1091(.a(N1448), .b(N943), .O(gate398inter0));
  nand2 gate1092(.a(gate398inter0), .b(s_30), .O(gate398inter1));
  and2  gate1093(.a(N1448), .b(N943), .O(gate398inter2));
  inv1  gate1094(.a(s_30), .O(gate398inter3));
  inv1  gate1095(.a(s_31), .O(gate398inter4));
  nand2 gate1096(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1097(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1098(.a(N943), .O(gate398inter7));
  inv1  gate1099(.a(N1448), .O(gate398inter8));
  nand2 gate1100(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1101(.a(s_31), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1102(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1103(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1104(.a(gate398inter12), .b(gate398inter1), .O(N1489));
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );

  xor2  gate1623(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate1624(.a(gate402inter0), .b(s_106), .O(gate402inter1));
  and2  gate1625(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate1626(.a(s_106), .O(gate402inter3));
  inv1  gate1627(.a(s_107), .O(gate402inter4));
  nand2 gate1628(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1629(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1630(.a(N955), .O(gate402inter7));
  inv1  gate1631(.a(N1454), .O(gate402inter8));
  nand2 gate1632(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1633(.a(s_107), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1634(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1635(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1636(.a(gate402inter12), .b(gate402inter1), .O(N1493));

  xor2  gate2183(.a(N1456), .b(N951), .O(gate403inter0));
  nand2 gate2184(.a(gate403inter0), .b(s_186), .O(gate403inter1));
  and2  gate2185(.a(N1456), .b(N951), .O(gate403inter2));
  inv1  gate2186(.a(s_186), .O(gate403inter3));
  inv1  gate2187(.a(s_187), .O(gate403inter4));
  nand2 gate2188(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2189(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2190(.a(N951), .O(gate403inter7));
  inv1  gate2191(.a(N1456), .O(gate403inter8));
  nand2 gate2192(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2193(.a(s_187), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2194(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2195(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2196(.a(gate403inter12), .b(gate403inter1), .O(N1494));

  xor2  gate951(.a(N1458), .b(N969), .O(gate404inter0));
  nand2 gate952(.a(gate404inter0), .b(s_10), .O(gate404inter1));
  and2  gate953(.a(N1458), .b(N969), .O(gate404inter2));
  inv1  gate954(.a(s_10), .O(gate404inter3));
  inv1  gate955(.a(s_11), .O(gate404inter4));
  nand2 gate956(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate957(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate958(.a(N969), .O(gate404inter7));
  inv1  gate959(.a(N1458), .O(gate404inter8));
  nand2 gate960(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate961(.a(s_11), .b(gate404inter3), .O(gate404inter10));
  nor2  gate962(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate963(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate964(.a(gate404inter12), .b(gate404inter1), .O(N1495));

  xor2  gate2603(.a(N1460), .b(N977), .O(gate405inter0));
  nand2 gate2604(.a(gate405inter0), .b(s_246), .O(gate405inter1));
  and2  gate2605(.a(N1460), .b(N977), .O(gate405inter2));
  inv1  gate2606(.a(s_246), .O(gate405inter3));
  inv1  gate2607(.a(s_247), .O(gate405inter4));
  nand2 gate2608(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2609(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2610(.a(N977), .O(gate405inter7));
  inv1  gate2611(.a(N1460), .O(gate405inter8));
  nand2 gate2612(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2613(.a(s_247), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2614(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2615(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2616(.a(gate405inter12), .b(gate405inter1), .O(N1496));

  xor2  gate2085(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate2086(.a(gate406inter0), .b(s_172), .O(gate406inter1));
  and2  gate2087(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate2088(.a(s_172), .O(gate406inter3));
  inv1  gate2089(.a(s_173), .O(gate406inter4));
  nand2 gate2090(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2091(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2092(.a(N998), .O(gate406inter7));
  inv1  gate2093(.a(N1463), .O(gate406inter8));
  nand2 gate2094(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2095(.a(s_173), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2096(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2097(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2098(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );

  xor2  gate1147(.a(N1468), .b(N965), .O(gate408inter0));
  nand2 gate1148(.a(gate408inter0), .b(s_38), .O(gate408inter1));
  and2  gate1149(.a(N1468), .b(N965), .O(gate408inter2));
  inv1  gate1150(.a(s_38), .O(gate408inter3));
  inv1  gate1151(.a(s_39), .O(gate408inter4));
  nand2 gate1152(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1153(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1154(.a(N965), .O(gate408inter7));
  inv1  gate1155(.a(N1468), .O(gate408inter8));
  nand2 gate1156(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1157(.a(s_39), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1158(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1159(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1160(.a(gate408inter12), .b(gate408inter1), .O(N1500));

  xor2  gate2435(.a(N1470), .b(N973), .O(gate409inter0));
  nand2 gate2436(.a(gate409inter0), .b(s_222), .O(gate409inter1));
  and2  gate2437(.a(N1470), .b(N973), .O(gate409inter2));
  inv1  gate2438(.a(s_222), .O(gate409inter3));
  inv1  gate2439(.a(s_223), .O(gate409inter4));
  nand2 gate2440(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2441(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2442(.a(N973), .O(gate409inter7));
  inv1  gate2443(.a(N1470), .O(gate409inter8));
  nand2 gate2444(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2445(.a(s_223), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2446(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2447(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2448(.a(gate409inter12), .b(gate409inter1), .O(N1501));

  xor2  gate1315(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate1316(.a(gate410inter0), .b(s_62), .O(gate410inter1));
  and2  gate1317(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate1318(.a(s_62), .O(gate410inter3));
  inv1  gate1319(.a(s_63), .O(gate410inter4));
  nand2 gate1320(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1321(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1322(.a(N994), .O(gate410inter7));
  inv1  gate1323(.a(N1475), .O(gate410inter8));
  nand2 gate1324(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1325(.a(s_63), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1326(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1327(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1328(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );

  xor2  gate2309(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate2310(.a(gate413inter0), .b(s_204), .O(gate413inter1));
  and2  gate2311(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate2312(.a(s_204), .O(gate413inter3));
  inv1  gate2313(.a(s_205), .O(gate413inter4));
  nand2 gate2314(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2315(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2316(.a(N1445), .O(gate413inter7));
  inv1  gate2317(.a(N1488), .O(gate413inter8));
  nand2 gate2318(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2319(.a(s_205), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2320(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2321(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2322(.a(gate413inter12), .b(gate413inter1), .O(N1514));

  xor2  gate1469(.a(N1489), .b(N1447), .O(gate414inter0));
  nand2 gate1470(.a(gate414inter0), .b(s_84), .O(gate414inter1));
  and2  gate1471(.a(N1489), .b(N1447), .O(gate414inter2));
  inv1  gate1472(.a(s_84), .O(gate414inter3));
  inv1  gate1473(.a(s_85), .O(gate414inter4));
  nand2 gate1474(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1475(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1476(.a(N1447), .O(gate414inter7));
  inv1  gate1477(.a(N1489), .O(gate414inter8));
  nand2 gate1478(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1479(.a(s_85), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1480(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1481(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1482(.a(gate414inter12), .b(gate414inter1), .O(N1517));

  xor2  gate1021(.a(N1492), .b(N1451), .O(gate415inter0));
  nand2 gate1022(.a(gate415inter0), .b(s_20), .O(gate415inter1));
  and2  gate1023(.a(N1492), .b(N1451), .O(gate415inter2));
  inv1  gate1024(.a(s_20), .O(gate415inter3));
  inv1  gate1025(.a(s_21), .O(gate415inter4));
  nand2 gate1026(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1027(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1028(.a(N1451), .O(gate415inter7));
  inv1  gate1029(.a(N1492), .O(gate415inter8));
  nand2 gate1030(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1031(.a(s_21), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1032(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1033(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1034(.a(gate415inter12), .b(gate415inter1), .O(N1520));
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );

  xor2  gate2617(.a(N1494), .b(N1455), .O(gate417inter0));
  nand2 gate2618(.a(gate417inter0), .b(s_248), .O(gate417inter1));
  and2  gate2619(.a(N1494), .b(N1455), .O(gate417inter2));
  inv1  gate2620(.a(s_248), .O(gate417inter3));
  inv1  gate2621(.a(s_249), .O(gate417inter4));
  nand2 gate2622(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2623(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2624(.a(N1455), .O(gate417inter7));
  inv1  gate2625(.a(N1494), .O(gate417inter8));
  nand2 gate2626(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2627(.a(s_249), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2628(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2629(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2630(.a(gate417inter12), .b(gate417inter1), .O(N1522));
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );

  xor2  gate1651(.a(N1496), .b(N1459), .O(gate419inter0));
  nand2 gate1652(.a(gate419inter0), .b(s_110), .O(gate419inter1));
  and2  gate1653(.a(N1496), .b(N1459), .O(gate419inter2));
  inv1  gate1654(.a(s_110), .O(gate419inter3));
  inv1  gate1655(.a(s_111), .O(gate419inter4));
  nand2 gate1656(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1657(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1658(.a(N1459), .O(gate419inter7));
  inv1  gate1659(.a(N1496), .O(gate419inter8));
  nand2 gate1660(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1661(.a(s_111), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1662(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1663(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1664(.a(gate419inter12), .b(gate419inter1), .O(N1527));
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );

  xor2  gate2393(.a(N1501), .b(N1471), .O(gate425inter0));
  nand2 gate2394(.a(gate425inter0), .b(s_216), .O(gate425inter1));
  and2  gate2395(.a(N1501), .b(N1471), .O(gate425inter2));
  inv1  gate2396(.a(s_216), .O(gate425inter3));
  inv1  gate2397(.a(s_217), .O(gate425inter4));
  nand2 gate2398(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2399(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2400(.a(N1471), .O(gate425inter7));
  inv1  gate2401(.a(N1501), .O(gate425inter8));
  nand2 gate2402(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2403(.a(s_217), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2404(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2405(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2406(.a(gate425inter12), .b(gate425inter1), .O(N1534));
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );

  xor2  gate1735(.a(N1531), .b(N1484), .O(gate432inter0));
  nand2 gate1736(.a(gate432inter0), .b(s_122), .O(gate432inter1));
  and2  gate1737(.a(N1531), .b(N1484), .O(gate432inter2));
  inv1  gate1738(.a(s_122), .O(gate432inter3));
  inv1  gate1739(.a(s_123), .O(gate432inter4));
  nand2 gate1740(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1741(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1742(.a(N1484), .O(gate432inter7));
  inv1  gate1743(.a(N1531), .O(gate432inter8));
  nand2 gate1744(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1745(.a(s_123), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1746(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1747(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1748(.a(gate432inter12), .b(gate432inter1), .O(N1567));
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );

  xor2  gate2687(.a(N1569), .b(N1576), .O(gate453inter0));
  nand2 gate2688(.a(gate453inter0), .b(s_258), .O(gate453inter1));
  and2  gate2689(.a(N1569), .b(N1576), .O(gate453inter2));
  inv1  gate2690(.a(s_258), .O(gate453inter3));
  inv1  gate2691(.a(s_259), .O(gate453inter4));
  nand2 gate2692(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2693(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2694(.a(N1576), .O(gate453inter7));
  inv1  gate2695(.a(N1569), .O(gate453inter8));
  nand2 gate2696(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2697(.a(s_259), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2698(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2699(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2700(.a(gate453inter12), .b(gate453inter1), .O(N1638));
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );

  xor2  gate2211(.a(N1217), .b(N1606), .O(gate466inter0));
  nand2 gate2212(.a(gate466inter0), .b(s_190), .O(gate466inter1));
  and2  gate2213(.a(N1217), .b(N1606), .O(gate466inter2));
  inv1  gate2214(.a(s_190), .O(gate466inter3));
  inv1  gate2215(.a(s_191), .O(gate466inter4));
  nand2 gate2216(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2217(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2218(.a(N1606), .O(gate466inter7));
  inv1  gate2219(.a(N1217), .O(gate466inter8));
  nand2 gate2220(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2221(.a(s_191), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2222(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2223(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2224(.a(gate466inter12), .b(gate466inter1), .O(N1678));
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );

  xor2  gate2477(.a(N1636), .b(N1594), .O(gate472inter0));
  nand2 gate2478(.a(gate472inter0), .b(s_228), .O(gate472inter1));
  and2  gate2479(.a(N1636), .b(N1594), .O(gate472inter2));
  inv1  gate2480(.a(s_228), .O(gate472inter3));
  inv1  gate2481(.a(s_229), .O(gate472inter4));
  nand2 gate2482(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2483(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2484(.a(N1594), .O(gate472inter7));
  inv1  gate2485(.a(N1636), .O(gate472inter8));
  nand2 gate2486(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2487(.a(s_229), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2488(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2489(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2490(.a(gate472inter12), .b(gate472inter1), .O(N1685));
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );

  xor2  gate2001(.a(N1679), .b(N1028), .O(gate482inter0));
  nand2 gate2002(.a(gate482inter0), .b(s_160), .O(gate482inter1));
  and2  gate2003(.a(N1679), .b(N1028), .O(gate482inter2));
  inv1  gate2004(.a(s_160), .O(gate482inter3));
  inv1  gate2005(.a(s_161), .O(gate482inter4));
  nand2 gate2006(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2007(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2008(.a(N1028), .O(gate482inter7));
  inv1  gate2009(.a(N1679), .O(gate482inter8));
  nand2 gate2010(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2011(.a(s_161), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2012(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2013(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2014(.a(gate482inter12), .b(gate482inter1), .O(N1712));

  xor2  gate1035(.a(N1681), .b(N1031), .O(gate483inter0));
  nand2 gate1036(.a(gate483inter0), .b(s_22), .O(gate483inter1));
  and2  gate1037(.a(N1681), .b(N1031), .O(gate483inter2));
  inv1  gate1038(.a(s_22), .O(gate483inter3));
  inv1  gate1039(.a(s_23), .O(gate483inter4));
  nand2 gate1040(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1041(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1042(.a(N1031), .O(gate483inter7));
  inv1  gate1043(.a(N1681), .O(gate483inter8));
  nand2 gate1044(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1045(.a(s_23), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1046(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1047(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1048(.a(gate483inter12), .b(gate483inter1), .O(N1713));
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );

  xor2  gate1805(.a(N1593), .b(N1658), .O(gate486inter0));
  nand2 gate1806(.a(gate486inter0), .b(s_132), .O(gate486inter1));
  and2  gate1807(.a(N1593), .b(N1658), .O(gate486inter2));
  inv1  gate1808(.a(s_132), .O(gate486inter3));
  inv1  gate1809(.a(s_133), .O(gate486inter4));
  nand2 gate1810(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1811(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1812(.a(N1658), .O(gate486inter7));
  inv1  gate1813(.a(N1593), .O(gate486inter8));
  nand2 gate1814(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1815(.a(s_133), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1816(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1817(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1818(.a(gate486inter12), .b(gate486inter1), .O(N1720));
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );

  xor2  gate1763(.a(N1711), .b(N1603), .O(gate498inter0));
  nand2 gate1764(.a(gate498inter0), .b(s_126), .O(gate498inter1));
  and2  gate1765(.a(N1711), .b(N1603), .O(gate498inter2));
  inv1  gate1766(.a(s_126), .O(gate498inter3));
  inv1  gate1767(.a(s_127), .O(gate498inter4));
  nand2 gate1768(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1769(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1770(.a(N1603), .O(gate498inter7));
  inv1  gate1771(.a(N1711), .O(gate498inter8));
  nand2 gate1772(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1773(.a(s_127), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1774(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1775(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1776(.a(gate498inter12), .b(gate498inter1), .O(N1747));
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );

  xor2  gate1721(.a(N1721), .b(N1537), .O(gate501inter0));
  nand2 gate1722(.a(gate501inter0), .b(s_120), .O(gate501inter1));
  and2  gate1723(.a(N1721), .b(N1537), .O(gate501inter2));
  inv1  gate1724(.a(s_120), .O(gate501inter3));
  inv1  gate1725(.a(s_121), .O(gate501inter4));
  nand2 gate1726(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1727(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1728(.a(N1537), .O(gate501inter7));
  inv1  gate1729(.a(N1721), .O(gate501inter8));
  nand2 gate1730(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1731(.a(s_121), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1732(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1733(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1734(.a(gate501inter12), .b(gate501inter1), .O(N1759));
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );

  xor2  gate1973(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate1974(.a(gate508inter0), .b(s_156), .O(gate508inter1));
  and2  gate1975(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate1976(.a(s_156), .O(gate508inter3));
  inv1  gate1977(.a(s_157), .O(gate508inter4));
  nand2 gate1978(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1979(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1980(.a(N1723), .O(gate508inter7));
  inv1  gate1981(.a(N1413), .O(gate508inter8));
  nand2 gate1982(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1983(.a(s_157), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1984(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1985(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1986(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );

  xor2  gate1399(.a(N1747), .b(N1710), .O(gate511inter0));
  nand2 gate1400(.a(gate511inter0), .b(s_74), .O(gate511inter1));
  and2  gate1401(.a(N1747), .b(N1710), .O(gate511inter2));
  inv1  gate1402(.a(s_74), .O(gate511inter3));
  inv1  gate1403(.a(s_75), .O(gate511inter4));
  nand2 gate1404(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1405(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1406(.a(N1710), .O(gate511inter7));
  inv1  gate1407(.a(N1747), .O(gate511inter8));
  nand2 gate1408(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1409(.a(s_75), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1410(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1411(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1412(.a(gate511inter12), .b(gate511inter1), .O(N1777));
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1861(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1862(.a(gate513inter0), .b(s_140), .O(gate513inter1));
  and2  gate1863(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1864(.a(s_140), .O(gate513inter3));
  inv1  gate1865(.a(s_141), .O(gate513inter4));
  nand2 gate1866(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1867(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1868(.a(N1731), .O(gate513inter7));
  inv1  gate1869(.a(N1682), .O(gate513inter8));
  nand2 gate1870(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1871(.a(s_141), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1872(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1873(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1874(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );

  xor2  gate1875(.a(N1683), .b(N1734), .O(gate516inter0));
  nand2 gate1876(.a(gate516inter0), .b(s_142), .O(gate516inter1));
  and2  gate1877(.a(N1683), .b(N1734), .O(gate516inter2));
  inv1  gate1878(.a(s_142), .O(gate516inter3));
  inv1  gate1879(.a(s_143), .O(gate516inter4));
  nand2 gate1880(.a(gate516inter4), .b(gate516inter3), .O(gate516inter5));
  nor2  gate1881(.a(gate516inter5), .b(gate516inter2), .O(gate516inter6));
  inv1  gate1882(.a(N1734), .O(gate516inter7));
  inv1  gate1883(.a(N1683), .O(gate516inter8));
  nand2 gate1884(.a(gate516inter8), .b(gate516inter7), .O(gate516inter9));
  nand2 gate1885(.a(s_143), .b(gate516inter3), .O(gate516inter10));
  nor2  gate1886(.a(gate516inter10), .b(gate516inter9), .O(gate516inter11));
  nor2  gate1887(.a(gate516inter11), .b(gate516inter6), .O(gate516inter12));
  nand2 gate1888(.a(gate516inter12), .b(gate516inter1), .O(N1787));
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );

  xor2  gate1343(.a(N1773), .b(N1334), .O(gate523inter0));
  nand2 gate1344(.a(gate523inter0), .b(s_66), .O(gate523inter1));
  and2  gate1345(.a(N1773), .b(N1334), .O(gate523inter2));
  inv1  gate1346(.a(s_66), .O(gate523inter3));
  inv1  gate1347(.a(s_67), .O(gate523inter4));
  nand2 gate1348(.a(gate523inter4), .b(gate523inter3), .O(gate523inter5));
  nor2  gate1349(.a(gate523inter5), .b(gate523inter2), .O(gate523inter6));
  inv1  gate1350(.a(N1334), .O(gate523inter7));
  inv1  gate1351(.a(N1773), .O(gate523inter8));
  nand2 gate1352(.a(gate523inter8), .b(gate523inter7), .O(gate523inter9));
  nand2 gate1353(.a(s_67), .b(gate523inter3), .O(gate523inter10));
  nor2  gate1354(.a(gate523inter10), .b(gate523inter9), .O(gate523inter11));
  nor2  gate1355(.a(gate523inter11), .b(gate523inter6), .O(gate523inter12));
  nand2 gate1356(.a(gate523inter12), .b(gate523inter1), .O(N1801));
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );

  xor2  gate1217(.a(N1783), .b(N1612), .O(gate527inter0));
  nand2 gate1218(.a(gate527inter0), .b(s_48), .O(gate527inter1));
  and2  gate1219(.a(N1783), .b(N1612), .O(gate527inter2));
  inv1  gate1220(.a(s_48), .O(gate527inter3));
  inv1  gate1221(.a(s_49), .O(gate527inter4));
  nand2 gate1222(.a(gate527inter4), .b(gate527inter3), .O(gate527inter5));
  nor2  gate1223(.a(gate527inter5), .b(gate527inter2), .O(gate527inter6));
  inv1  gate1224(.a(N1612), .O(gate527inter7));
  inv1  gate1225(.a(N1783), .O(gate527inter8));
  nand2 gate1226(.a(gate527inter8), .b(gate527inter7), .O(gate527inter9));
  nand2 gate1227(.a(s_49), .b(gate527inter3), .O(gate527inter10));
  nor2  gate1228(.a(gate527inter10), .b(gate527inter9), .O(gate527inter11));
  nor2  gate1229(.a(gate527inter11), .b(gate527inter6), .O(gate527inter12));
  nand2 gate1230(.a(gate527inter12), .b(gate527inter1), .O(N1809));

  xor2  gate2253(.a(N1786), .b(N1615), .O(gate528inter0));
  nand2 gate2254(.a(gate528inter0), .b(s_196), .O(gate528inter1));
  and2  gate2255(.a(N1786), .b(N1615), .O(gate528inter2));
  inv1  gate2256(.a(s_196), .O(gate528inter3));
  inv1  gate2257(.a(s_197), .O(gate528inter4));
  nand2 gate2258(.a(gate528inter4), .b(gate528inter3), .O(gate528inter5));
  nor2  gate2259(.a(gate528inter5), .b(gate528inter2), .O(gate528inter6));
  inv1  gate2260(.a(N1615), .O(gate528inter7));
  inv1  gate2261(.a(N1786), .O(gate528inter8));
  nand2 gate2262(.a(gate528inter8), .b(gate528inter7), .O(gate528inter9));
  nand2 gate2263(.a(s_197), .b(gate528inter3), .O(gate528inter10));
  nor2  gate2264(.a(gate528inter10), .b(gate528inter9), .O(gate528inter11));
  nor2  gate2265(.a(gate528inter11), .b(gate528inter6), .O(gate528inter12));
  nand2 gate2266(.a(gate528inter12), .b(gate528inter1), .O(N1810));

  xor2  gate1301(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate1302(.a(gate529inter0), .b(s_60), .O(gate529inter1));
  and2  gate1303(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate1304(.a(s_60), .O(gate529inter3));
  inv1  gate1305(.a(s_61), .O(gate529inter4));
  nand2 gate1306(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate1307(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate1308(.a(N1791), .O(gate529inter7));
  inv1  gate1309(.a(N1762), .O(gate529inter8));
  nand2 gate1310(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate1311(.a(s_61), .b(gate529inter3), .O(gate529inter10));
  nor2  gate1312(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate1313(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate1314(.a(gate529inter12), .b(gate529inter1), .O(N1812));
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );

  xor2  gate1455(.a(N1801), .b(N1772), .O(gate539inter0));
  nand2 gate1456(.a(gate539inter0), .b(s_82), .O(gate539inter1));
  and2  gate1457(.a(N1801), .b(N1772), .O(gate539inter2));
  inv1  gate1458(.a(s_82), .O(gate539inter3));
  inv1  gate1459(.a(s_83), .O(gate539inter4));
  nand2 gate1460(.a(gate539inter4), .b(gate539inter3), .O(gate539inter5));
  nor2  gate1461(.a(gate539inter5), .b(gate539inter2), .O(gate539inter6));
  inv1  gate1462(.a(N1772), .O(gate539inter7));
  inv1  gate1463(.a(N1801), .O(gate539inter8));
  nand2 gate1464(.a(gate539inter8), .b(gate539inter7), .O(gate539inter9));
  nand2 gate1465(.a(s_83), .b(gate539inter3), .O(gate539inter10));
  nor2  gate1466(.a(gate539inter10), .b(gate539inter9), .O(gate539inter11));
  nor2  gate1467(.a(gate539inter11), .b(gate539inter6), .O(gate539inter12));
  nand2 gate1468(.a(gate539inter12), .b(gate539inter1), .O(N1830));
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );

  xor2  gate1777(.a(N1822), .b(N1419), .O(gate543inter0));
  nand2 gate1778(.a(gate543inter0), .b(s_128), .O(gate543inter1));
  and2  gate1779(.a(N1822), .b(N1419), .O(gate543inter2));
  inv1  gate1780(.a(s_128), .O(gate543inter3));
  inv1  gate1781(.a(s_129), .O(gate543inter4));
  nand2 gate1782(.a(gate543inter4), .b(gate543inter3), .O(gate543inter5));
  nor2  gate1783(.a(gate543inter5), .b(gate543inter2), .O(gate543inter6));
  inv1  gate1784(.a(N1419), .O(gate543inter7));
  inv1  gate1785(.a(N1822), .O(gate543inter8));
  nand2 gate1786(.a(gate543inter8), .b(gate543inter7), .O(gate543inter9));
  nand2 gate1787(.a(s_129), .b(gate543inter3), .O(gate543inter10));
  nor2  gate1788(.a(gate543inter10), .b(gate543inter9), .O(gate543inter11));
  nor2  gate1789(.a(gate543inter11), .b(gate543inter6), .O(gate543inter12));
  nand2 gate1790(.a(gate543inter12), .b(gate543inter1), .O(N1848));
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );

  xor2  gate1581(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate1582(.a(gate546inter0), .b(s_100), .O(gate546inter1));
  and2  gate1583(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate1584(.a(s_100), .O(gate546inter3));
  inv1  gate1585(.a(s_101), .O(gate546inter4));
  nand2 gate1586(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate1587(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate1588(.a(N1319), .O(gate546inter7));
  inv1  gate1589(.a(N1827), .O(gate546inter8));
  nand2 gate1590(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate1591(.a(s_101), .b(gate546inter3), .O(gate546inter10));
  nor2  gate1592(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate1593(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate1594(.a(gate546inter12), .b(gate546inter1), .O(N1852));
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );

  xor2  gate1567(.a(N1848), .b(N1821), .O(gate557inter0));
  nand2 gate1568(.a(gate557inter0), .b(s_98), .O(gate557inter1));
  and2  gate1569(.a(N1848), .b(N1821), .O(gate557inter2));
  inv1  gate1570(.a(s_98), .O(gate557inter3));
  inv1  gate1571(.a(s_99), .O(gate557inter4));
  nand2 gate1572(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate1573(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate1574(.a(N1821), .O(gate557inter7));
  inv1  gate1575(.a(N1848), .O(gate557inter8));
  nand2 gate1576(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate1577(.a(s_99), .b(gate557inter3), .O(gate557inter10));
  nor2  gate1578(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate1579(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate1580(.a(gate557inter12), .b(gate557inter1), .O(N1878));

  xor2  gate2057(.a(N1849), .b(N1823), .O(gate558inter0));
  nand2 gate2058(.a(gate558inter0), .b(s_168), .O(gate558inter1));
  and2  gate2059(.a(N1849), .b(N1823), .O(gate558inter2));
  inv1  gate2060(.a(s_168), .O(gate558inter3));
  inv1  gate2061(.a(s_169), .O(gate558inter4));
  nand2 gate2062(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate2063(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate2064(.a(N1823), .O(gate558inter7));
  inv1  gate2065(.a(N1849), .O(gate558inter8));
  nand2 gate2066(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate2067(.a(s_169), .b(gate558inter3), .O(gate558inter10));
  nor2  gate2068(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate2069(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate2070(.a(gate558inter12), .b(gate558inter1), .O(N1879));
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );

  xor2  gate2701(.a(N1852), .b(N1826), .O(gate561inter0));
  nand2 gate2702(.a(gate561inter0), .b(s_260), .O(gate561inter1));
  and2  gate2703(.a(N1852), .b(N1826), .O(gate561inter2));
  inv1  gate2704(.a(s_260), .O(gate561inter3));
  inv1  gate2705(.a(s_261), .O(gate561inter4));
  nand2 gate2706(.a(gate561inter4), .b(gate561inter3), .O(gate561inter5));
  nor2  gate2707(.a(gate561inter5), .b(gate561inter2), .O(gate561inter6));
  inv1  gate2708(.a(N1826), .O(gate561inter7));
  inv1  gate2709(.a(N1852), .O(gate561inter8));
  nand2 gate2710(.a(gate561inter8), .b(gate561inter7), .O(gate561inter9));
  nand2 gate2711(.a(s_261), .b(gate561inter3), .O(gate561inter10));
  nor2  gate2712(.a(gate561inter10), .b(gate561inter9), .O(gate561inter11));
  nor2  gate2713(.a(gate561inter11), .b(gate561inter6), .O(gate561inter12));
  nand2 gate2714(.a(gate561inter12), .b(gate561inter1), .O(N1884));
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );

  xor2  gate2323(.a(N1864), .b(N1640), .O(gate566inter0));
  nand2 gate2324(.a(gate566inter0), .b(s_206), .O(gate566inter1));
  and2  gate2325(.a(N1864), .b(N1640), .O(gate566inter2));
  inv1  gate2326(.a(s_206), .O(gate566inter3));
  inv1  gate2327(.a(s_207), .O(gate566inter4));
  nand2 gate2328(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate2329(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate2330(.a(N1640), .O(gate566inter7));
  inv1  gate2331(.a(N1864), .O(gate566inter8));
  nand2 gate2332(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate2333(.a(s_207), .b(gate566inter3), .O(gate566inter10));
  nor2  gate2334(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate2335(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate2336(.a(gate566inter12), .b(gate566inter1), .O(N1897));
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate1049(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate1050(.a(gate579inter0), .b(s_24), .O(gate579inter1));
  and2  gate1051(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate1052(.a(s_24), .O(gate579inter3));
  inv1  gate1053(.a(s_25), .O(gate579inter4));
  nand2 gate1054(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate1055(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate1056(.a(N1714), .O(gate579inter7));
  inv1  gate1057(.a(N1895), .O(gate579inter8));
  nand2 gate1058(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate1059(.a(s_25), .b(gate579inter3), .O(gate579inter10));
  nor2  gate1060(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate1061(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate1062(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );

  xor2  gate1077(.a(N1924), .b(N1896), .O(gate593inter0));
  nand2 gate1078(.a(gate593inter0), .b(s_28), .O(gate593inter1));
  and2  gate1079(.a(N1924), .b(N1896), .O(gate593inter2));
  inv1  gate1080(.a(s_28), .O(gate593inter3));
  inv1  gate1081(.a(s_29), .O(gate593inter4));
  nand2 gate1082(.a(gate593inter4), .b(gate593inter3), .O(gate593inter5));
  nor2  gate1083(.a(gate593inter5), .b(gate593inter2), .O(gate593inter6));
  inv1  gate1084(.a(N1896), .O(gate593inter7));
  inv1  gate1085(.a(N1924), .O(gate593inter8));
  nand2 gate1086(.a(gate593inter8), .b(gate593inter7), .O(gate593inter9));
  nand2 gate1087(.a(s_29), .b(gate593inter3), .O(gate593inter10));
  nor2  gate1088(.a(gate593inter10), .b(gate593inter9), .O(gate593inter11));
  nor2  gate1089(.a(gate593inter11), .b(gate593inter6), .O(gate593inter12));
  nand2 gate1090(.a(gate593inter12), .b(gate593inter1), .O(N1961));
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );

  xor2  gate2449(.a(N918), .b(N1927), .O(gate598inter0));
  nand2 gate2450(.a(gate598inter0), .b(s_224), .O(gate598inter1));
  and2  gate2451(.a(N918), .b(N1927), .O(gate598inter2));
  inv1  gate2452(.a(s_224), .O(gate598inter3));
  inv1  gate2453(.a(s_225), .O(gate598inter4));
  nand2 gate2454(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate2455(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate2456(.a(N1927), .O(gate598inter7));
  inv1  gate2457(.a(N918), .O(gate598inter8));
  nand2 gate2458(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate2459(.a(s_225), .b(gate598inter3), .O(gate598inter10));
  nor2  gate2460(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate2461(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate2462(.a(gate598inter12), .b(gate598inter1), .O(N1977));
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );

  xor2  gate1105(.a(N1499), .b(N1947), .O(gate607inter0));
  nand2 gate1106(.a(gate607inter0), .b(s_32), .O(gate607inter1));
  and2  gate1107(.a(N1499), .b(N1947), .O(gate607inter2));
  inv1  gate1108(.a(s_32), .O(gate607inter3));
  inv1  gate1109(.a(s_33), .O(gate607inter4));
  nand2 gate1110(.a(gate607inter4), .b(gate607inter3), .O(gate607inter5));
  nor2  gate1111(.a(gate607inter5), .b(gate607inter2), .O(gate607inter6));
  inv1  gate1112(.a(N1947), .O(gate607inter7));
  inv1  gate1113(.a(N1499), .O(gate607inter8));
  nand2 gate1114(.a(gate607inter8), .b(gate607inter7), .O(gate607inter9));
  nand2 gate1115(.a(s_33), .b(gate607inter3), .O(gate607inter10));
  nor2  gate1116(.a(gate607inter10), .b(gate607inter9), .O(gate607inter11));
  nor2  gate1117(.a(gate607inter11), .b(gate607inter6), .O(gate607inter12));
  nand2 gate1118(.a(gate607inter12), .b(gate607inter1), .O(N2003));

  xor2  gate2533(.a(N1350), .b(N1953), .O(gate608inter0));
  nand2 gate2534(.a(gate608inter0), .b(s_236), .O(gate608inter1));
  and2  gate2535(.a(N1350), .b(N1953), .O(gate608inter2));
  inv1  gate2536(.a(s_236), .O(gate608inter3));
  inv1  gate2537(.a(s_237), .O(gate608inter4));
  nand2 gate2538(.a(gate608inter4), .b(gate608inter3), .O(gate608inter5));
  nor2  gate2539(.a(gate608inter5), .b(gate608inter2), .O(gate608inter6));
  inv1  gate2540(.a(N1953), .O(gate608inter7));
  inv1  gate2541(.a(N1350), .O(gate608inter8));
  nand2 gate2542(.a(gate608inter8), .b(gate608inter7), .O(gate608inter9));
  nand2 gate2543(.a(s_237), .b(gate608inter3), .O(gate608inter10));
  nor2  gate2544(.a(gate608inter10), .b(gate608inter9), .O(gate608inter11));
  nor2  gate2545(.a(gate608inter11), .b(gate608inter6), .O(gate608inter12));
  nand2 gate2546(.a(gate608inter12), .b(gate608inter1), .O(N2004));
inv1 gate609( .a(N1953), .O(N2005) );

  xor2  gate2519(.a(N1351), .b(N1950), .O(gate610inter0));
  nand2 gate2520(.a(gate610inter0), .b(s_234), .O(gate610inter1));
  and2  gate2521(.a(N1351), .b(N1950), .O(gate610inter2));
  inv1  gate2522(.a(s_234), .O(gate610inter3));
  inv1  gate2523(.a(s_235), .O(gate610inter4));
  nand2 gate2524(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate2525(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate2526(.a(N1950), .O(gate610inter7));
  inv1  gate2527(.a(N1351), .O(gate610inter8));
  nand2 gate2528(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate2529(.a(s_235), .b(gate610inter3), .O(gate610inter10));
  nor2  gate2530(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate2531(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate2532(.a(gate610inter12), .b(gate610inter1), .O(N2006));
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate1903(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate1904(.a(gate612inter0), .b(s_146), .O(gate612inter1));
  and2  gate1905(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate1906(.a(s_146), .O(gate612inter3));
  inv1  gate1907(.a(s_147), .O(gate612inter4));
  nand2 gate1908(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate1909(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate1910(.a(N673), .O(gate612inter7));
  inv1  gate1911(.a(N1976), .O(gate612inter8));
  nand2 gate1912(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate1913(.a(s_147), .b(gate612inter3), .O(gate612inter10));
  nor2  gate1914(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate1915(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate1916(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );

  xor2  gate2239(.a(N1591), .b(N1987), .O(gate623inter0));
  nand2 gate2240(.a(gate623inter0), .b(s_194), .O(gate623inter1));
  and2  gate2241(.a(N1591), .b(N1987), .O(gate623inter2));
  inv1  gate2242(.a(s_194), .O(gate623inter3));
  inv1  gate2243(.a(s_195), .O(gate623inter4));
  nand2 gate2244(.a(gate623inter4), .b(gate623inter3), .O(gate623inter5));
  nor2  gate2245(.a(gate623inter5), .b(gate623inter2), .O(gate623inter6));
  inv1  gate2246(.a(N1987), .O(gate623inter7));
  inv1  gate2247(.a(N1591), .O(gate623inter8));
  nand2 gate2248(.a(gate623inter8), .b(gate623inter7), .O(gate623inter9));
  nand2 gate2249(.a(s_195), .b(gate623inter3), .O(gate623inter10));
  nor2  gate2250(.a(gate623inter10), .b(gate623inter9), .O(gate623inter11));
  nor2  gate2251(.a(gate623inter11), .b(gate623inter6), .O(gate623inter12));
  nand2 gate2252(.a(gate623inter12), .b(gate623inter1), .O(N2022));
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );

  xor2  gate1637(.a(N2005), .b(N1261), .O(gate625inter0));
  nand2 gate1638(.a(gate625inter0), .b(s_108), .O(gate625inter1));
  and2  gate1639(.a(N2005), .b(N1261), .O(gate625inter2));
  inv1  gate1640(.a(s_108), .O(gate625inter3));
  inv1  gate1641(.a(s_109), .O(gate625inter4));
  nand2 gate1642(.a(gate625inter4), .b(gate625inter3), .O(gate625inter5));
  nor2  gate1643(.a(gate625inter5), .b(gate625inter2), .O(gate625inter6));
  inv1  gate1644(.a(N1261), .O(gate625inter7));
  inv1  gate1645(.a(N2005), .O(gate625inter8));
  nand2 gate1646(.a(gate625inter8), .b(gate625inter7), .O(gate625inter9));
  nand2 gate1647(.a(s_109), .b(gate625inter3), .O(gate625inter10));
  nor2  gate1648(.a(gate625inter10), .b(gate625inter9), .O(gate625inter11));
  nor2  gate1649(.a(gate625inter11), .b(gate625inter6), .O(gate625inter12));
  nand2 gate1650(.a(gate625inter12), .b(gate625inter1), .O(N2024));
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );

  xor2  gate1679(.a(N2013), .b(N1875), .O(gate631inter0));
  nand2 gate1680(.a(gate631inter0), .b(s_114), .O(gate631inter1));
  and2  gate1681(.a(N2013), .b(N1875), .O(gate631inter2));
  inv1  gate1682(.a(s_114), .O(gate631inter3));
  inv1  gate1683(.a(s_115), .O(gate631inter4));
  nand2 gate1684(.a(gate631inter4), .b(gate631inter3), .O(gate631inter5));
  nor2  gate1685(.a(gate631inter5), .b(gate631inter2), .O(gate631inter6));
  inv1  gate1686(.a(N1875), .O(gate631inter7));
  inv1  gate1687(.a(N2013), .O(gate631inter8));
  nand2 gate1688(.a(gate631inter8), .b(gate631inter7), .O(gate631inter9));
  nand2 gate1689(.a(s_115), .b(gate631inter3), .O(gate631inter10));
  nor2  gate1690(.a(gate631inter10), .b(gate631inter9), .O(gate631inter11));
  nor2  gate1691(.a(gate631inter11), .b(gate631inter6), .O(gate631inter12));
  nand2 gate1692(.a(gate631inter12), .b(gate631inter1), .O(N2036));

  xor2  gate1553(.a(N2015), .b(N1571), .O(gate632inter0));
  nand2 gate1554(.a(gate632inter0), .b(s_96), .O(gate632inter1));
  and2  gate1555(.a(N2015), .b(N1571), .O(gate632inter2));
  inv1  gate1556(.a(s_96), .O(gate632inter3));
  inv1  gate1557(.a(s_97), .O(gate632inter4));
  nand2 gate1558(.a(gate632inter4), .b(gate632inter3), .O(gate632inter5));
  nor2  gate1559(.a(gate632inter5), .b(gate632inter2), .O(gate632inter6));
  inv1  gate1560(.a(N1571), .O(gate632inter7));
  inv1  gate1561(.a(N2015), .O(gate632inter8));
  nand2 gate1562(.a(gate632inter8), .b(gate632inter7), .O(gate632inter9));
  nand2 gate1563(.a(s_97), .b(gate632inter3), .O(gate632inter10));
  nor2  gate1564(.a(gate632inter10), .b(gate632inter9), .O(gate632inter11));
  nor2  gate1565(.a(gate632inter11), .b(gate632inter6), .O(gate632inter12));
  nand2 gate1566(.a(gate632inter12), .b(gate632inter1), .O(N2037));
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );

  xor2  gate1357(.a(N2003), .b(N2023), .O(gate635inter0));
  nand2 gate1358(.a(gate635inter0), .b(s_68), .O(gate635inter1));
  and2  gate1359(.a(N2003), .b(N2023), .O(gate635inter2));
  inv1  gate1360(.a(s_68), .O(gate635inter3));
  inv1  gate1361(.a(s_69), .O(gate635inter4));
  nand2 gate1362(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate1363(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate1364(.a(N2023), .O(gate635inter7));
  inv1  gate1365(.a(N2003), .O(gate635inter8));
  nand2 gate1366(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate1367(.a(s_69), .b(gate635inter3), .O(gate635inter10));
  nor2  gate1368(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate1369(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate1370(.a(gate635inter12), .b(gate635inter1), .O(N2040));
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );

  xor2  gate2631(.a(N2025), .b(N2006), .O(gate637inter0));
  nand2 gate2632(.a(gate637inter0), .b(s_250), .O(gate637inter1));
  and2  gate2633(.a(N2025), .b(N2006), .O(gate637inter2));
  inv1  gate2634(.a(s_250), .O(gate637inter3));
  inv1  gate2635(.a(s_251), .O(gate637inter4));
  nand2 gate2636(.a(gate637inter4), .b(gate637inter3), .O(gate637inter5));
  nor2  gate2637(.a(gate637inter5), .b(gate637inter2), .O(gate637inter6));
  inv1  gate2638(.a(N2006), .O(gate637inter7));
  inv1  gate2639(.a(N2025), .O(gate637inter8));
  nand2 gate2640(.a(gate637inter8), .b(gate637inter7), .O(gate637inter9));
  nand2 gate2641(.a(s_251), .b(gate637inter3), .O(gate637inter10));
  nor2  gate2642(.a(gate637inter10), .b(gate637inter9), .O(gate637inter11));
  nor2  gate2643(.a(gate637inter11), .b(gate637inter6), .O(gate637inter12));
  nand2 gate2644(.a(gate637inter12), .b(gate637inter1), .O(N2042));
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );

  xor2  gate2197(.a(N2022), .b(N2039), .O(gate642inter0));
  nand2 gate2198(.a(gate642inter0), .b(s_188), .O(gate642inter1));
  and2  gate2199(.a(N2022), .b(N2039), .O(gate642inter2));
  inv1  gate2200(.a(s_188), .O(gate642inter3));
  inv1  gate2201(.a(s_189), .O(gate642inter4));
  nand2 gate2202(.a(gate642inter4), .b(gate642inter3), .O(gate642inter5));
  nor2  gate2203(.a(gate642inter5), .b(gate642inter2), .O(gate642inter6));
  inv1  gate2204(.a(N2039), .O(gate642inter7));
  inv1  gate2205(.a(N2022), .O(gate642inter8));
  nand2 gate2206(.a(gate642inter8), .b(gate642inter7), .O(gate642inter9));
  nand2 gate2207(.a(s_189), .b(gate642inter3), .O(gate642inter10));
  nor2  gate2208(.a(gate642inter10), .b(gate642inter9), .O(gate642inter11));
  nor2  gate2209(.a(gate642inter11), .b(gate642inter6), .O(gate642inter12));
  nand2 gate2210(.a(gate642inter12), .b(gate642inter1), .O(N2061));
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );

  xor2  gate1371(.a(N915), .b(N2151), .O(gate663inter0));
  nand2 gate1372(.a(gate663inter0), .b(s_70), .O(gate663inter1));
  and2  gate1373(.a(N915), .b(N2151), .O(gate663inter2));
  inv1  gate1374(.a(s_70), .O(gate663inter3));
  inv1  gate1375(.a(s_71), .O(gate663inter4));
  nand2 gate1376(.a(gate663inter4), .b(gate663inter3), .O(gate663inter5));
  nor2  gate1377(.a(gate663inter5), .b(gate663inter2), .O(gate663inter6));
  inv1  gate1378(.a(N2151), .O(gate663inter7));
  inv1  gate1379(.a(N915), .O(gate663inter8));
  nand2 gate1380(.a(gate663inter8), .b(gate663inter7), .O(gate663inter9));
  nand2 gate1381(.a(s_71), .b(gate663inter3), .O(gate663inter10));
  nor2  gate1382(.a(gate663inter10), .b(gate663inter9), .O(gate663inter11));
  nor2  gate1383(.a(gate663inter11), .b(gate663inter6), .O(gate663inter12));
  nand2 gate1384(.a(gate663inter12), .b(gate663inter1), .O(N2214));
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate2505(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate2506(.a(gate667inter0), .b(s_232), .O(gate667inter1));
  and2  gate2507(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate2508(.a(s_232), .O(gate667inter3));
  inv1  gate2509(.a(s_233), .O(gate667inter4));
  nand2 gate2510(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate2511(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate2512(.a(N2199), .O(gate667inter7));
  inv1  gate2513(.a(N1348), .O(gate667inter8));
  nand2 gate2514(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate2515(.a(s_233), .b(gate667inter3), .O(gate667inter10));
  nor2  gate2516(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate2517(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate2518(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );

  xor2  gate1833(.a(N1349), .b(N2196), .O(gate669inter0));
  nand2 gate1834(.a(gate669inter0), .b(s_136), .O(gate669inter1));
  and2  gate1835(.a(N1349), .b(N2196), .O(gate669inter2));
  inv1  gate1836(.a(s_136), .O(gate669inter3));
  inv1  gate1837(.a(s_137), .O(gate669inter4));
  nand2 gate1838(.a(gate669inter4), .b(gate669inter3), .O(gate669inter5));
  nor2  gate1839(.a(gate669inter5), .b(gate669inter2), .O(gate669inter6));
  inv1  gate1840(.a(N2196), .O(gate669inter7));
  inv1  gate1841(.a(N1349), .O(gate669inter8));
  nand2 gate1842(.a(gate669inter8), .b(gate669inter7), .O(gate669inter9));
  nand2 gate1843(.a(s_137), .b(gate669inter3), .O(gate669inter10));
  nor2  gate1844(.a(gate669inter10), .b(gate669inter9), .O(gate669inter11));
  nor2  gate1845(.a(gate669inter11), .b(gate669inter6), .O(gate669inter12));
  nand2 gate1846(.a(gate669inter12), .b(gate669inter1), .O(N2224));
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate1945(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate1946(.a(gate671inter0), .b(s_152), .O(gate671inter1));
  and2  gate1947(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate1948(.a(s_152), .O(gate671inter3));
  inv1  gate1949(.a(s_153), .O(gate671inter4));
  nand2 gate1950(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate1951(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate1952(.a(N2205), .O(gate671inter7));
  inv1  gate1953(.a(N913), .O(gate671inter8));
  nand2 gate1954(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate1955(.a(s_153), .b(gate671inter3), .O(gate671inter10));
  nor2  gate1956(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate1957(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate1958(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );

  xor2  gate923(.a(N914), .b(N2202), .O(gate673inter0));
  nand2 gate924(.a(gate673inter0), .b(s_6), .O(gate673inter1));
  and2  gate925(.a(N914), .b(N2202), .O(gate673inter2));
  inv1  gate926(.a(s_6), .O(gate673inter3));
  inv1  gate927(.a(s_7), .O(gate673inter4));
  nand2 gate928(.a(gate673inter4), .b(gate673inter3), .O(gate673inter5));
  nor2  gate929(.a(gate673inter5), .b(gate673inter2), .O(gate673inter6));
  inv1  gate930(.a(N2202), .O(gate673inter7));
  inv1  gate931(.a(N914), .O(gate673inter8));
  nand2 gate932(.a(gate673inter8), .b(gate673inter7), .O(gate673inter9));
  nand2 gate933(.a(s_7), .b(gate673inter3), .O(gate673inter10));
  nor2  gate934(.a(gate673inter10), .b(gate673inter9), .O(gate673inter11));
  nor2  gate935(.a(gate673inter11), .b(gate673inter6), .O(gate673inter12));
  nand2 gate936(.a(gate673inter12), .b(gate673inter1), .O(N2228));
inv1 gate674( .a(N2202), .O(N2229) );

  xor2  gate2141(.a(N2215), .b(N667), .O(gate675inter0));
  nand2 gate2142(.a(gate675inter0), .b(s_180), .O(gate675inter1));
  and2  gate2143(.a(N2215), .b(N667), .O(gate675inter2));
  inv1  gate2144(.a(s_180), .O(gate675inter3));
  inv1  gate2145(.a(s_181), .O(gate675inter4));
  nand2 gate2146(.a(gate675inter4), .b(gate675inter3), .O(gate675inter5));
  nor2  gate2147(.a(gate675inter5), .b(gate675inter2), .O(gate675inter6));
  inv1  gate2148(.a(N667), .O(gate675inter7));
  inv1  gate2149(.a(N2215), .O(gate675inter8));
  nand2 gate2150(.a(gate675inter8), .b(gate675inter7), .O(gate675inter9));
  nand2 gate2151(.a(s_181), .b(gate675inter3), .O(gate675inter10));
  nor2  gate2152(.a(gate675inter10), .b(gate675inter9), .O(gate675inter11));
  nor2  gate2153(.a(gate675inter11), .b(gate675inter6), .O(gate675inter12));
  nand2 gate2154(.a(gate675inter12), .b(gate675inter1), .O(N2230));

  xor2  gate2169(.a(N2217), .b(N664), .O(gate676inter0));
  nand2 gate2170(.a(gate676inter0), .b(s_184), .O(gate676inter1));
  and2  gate2171(.a(N2217), .b(N664), .O(gate676inter2));
  inv1  gate2172(.a(s_184), .O(gate676inter3));
  inv1  gate2173(.a(s_185), .O(gate676inter4));
  nand2 gate2174(.a(gate676inter4), .b(gate676inter3), .O(gate676inter5));
  nor2  gate2175(.a(gate676inter5), .b(gate676inter2), .O(gate676inter6));
  inv1  gate2176(.a(N664), .O(gate676inter7));
  inv1  gate2177(.a(N2217), .O(gate676inter8));
  nand2 gate2178(.a(gate676inter8), .b(gate676inter7), .O(gate676inter9));
  nand2 gate2179(.a(s_185), .b(gate676inter3), .O(gate676inter10));
  nor2  gate2180(.a(gate676inter10), .b(gate676inter9), .O(gate676inter11));
  nor2  gate2181(.a(gate676inter11), .b(gate676inter6), .O(gate676inter12));
  nand2 gate2182(.a(gate676inter12), .b(gate676inter1), .O(N2231));
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );

  xor2  gate1427(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate1428(.a(gate678inter0), .b(s_78), .O(gate678inter1));
  and2  gate1429(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate1430(.a(s_78), .O(gate678inter3));
  inv1  gate1431(.a(s_79), .O(gate678inter4));
  nand2 gate1432(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate1433(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate1434(.a(N1252), .O(gate678inter7));
  inv1  gate1435(.a(N2225), .O(gate678inter8));
  nand2 gate1436(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate1437(.a(s_79), .b(gate678inter3), .O(gate678inter10));
  nor2  gate1438(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate1439(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate1440(.a(gate678inter12), .b(gate678inter1), .O(N2233));
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );

  xor2  gate2043(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate2044(.a(gate684inter0), .b(s_166), .O(gate684inter1));
  and2  gate2045(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate2046(.a(s_166), .O(gate684inter3));
  inv1  gate2047(.a(s_167), .O(gate684inter4));
  nand2 gate2048(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate2049(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate2050(.a(N2224), .O(gate684inter7));
  inv1  gate2051(.a(N2233), .O(gate684inter8));
  nand2 gate2052(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate2053(.a(s_167), .b(gate684inter3), .O(gate684inter10));
  nor2  gate2054(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate2055(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate2056(.a(gate684inter12), .b(gate684inter1), .O(N2241));
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );

  xor2  gate1497(.a(N2235), .b(N2228), .O(gate686inter0));
  nand2 gate1498(.a(gate686inter0), .b(s_88), .O(gate686inter1));
  and2  gate1499(.a(N2235), .b(N2228), .O(gate686inter2));
  inv1  gate1500(.a(s_88), .O(gate686inter3));
  inv1  gate1501(.a(s_89), .O(gate686inter4));
  nand2 gate1502(.a(gate686inter4), .b(gate686inter3), .O(gate686inter5));
  nor2  gate1503(.a(gate686inter5), .b(gate686inter2), .O(gate686inter6));
  inv1  gate1504(.a(N2228), .O(gate686inter7));
  inv1  gate1505(.a(N2235), .O(gate686inter8));
  nand2 gate1506(.a(gate686inter8), .b(gate686inter7), .O(gate686inter9));
  nand2 gate1507(.a(s_89), .b(gate686inter3), .O(gate686inter10));
  nor2  gate1508(.a(gate686inter10), .b(gate686inter9), .O(gate686inter11));
  nor2  gate1509(.a(gate686inter11), .b(gate686inter6), .O(gate686inter12));
  nand2 gate1510(.a(gate686inter12), .b(gate686inter1), .O(N2245));
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate1329(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate1330(.a(gate754inter0), .b(s_64), .O(gate754inter1));
  and2  gate1331(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate1332(.a(s_64), .O(gate754inter3));
  inv1  gate1333(.a(s_65), .O(gate754inter4));
  nand2 gate1334(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1335(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1336(.a(N2564), .O(gate754inter7));
  inv1  gate1337(.a(N536), .O(gate754inter8));
  nand2 gate1338(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1339(.a(s_65), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1340(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1341(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1342(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );

  xor2  gate1693(.a(N543), .b(N2570), .O(gate758inter0));
  nand2 gate1694(.a(gate758inter0), .b(s_116), .O(gate758inter1));
  and2  gate1695(.a(N543), .b(N2570), .O(gate758inter2));
  inv1  gate1696(.a(s_116), .O(gate758inter3));
  inv1  gate1697(.a(s_117), .O(gate758inter4));
  nand2 gate1698(.a(gate758inter4), .b(gate758inter3), .O(gate758inter5));
  nor2  gate1699(.a(gate758inter5), .b(gate758inter2), .O(gate758inter6));
  inv1  gate1700(.a(N2570), .O(gate758inter7));
  inv1  gate1701(.a(N543), .O(gate758inter8));
  nand2 gate1702(.a(gate758inter8), .b(gate758inter7), .O(gate758inter9));
  nand2 gate1703(.a(s_117), .b(gate758inter3), .O(gate758inter10));
  nor2  gate1704(.a(gate758inter10), .b(gate758inter9), .O(gate758inter11));
  nor2  gate1705(.a(gate758inter11), .b(gate758inter6), .O(gate758inter12));
  nand2 gate1706(.a(gate758inter12), .b(gate758inter1), .O(N2682));
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );

  xor2  gate1119(.a(N2670), .b(N343), .O(gate765inter0));
  nand2 gate1120(.a(gate765inter0), .b(s_34), .O(gate765inter1));
  and2  gate1121(.a(N2670), .b(N343), .O(gate765inter2));
  inv1  gate1122(.a(s_34), .O(gate765inter3));
  inv1  gate1123(.a(s_35), .O(gate765inter4));
  nand2 gate1124(.a(gate765inter4), .b(gate765inter3), .O(gate765inter5));
  nor2  gate1125(.a(gate765inter5), .b(gate765inter2), .O(gate765inter6));
  inv1  gate1126(.a(N343), .O(gate765inter7));
  inv1  gate1127(.a(N2670), .O(gate765inter8));
  nand2 gate1128(.a(gate765inter8), .b(gate765inter7), .O(gate765inter9));
  nand2 gate1129(.a(s_35), .b(gate765inter3), .O(gate765inter10));
  nor2  gate1130(.a(gate765inter10), .b(gate765inter9), .O(gate765inter11));
  nor2  gate1131(.a(gate765inter11), .b(gate765inter6), .O(gate765inter12));
  nand2 gate1132(.a(gate765inter12), .b(gate765inter1), .O(N2720));
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );

  xor2  gate1203(.a(N2674), .b(N349), .O(gate767inter0));
  nand2 gate1204(.a(gate767inter0), .b(s_46), .O(gate767inter1));
  and2  gate1205(.a(N2674), .b(N349), .O(gate767inter2));
  inv1  gate1206(.a(s_46), .O(gate767inter3));
  inv1  gate1207(.a(s_47), .O(gate767inter4));
  nand2 gate1208(.a(gate767inter4), .b(gate767inter3), .O(gate767inter5));
  nor2  gate1209(.a(gate767inter5), .b(gate767inter2), .O(gate767inter6));
  inv1  gate1210(.a(N349), .O(gate767inter7));
  inv1  gate1211(.a(N2674), .O(gate767inter8));
  nand2 gate1212(.a(gate767inter8), .b(gate767inter7), .O(gate767inter9));
  nand2 gate1213(.a(s_47), .b(gate767inter3), .O(gate767inter10));
  nor2  gate1214(.a(gate767inter10), .b(gate767inter9), .O(gate767inter11));
  nor2  gate1215(.a(gate767inter11), .b(gate767inter6), .O(gate767inter12));
  nand2 gate1216(.a(gate767inter12), .b(gate767inter1), .O(N2722));
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );

  xor2  gate2029(.a(N539), .b(N2642), .O(gate771inter0));
  nand2 gate2030(.a(gate771inter0), .b(s_164), .O(gate771inter1));
  and2  gate2031(.a(N539), .b(N2642), .O(gate771inter2));
  inv1  gate2032(.a(s_164), .O(gate771inter3));
  inv1  gate2033(.a(s_165), .O(gate771inter4));
  nand2 gate2034(.a(gate771inter4), .b(gate771inter3), .O(gate771inter5));
  nor2  gate2035(.a(gate771inter5), .b(gate771inter2), .O(gate771inter6));
  inv1  gate2036(.a(N2642), .O(gate771inter7));
  inv1  gate2037(.a(N539), .O(gate771inter8));
  nand2 gate2038(.a(gate771inter8), .b(gate771inter7), .O(gate771inter9));
  nand2 gate2039(.a(s_165), .b(gate771inter3), .O(gate771inter10));
  nor2  gate2040(.a(gate771inter10), .b(gate771inter9), .O(gate771inter11));
  nor2  gate2041(.a(gate771inter11), .b(gate771inter6), .O(gate771inter12));
  nand2 gate2042(.a(gate771inter12), .b(gate771inter1), .O(N2726));
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate2071(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate2072(.a(gate773inter0), .b(s_170), .O(gate773inter1));
  and2  gate2073(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate2074(.a(s_170), .O(gate773inter3));
  inv1  gate2075(.a(s_171), .O(gate773inter4));
  nand2 gate2076(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate2077(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate2078(.a(N2645), .O(gate773inter7));
  inv1  gate2079(.a(N540), .O(gate773inter8));
  nand2 gate2080(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate2081(.a(s_171), .b(gate773inter3), .O(gate773inter10));
  nor2  gate2082(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate2083(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate2084(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );

  xor2  gate1917(.a(N541), .b(N2648), .O(gate775inter0));
  nand2 gate1918(.a(gate775inter0), .b(s_148), .O(gate775inter1));
  and2  gate1919(.a(N541), .b(N2648), .O(gate775inter2));
  inv1  gate1920(.a(s_148), .O(gate775inter3));
  inv1  gate1921(.a(s_149), .O(gate775inter4));
  nand2 gate1922(.a(gate775inter4), .b(gate775inter3), .O(gate775inter5));
  nor2  gate1923(.a(gate775inter5), .b(gate775inter2), .O(gate775inter6));
  inv1  gate1924(.a(N2648), .O(gate775inter7));
  inv1  gate1925(.a(N541), .O(gate775inter8));
  nand2 gate1926(.a(gate775inter8), .b(gate775inter7), .O(gate775inter9));
  nand2 gate1927(.a(s_149), .b(gate775inter3), .O(gate775inter10));
  nor2  gate1928(.a(gate775inter10), .b(gate775inter9), .O(gate775inter11));
  nor2  gate1929(.a(gate775inter11), .b(gate775inter6), .O(gate775inter12));
  nand2 gate1930(.a(gate775inter12), .b(gate775inter1), .O(N2730));
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );

  xor2  gate1665(.a(N544), .b(N2655), .O(gate780inter0));
  nand2 gate1666(.a(gate780inter0), .b(s_112), .O(gate780inter1));
  and2  gate1667(.a(N544), .b(N2655), .O(gate780inter2));
  inv1  gate1668(.a(s_112), .O(gate780inter3));
  inv1  gate1669(.a(s_113), .O(gate780inter4));
  nand2 gate1670(.a(gate780inter4), .b(gate780inter3), .O(gate780inter5));
  nor2  gate1671(.a(gate780inter5), .b(gate780inter2), .O(gate780inter6));
  inv1  gate1672(.a(N2655), .O(gate780inter7));
  inv1  gate1673(.a(N544), .O(gate780inter8));
  nand2 gate1674(.a(gate780inter8), .b(gate780inter7), .O(gate780inter9));
  nand2 gate1675(.a(s_113), .b(gate780inter3), .O(gate780inter10));
  nor2  gate1676(.a(gate780inter10), .b(gate780inter9), .O(gate780inter11));
  nor2  gate1677(.a(gate780inter11), .b(gate780inter6), .O(gate780inter12));
  nand2 gate1678(.a(gate780inter12), .b(gate780inter1), .O(N2735));
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate2127(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate2128(.a(gate788inter0), .b(s_178), .O(gate788inter1));
  and2  gate2129(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate2130(.a(s_178), .O(gate788inter3));
  inv1  gate2131(.a(s_179), .O(gate788inter4));
  nand2 gate2132(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate2133(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate2134(.a(N385), .O(gate788inter7));
  inv1  gate2135(.a(N2689), .O(gate788inter8));
  nand2 gate2136(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate2137(.a(s_179), .b(gate788inter3), .O(gate788inter10));
  nor2  gate2138(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate2139(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate2140(.a(gate788inter12), .b(gate788inter1), .O(N2743));
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );

  xor2  gate1175(.a(N2720), .b(N2669), .O(gate794inter0));
  nand2 gate1176(.a(gate794inter0), .b(s_42), .O(gate794inter1));
  and2  gate1177(.a(N2720), .b(N2669), .O(gate794inter2));
  inv1  gate1178(.a(s_42), .O(gate794inter3));
  inv1  gate1179(.a(s_43), .O(gate794inter4));
  nand2 gate1180(.a(gate794inter4), .b(gate794inter3), .O(gate794inter5));
  nor2  gate1181(.a(gate794inter5), .b(gate794inter2), .O(gate794inter6));
  inv1  gate1182(.a(N2669), .O(gate794inter7));
  inv1  gate1183(.a(N2720), .O(gate794inter8));
  nand2 gate1184(.a(gate794inter8), .b(gate794inter7), .O(gate794inter9));
  nand2 gate1185(.a(s_43), .b(gate794inter3), .O(gate794inter10));
  nor2  gate1186(.a(gate794inter10), .b(gate794inter9), .O(gate794inter11));
  nor2  gate1187(.a(gate794inter11), .b(gate794inter6), .O(gate794inter12));
  nand2 gate1188(.a(gate794inter12), .b(gate794inter1), .O(N2753));

  xor2  gate2421(.a(N2721), .b(N2671), .O(gate795inter0));
  nand2 gate2422(.a(gate795inter0), .b(s_220), .O(gate795inter1));
  and2  gate2423(.a(N2721), .b(N2671), .O(gate795inter2));
  inv1  gate2424(.a(s_220), .O(gate795inter3));
  inv1  gate2425(.a(s_221), .O(gate795inter4));
  nand2 gate2426(.a(gate795inter4), .b(gate795inter3), .O(gate795inter5));
  nor2  gate2427(.a(gate795inter5), .b(gate795inter2), .O(gate795inter6));
  inv1  gate2428(.a(N2671), .O(gate795inter7));
  inv1  gate2429(.a(N2721), .O(gate795inter8));
  nand2 gate2430(.a(gate795inter8), .b(gate795inter7), .O(gate795inter9));
  nand2 gate2431(.a(s_221), .b(gate795inter3), .O(gate795inter10));
  nor2  gate2432(.a(gate795inter10), .b(gate795inter9), .O(gate795inter11));
  nor2  gate2433(.a(gate795inter11), .b(gate795inter6), .O(gate795inter12));
  nand2 gate2434(.a(gate795inter12), .b(gate795inter1), .O(N2754));
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );

  xor2  gate1385(.a(N2723), .b(N2675), .O(gate797inter0));
  nand2 gate1386(.a(gate797inter0), .b(s_72), .O(gate797inter1));
  and2  gate1387(.a(N2723), .b(N2675), .O(gate797inter2));
  inv1  gate1388(.a(s_72), .O(gate797inter3));
  inv1  gate1389(.a(s_73), .O(gate797inter4));
  nand2 gate1390(.a(gate797inter4), .b(gate797inter3), .O(gate797inter5));
  nor2  gate1391(.a(gate797inter5), .b(gate797inter2), .O(gate797inter6));
  inv1  gate1392(.a(N2675), .O(gate797inter7));
  inv1  gate1393(.a(N2723), .O(gate797inter8));
  nand2 gate1394(.a(gate797inter8), .b(gate797inter7), .O(gate797inter9));
  nand2 gate1395(.a(s_73), .b(gate797inter3), .O(gate797inter10));
  nor2  gate1396(.a(gate797inter10), .b(gate797inter9), .O(gate797inter11));
  nor2  gate1397(.a(gate797inter11), .b(gate797inter6), .O(gate797inter12));
  nand2 gate1398(.a(gate797inter12), .b(gate797inter1), .O(N2756));

  xor2  gate2365(.a(N2725), .b(N355), .O(gate798inter0));
  nand2 gate2366(.a(gate798inter0), .b(s_212), .O(gate798inter1));
  and2  gate2367(.a(N2725), .b(N355), .O(gate798inter2));
  inv1  gate2368(.a(s_212), .O(gate798inter3));
  inv1  gate2369(.a(s_213), .O(gate798inter4));
  nand2 gate2370(.a(gate798inter4), .b(gate798inter3), .O(gate798inter5));
  nor2  gate2371(.a(gate798inter5), .b(gate798inter2), .O(gate798inter6));
  inv1  gate2372(.a(N355), .O(gate798inter7));
  inv1  gate2373(.a(N2725), .O(gate798inter8));
  nand2 gate2374(.a(gate798inter8), .b(gate798inter7), .O(gate798inter9));
  nand2 gate2375(.a(s_213), .b(gate798inter3), .O(gate798inter10));
  nor2  gate2376(.a(gate798inter10), .b(gate798inter9), .O(gate798inter11));
  nor2  gate2377(.a(gate798inter11), .b(gate798inter6), .O(gate798inter12));
  nand2 gate2378(.a(gate798inter12), .b(gate798inter1), .O(N2757));
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );

  xor2  gate979(.a(N2731), .b(N364), .O(gate801inter0));
  nand2 gate980(.a(gate801inter0), .b(s_14), .O(gate801inter1));
  and2  gate981(.a(N2731), .b(N364), .O(gate801inter2));
  inv1  gate982(.a(s_14), .O(gate801inter3));
  inv1  gate983(.a(s_15), .O(gate801inter4));
  nand2 gate984(.a(gate801inter4), .b(gate801inter3), .O(gate801inter5));
  nor2  gate985(.a(gate801inter5), .b(gate801inter2), .O(gate801inter6));
  inv1  gate986(.a(N364), .O(gate801inter7));
  inv1  gate987(.a(N2731), .O(gate801inter8));
  nand2 gate988(.a(gate801inter8), .b(gate801inter7), .O(gate801inter9));
  nand2 gate989(.a(s_15), .b(gate801inter3), .O(gate801inter10));
  nor2  gate990(.a(gate801inter10), .b(gate801inter9), .O(gate801inter11));
  nor2  gate991(.a(gate801inter11), .b(gate801inter6), .O(gate801inter12));
  nand2 gate992(.a(gate801inter12), .b(gate801inter1), .O(N2760));

  xor2  gate2351(.a(N2733), .b(N367), .O(gate802inter0));
  nand2 gate2352(.a(gate802inter0), .b(s_210), .O(gate802inter1));
  and2  gate2353(.a(N2733), .b(N367), .O(gate802inter2));
  inv1  gate2354(.a(s_210), .O(gate802inter3));
  inv1  gate2355(.a(s_211), .O(gate802inter4));
  nand2 gate2356(.a(gate802inter4), .b(gate802inter3), .O(gate802inter5));
  nor2  gate2357(.a(gate802inter5), .b(gate802inter2), .O(gate802inter6));
  inv1  gate2358(.a(N367), .O(gate802inter7));
  inv1  gate2359(.a(N2733), .O(gate802inter8));
  nand2 gate2360(.a(gate802inter8), .b(gate802inter7), .O(gate802inter9));
  nand2 gate2361(.a(s_211), .b(gate802inter3), .O(gate802inter10));
  nor2  gate2362(.a(gate802inter10), .b(gate802inter9), .O(gate802inter11));
  nor2  gate2363(.a(gate802inter11), .b(gate802inter6), .O(gate802inter12));
  nand2 gate2364(.a(gate802inter12), .b(gate802inter1), .O(N2761));
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );

  xor2  gate1007(.a(N2738), .b(N376), .O(gate805inter0));
  nand2 gate1008(.a(gate805inter0), .b(s_18), .O(gate805inter1));
  and2  gate1009(.a(N2738), .b(N376), .O(gate805inter2));
  inv1  gate1010(.a(s_18), .O(gate805inter3));
  inv1  gate1011(.a(s_19), .O(gate805inter4));
  nand2 gate1012(.a(gate805inter4), .b(gate805inter3), .O(gate805inter5));
  nor2  gate1013(.a(gate805inter5), .b(gate805inter2), .O(gate805inter6));
  inv1  gate1014(.a(N376), .O(gate805inter7));
  inv1  gate1015(.a(N2738), .O(gate805inter8));
  nand2 gate1016(.a(gate805inter8), .b(gate805inter7), .O(gate805inter9));
  nand2 gate1017(.a(s_19), .b(gate805inter3), .O(gate805inter10));
  nor2  gate1018(.a(gate805inter10), .b(gate805inter9), .O(gate805inter11));
  nor2  gate1019(.a(gate805inter11), .b(gate805inter6), .O(gate805inter12));
  nand2 gate1020(.a(gate805inter12), .b(gate805inter1), .O(N2764));
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );

  xor2  gate1959(.a(N2742), .b(N382), .O(gate807inter0));
  nand2 gate1960(.a(gate807inter0), .b(s_154), .O(gate807inter1));
  and2  gate1961(.a(N2742), .b(N382), .O(gate807inter2));
  inv1  gate1962(.a(s_154), .O(gate807inter3));
  inv1  gate1963(.a(s_155), .O(gate807inter4));
  nand2 gate1964(.a(gate807inter4), .b(gate807inter3), .O(gate807inter5));
  nor2  gate1965(.a(gate807inter5), .b(gate807inter2), .O(gate807inter6));
  inv1  gate1966(.a(N382), .O(gate807inter7));
  inv1  gate1967(.a(N2742), .O(gate807inter8));
  nand2 gate1968(.a(gate807inter8), .b(gate807inter7), .O(gate807inter9));
  nand2 gate1969(.a(s_155), .b(gate807inter3), .O(gate807inter10));
  nor2  gate1970(.a(gate807inter10), .b(gate807inter9), .O(gate807inter11));
  nor2  gate1971(.a(gate807inter11), .b(gate807inter6), .O(gate807inter12));
  nand2 gate1972(.a(gate807inter12), .b(gate807inter1), .O(N2766));
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );

  xor2  gate2561(.a(N2757), .b(N2724), .O(gate812inter0));
  nand2 gate2562(.a(gate812inter0), .b(s_240), .O(gate812inter1));
  and2  gate2563(.a(N2757), .b(N2724), .O(gate812inter2));
  inv1  gate2564(.a(s_240), .O(gate812inter3));
  inv1  gate2565(.a(s_241), .O(gate812inter4));
  nand2 gate2566(.a(gate812inter4), .b(gate812inter3), .O(gate812inter5));
  nor2  gate2567(.a(gate812inter5), .b(gate812inter2), .O(gate812inter6));
  inv1  gate2568(.a(N2724), .O(gate812inter7));
  inv1  gate2569(.a(N2757), .O(gate812inter8));
  nand2 gate2570(.a(gate812inter8), .b(gate812inter7), .O(gate812inter9));
  nand2 gate2571(.a(s_241), .b(gate812inter3), .O(gate812inter10));
  nor2  gate2572(.a(gate812inter10), .b(gate812inter9), .O(gate812inter11));
  nor2  gate2573(.a(gate812inter11), .b(gate812inter6), .O(gate812inter12));
  nand2 gate2574(.a(gate812inter12), .b(gate812inter1), .O(N2779));
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );

  xor2  gate965(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate966(.a(gate815inter0), .b(s_12), .O(gate815inter1));
  and2  gate967(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate968(.a(s_12), .O(gate815inter3));
  inv1  gate969(.a(s_13), .O(gate815inter4));
  nand2 gate970(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate971(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate972(.a(N2730), .O(gate815inter7));
  inv1  gate973(.a(N2760), .O(gate815inter8));
  nand2 gate974(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate975(.a(s_13), .b(gate815inter3), .O(gate815inter10));
  nor2  gate976(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate977(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate978(.a(gate815inter12), .b(gate815inter1), .O(N2782));
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );

  xor2  gate2337(.a(N2763), .b(N2735), .O(gate817inter0));
  nand2 gate2338(.a(gate817inter0), .b(s_208), .O(gate817inter1));
  and2  gate2339(.a(N2763), .b(N2735), .O(gate817inter2));
  inv1  gate2340(.a(s_208), .O(gate817inter3));
  inv1  gate2341(.a(s_209), .O(gate817inter4));
  nand2 gate2342(.a(gate817inter4), .b(gate817inter3), .O(gate817inter5));
  nor2  gate2343(.a(gate817inter5), .b(gate817inter2), .O(gate817inter6));
  inv1  gate2344(.a(N2735), .O(gate817inter7));
  inv1  gate2345(.a(N2763), .O(gate817inter8));
  nand2 gate2346(.a(gate817inter8), .b(gate817inter7), .O(gate817inter9));
  nand2 gate2347(.a(s_209), .b(gate817inter3), .O(gate817inter10));
  nor2  gate2348(.a(gate817inter10), .b(gate817inter9), .O(gate817inter11));
  nor2  gate2349(.a(gate817inter11), .b(gate817inter6), .O(gate817inter12));
  nand2 gate2350(.a(gate817inter12), .b(gate817inter1), .O(N2784));

  xor2  gate2113(.a(N2764), .b(N2737), .O(gate818inter0));
  nand2 gate2114(.a(gate818inter0), .b(s_176), .O(gate818inter1));
  and2  gate2115(.a(N2764), .b(N2737), .O(gate818inter2));
  inv1  gate2116(.a(s_176), .O(gate818inter3));
  inv1  gate2117(.a(s_177), .O(gate818inter4));
  nand2 gate2118(.a(gate818inter4), .b(gate818inter3), .O(gate818inter5));
  nor2  gate2119(.a(gate818inter5), .b(gate818inter2), .O(gate818inter6));
  inv1  gate2120(.a(N2737), .O(gate818inter7));
  inv1  gate2121(.a(N2764), .O(gate818inter8));
  nand2 gate2122(.a(gate818inter8), .b(gate818inter7), .O(gate818inter9));
  nand2 gate2123(.a(s_177), .b(gate818inter3), .O(gate818inter10));
  nor2  gate2124(.a(gate818inter10), .b(gate818inter9), .O(gate818inter11));
  nor2  gate2125(.a(gate818inter11), .b(gate818inter6), .O(gate818inter12));
  nand2 gate2126(.a(gate818inter12), .b(gate818inter1), .O(N2785));
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );

  xor2  gate881(.a(N2018), .b(N2773), .O(gate824inter0));
  nand2 gate882(.a(gate824inter0), .b(s_0), .O(gate824inter1));
  and2  gate883(.a(N2018), .b(N2773), .O(gate824inter2));
  inv1  gate884(.a(s_0), .O(gate824inter3));
  inv1  gate885(.a(s_1), .O(gate824inter4));
  nand2 gate886(.a(gate824inter4), .b(gate824inter3), .O(gate824inter5));
  nor2  gate887(.a(gate824inter5), .b(gate824inter2), .O(gate824inter6));
  inv1  gate888(.a(N2773), .O(gate824inter7));
  inv1  gate889(.a(N2018), .O(gate824inter8));
  nand2 gate890(.a(gate824inter8), .b(gate824inter7), .O(gate824inter9));
  nand2 gate891(.a(s_1), .b(gate824inter3), .O(gate824inter10));
  nor2  gate892(.a(gate824inter10), .b(gate824inter9), .O(gate824inter11));
  nor2  gate893(.a(gate824inter11), .b(gate824inter6), .O(gate824inter12));
  nand2 gate894(.a(gate824inter12), .b(gate824inter1), .O(N2807));
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );

  xor2  gate1539(.a(N2857), .b(N2052), .O(gate851inter0));
  nand2 gate1540(.a(gate851inter0), .b(s_94), .O(gate851inter1));
  and2  gate1541(.a(N2857), .b(N2052), .O(gate851inter2));
  inv1  gate1542(.a(s_94), .O(gate851inter3));
  inv1  gate1543(.a(s_95), .O(gate851inter4));
  nand2 gate1544(.a(gate851inter4), .b(gate851inter3), .O(gate851inter5));
  nor2  gate1545(.a(gate851inter5), .b(gate851inter2), .O(gate851inter6));
  inv1  gate1546(.a(N2052), .O(gate851inter7));
  inv1  gate1547(.a(N2857), .O(gate851inter8));
  nand2 gate1548(.a(gate851inter8), .b(gate851inter7), .O(gate851inter9));
  nand2 gate1549(.a(s_95), .b(gate851inter3), .O(gate851inter10));
  nor2  gate1550(.a(gate851inter10), .b(gate851inter9), .O(gate851inter11));
  nor2  gate1551(.a(gate851inter11), .b(gate851inter6), .O(gate851inter12));
  nand2 gate1552(.a(gate851inter12), .b(gate851inter1), .O(N2866));
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );

  xor2  gate1161(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1162(.a(gate856inter0), .b(s_40), .O(gate856inter1));
  and2  gate1163(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1164(.a(s_40), .O(gate856inter3));
  inv1  gate1165(.a(s_41), .O(gate856inter4));
  nand2 gate1166(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1167(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1168(.a(N2843), .O(gate856inter7));
  inv1  gate1169(.a(N886), .O(gate856inter8));
  nand2 gate1170(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1171(.a(s_41), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1172(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1173(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1174(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );

  xor2  gate1483(.a(N2851), .b(N2867), .O(gate862inter0));
  nand2 gate1484(.a(gate862inter0), .b(s_86), .O(gate862inter1));
  and2  gate1485(.a(N2851), .b(N2867), .O(gate862inter2));
  inv1  gate1486(.a(s_86), .O(gate862inter3));
  inv1  gate1487(.a(s_87), .O(gate862inter4));
  nand2 gate1488(.a(gate862inter4), .b(gate862inter3), .O(gate862inter5));
  nor2  gate1489(.a(gate862inter5), .b(gate862inter2), .O(gate862inter6));
  inv1  gate1490(.a(N2867), .O(gate862inter7));
  inv1  gate1491(.a(N2851), .O(gate862inter8));
  nand2 gate1492(.a(gate862inter8), .b(gate862inter7), .O(gate862inter9));
  nand2 gate1493(.a(s_87), .b(gate862inter3), .O(gate862inter10));
  nor2  gate1494(.a(gate862inter10), .b(gate862inter9), .O(gate862inter11));
  nor2  gate1495(.a(gate862inter11), .b(gate862inter6), .O(gate862inter12));
  nand2 gate1496(.a(gate862inter12), .b(gate862inter1), .O(N2877));

  xor2  gate1287(.a(N2852), .b(N2868), .O(gate863inter0));
  nand2 gate1288(.a(gate863inter0), .b(s_58), .O(gate863inter1));
  and2  gate1289(.a(N2852), .b(N2868), .O(gate863inter2));
  inv1  gate1290(.a(s_58), .O(gate863inter3));
  inv1  gate1291(.a(s_59), .O(gate863inter4));
  nand2 gate1292(.a(gate863inter4), .b(gate863inter3), .O(gate863inter5));
  nor2  gate1293(.a(gate863inter5), .b(gate863inter2), .O(gate863inter6));
  inv1  gate1294(.a(N2868), .O(gate863inter7));
  inv1  gate1295(.a(N2852), .O(gate863inter8));
  nand2 gate1296(.a(gate863inter8), .b(gate863inter7), .O(gate863inter9));
  nand2 gate1297(.a(s_59), .b(gate863inter3), .O(gate863inter10));
  nor2  gate1298(.a(gate863inter10), .b(gate863inter9), .O(gate863inter11));
  nor2  gate1299(.a(gate863inter11), .b(gate863inter6), .O(gate863inter12));
  nand2 gate1300(.a(gate863inter12), .b(gate863inter1), .O(N2878));
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );

  xor2  gate1791(.a(N2872), .b(N682), .O(gate866inter0));
  nand2 gate1792(.a(gate866inter0), .b(s_130), .O(gate866inter1));
  and2  gate1793(.a(N2872), .b(N682), .O(gate866inter2));
  inv1  gate1794(.a(s_130), .O(gate866inter3));
  inv1  gate1795(.a(s_131), .O(gate866inter4));
  nand2 gate1796(.a(gate866inter4), .b(gate866inter3), .O(gate866inter5));
  nor2  gate1797(.a(gate866inter5), .b(gate866inter2), .O(gate866inter6));
  inv1  gate1798(.a(N682), .O(gate866inter7));
  inv1  gate1799(.a(N2872), .O(gate866inter8));
  nand2 gate1800(.a(gate866inter8), .b(gate866inter7), .O(gate866inter9));
  nand2 gate1801(.a(s_131), .b(gate866inter3), .O(gate866inter10));
  nor2  gate1802(.a(gate866inter10), .b(gate866inter9), .O(gate866inter11));
  nor2  gate1803(.a(gate866inter11), .b(gate866inter6), .O(gate866inter12));
  nand2 gate1804(.a(gate866inter12), .b(gate866inter1), .O(N2881));
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );

  xor2  gate1931(.a(N2882), .b(N2873), .O(gate875inter0));
  nand2 gate1932(.a(gate875inter0), .b(s_150), .O(gate875inter1));
  and2  gate1933(.a(N2882), .b(N2873), .O(gate875inter2));
  inv1  gate1934(.a(s_150), .O(gate875inter3));
  inv1  gate1935(.a(s_151), .O(gate875inter4));
  nand2 gate1936(.a(gate875inter4), .b(gate875inter3), .O(gate875inter5));
  nor2  gate1937(.a(gate875inter5), .b(gate875inter2), .O(gate875inter6));
  inv1  gate1938(.a(N2873), .O(gate875inter7));
  inv1  gate1939(.a(N2882), .O(gate875inter8));
  nand2 gate1940(.a(gate875inter8), .b(gate875inter7), .O(gate875inter9));
  nand2 gate1941(.a(s_151), .b(gate875inter3), .O(gate875inter10));
  nor2  gate1942(.a(gate875inter10), .b(gate875inter9), .O(gate875inter11));
  nor2  gate1943(.a(gate875inter11), .b(gate875inter6), .O(gate875inter12));
  nand2 gate1944(.a(gate875inter12), .b(gate875inter1), .O(N2892));

  xor2  gate909(.a(N1461), .b(N2883), .O(gate876inter0));
  nand2 gate910(.a(gate876inter0), .b(s_4), .O(gate876inter1));
  and2  gate911(.a(N1461), .b(N2883), .O(gate876inter2));
  inv1  gate912(.a(s_4), .O(gate876inter3));
  inv1  gate913(.a(s_5), .O(gate876inter4));
  nand2 gate914(.a(gate876inter4), .b(gate876inter3), .O(gate876inter5));
  nor2  gate915(.a(gate876inter5), .b(gate876inter2), .O(gate876inter6));
  inv1  gate916(.a(N2883), .O(gate876inter7));
  inv1  gate917(.a(N1461), .O(gate876inter8));
  nand2 gate918(.a(gate876inter8), .b(gate876inter7), .O(gate876inter9));
  nand2 gate919(.a(s_5), .b(gate876inter3), .O(gate876inter10));
  nor2  gate920(.a(gate876inter10), .b(gate876inter9), .O(gate876inter11));
  nor2  gate921(.a(gate876inter11), .b(gate876inter6), .O(gate876inter12));
  nand2 gate922(.a(gate876inter12), .b(gate876inter1), .O(N2895));
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );

  xor2  gate2491(.a(N2897), .b(N2895), .O(gate879inter0));
  nand2 gate2492(.a(gate879inter0), .b(s_230), .O(gate879inter1));
  and2  gate2493(.a(N2897), .b(N2895), .O(gate879inter2));
  inv1  gate2494(.a(s_230), .O(gate879inter3));
  inv1  gate2495(.a(s_231), .O(gate879inter4));
  nand2 gate2496(.a(gate879inter4), .b(gate879inter3), .O(gate879inter5));
  nor2  gate2497(.a(gate879inter5), .b(gate879inter2), .O(gate879inter6));
  inv1  gate2498(.a(N2895), .O(gate879inter7));
  inv1  gate2499(.a(N2897), .O(gate879inter8));
  nand2 gate2500(.a(gate879inter8), .b(gate879inter7), .O(gate879inter9));
  nand2 gate2501(.a(s_231), .b(gate879inter3), .O(gate879inter10));
  nor2  gate2502(.a(gate879inter10), .b(gate879inter9), .O(gate879inter11));
  nor2  gate2503(.a(gate879inter11), .b(gate879inter6), .O(gate879inter12));
  nand2 gate2504(.a(gate879inter12), .b(gate879inter1), .O(N2898));
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule