module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12;


  xor2  gate455(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate456(.a(gate1inter0), .b(s_36), .O(gate1inter1));
  and2  gate457(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate458(.a(s_36), .O(gate1inter3));
  inv1  gate459(.a(s_37), .O(gate1inter4));
  nand2 gate460(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate461(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate462(.a(N1), .O(gate1inter7));
  inv1  gate463(.a(N5), .O(gate1inter8));
  nand2 gate464(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate465(.a(s_37), .b(gate1inter3), .O(gate1inter10));
  nor2  gate466(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate467(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate468(.a(gate1inter12), .b(gate1inter1), .O(N250));
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate343(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate344(.a(gate3inter0), .b(s_20), .O(gate3inter1));
  and2  gate345(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate346(.a(s_20), .O(gate3inter3));
  inv1  gate347(.a(s_21), .O(gate3inter4));
  nand2 gate348(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate349(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate350(.a(N17), .O(gate3inter7));
  inv1  gate351(.a(N21), .O(gate3inter8));
  nand2 gate352(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate353(.a(s_21), .b(gate3inter3), .O(gate3inter10));
  nor2  gate354(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate355(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate356(.a(gate3inter12), .b(gate3inter1), .O(N252));

  xor2  gate231(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate232(.a(gate4inter0), .b(s_4), .O(gate4inter1));
  and2  gate233(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate234(.a(s_4), .O(gate4inter3));
  inv1  gate235(.a(s_5), .O(gate4inter4));
  nand2 gate236(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate237(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate238(.a(N25), .O(gate4inter7));
  inv1  gate239(.a(N29), .O(gate4inter8));
  nand2 gate240(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate241(.a(s_5), .b(gate4inter3), .O(gate4inter10));
  nor2  gate242(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate243(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate244(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate273(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate274(.a(gate6inter0), .b(s_10), .O(gate6inter1));
  and2  gate275(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate276(.a(s_10), .O(gate6inter3));
  inv1  gate277(.a(s_11), .O(gate6inter4));
  nand2 gate278(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate279(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate280(.a(N41), .O(gate6inter7));
  inv1  gate281(.a(N45), .O(gate6inter8));
  nand2 gate282(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate283(.a(s_11), .b(gate6inter3), .O(gate6inter10));
  nor2  gate284(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate285(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate286(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );

  xor2  gate385(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate386(.a(gate10inter0), .b(s_26), .O(gate10inter1));
  and2  gate387(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate388(.a(s_26), .O(gate10inter3));
  inv1  gate389(.a(s_27), .O(gate10inter4));
  nand2 gate390(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate391(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate392(.a(N73), .O(gate10inter7));
  inv1  gate393(.a(N77), .O(gate10inter8));
  nand2 gate394(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate395(.a(s_27), .b(gate10inter3), .O(gate10inter10));
  nor2  gate396(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate397(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate398(.a(gate10inter12), .b(gate10inter1), .O(N259));
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );

  xor2  gate609(.a(N21), .b(N5), .O(gate27inter0));
  nand2 gate610(.a(gate27inter0), .b(s_58), .O(gate27inter1));
  and2  gate611(.a(N21), .b(N5), .O(gate27inter2));
  inv1  gate612(.a(s_58), .O(gate27inter3));
  inv1  gate613(.a(s_59), .O(gate27inter4));
  nand2 gate614(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate615(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate616(.a(N5), .O(gate27inter7));
  inv1  gate617(.a(N21), .O(gate27inter8));
  nand2 gate618(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate619(.a(s_59), .b(gate27inter3), .O(gate27inter10));
  nor2  gate620(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate621(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate622(.a(gate27inter12), .b(gate27inter1), .O(N276));

  xor2  gate539(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate540(.a(gate28inter0), .b(s_48), .O(gate28inter1));
  and2  gate541(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate542(.a(s_48), .O(gate28inter3));
  inv1  gate543(.a(s_49), .O(gate28inter4));
  nand2 gate544(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate545(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate546(.a(N37), .O(gate28inter7));
  inv1  gate547(.a(N53), .O(gate28inter8));
  nand2 gate548(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate549(.a(s_49), .b(gate28inter3), .O(gate28inter10));
  nor2  gate550(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate551(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate552(.a(gate28inter12), .b(gate28inter1), .O(N277));

  xor2  gate329(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate330(.a(gate29inter0), .b(s_18), .O(gate29inter1));
  and2  gate331(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate332(.a(s_18), .O(gate29inter3));
  inv1  gate333(.a(s_19), .O(gate29inter4));
  nand2 gate334(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate335(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate336(.a(N9), .O(gate29inter7));
  inv1  gate337(.a(N25), .O(gate29inter8));
  nand2 gate338(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate339(.a(s_19), .b(gate29inter3), .O(gate29inter10));
  nor2  gate340(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate341(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate342(.a(gate29inter12), .b(gate29inter1), .O(N278));
xor2 gate30( .a(N41), .b(N57), .O(N279) );

  xor2  gate581(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate582(.a(gate31inter0), .b(s_54), .O(gate31inter1));
  and2  gate583(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate584(.a(s_54), .O(gate31inter3));
  inv1  gate585(.a(s_55), .O(gate31inter4));
  nand2 gate586(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate587(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate588(.a(N13), .O(gate31inter7));
  inv1  gate589(.a(N29), .O(gate31inter8));
  nand2 gate590(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate591(.a(s_55), .b(gate31inter3), .O(gate31inter10));
  nor2  gate592(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate593(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate594(.a(gate31inter12), .b(gate31inter1), .O(N280));
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );

  xor2  gate301(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate302(.a(gate34inter0), .b(s_14), .O(gate34inter1));
  and2  gate303(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate304(.a(s_14), .O(gate34inter3));
  inv1  gate305(.a(s_15), .O(gate34inter4));
  nand2 gate306(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate307(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate308(.a(N97), .O(gate34inter7));
  inv1  gate309(.a(N113), .O(gate34inter8));
  nand2 gate310(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate311(.a(s_15), .b(gate34inter3), .O(gate34inter10));
  nor2  gate312(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate313(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate314(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );

  xor2  gate441(.a(N93), .b(N77), .O(gate39inter0));
  nand2 gate442(.a(gate39inter0), .b(s_34), .O(gate39inter1));
  and2  gate443(.a(N93), .b(N77), .O(gate39inter2));
  inv1  gate444(.a(s_34), .O(gate39inter3));
  inv1  gate445(.a(s_35), .O(gate39inter4));
  nand2 gate446(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate447(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate448(.a(N77), .O(gate39inter7));
  inv1  gate449(.a(N93), .O(gate39inter8));
  nand2 gate450(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate451(.a(s_35), .b(gate39inter3), .O(gate39inter10));
  nor2  gate452(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate453(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate454(.a(gate39inter12), .b(gate39inter1), .O(N288));
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );

  xor2  gate399(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate400(.a(gate43inter0), .b(s_28), .O(gate43inter1));
  and2  gate401(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate402(.a(s_28), .O(gate43inter3));
  inv1  gate403(.a(s_29), .O(gate43inter4));
  nand2 gate404(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate405(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate406(.a(N254), .O(gate43inter7));
  inv1  gate407(.a(N255), .O(gate43inter8));
  nand2 gate408(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate409(.a(s_29), .b(gate43inter3), .O(gate43inter10));
  nor2  gate410(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate411(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate412(.a(gate43inter12), .b(gate43inter1), .O(N296));
xor2 gate44( .a(N256), .b(N257), .O(N299) );

  xor2  gate469(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate470(.a(gate45inter0), .b(s_38), .O(gate45inter1));
  and2  gate471(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate472(.a(s_38), .O(gate45inter3));
  inv1  gate473(.a(s_39), .O(gate45inter4));
  nand2 gate474(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate475(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate476(.a(N258), .O(gate45inter7));
  inv1  gate477(.a(N259), .O(gate45inter8));
  nand2 gate478(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate479(.a(s_39), .b(gate45inter3), .O(gate45inter10));
  nor2  gate480(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate481(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate482(.a(gate45inter12), .b(gate45inter1), .O(N302));

  xor2  gate427(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate428(.a(gate46inter0), .b(s_32), .O(gate46inter1));
  and2  gate429(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate430(.a(s_32), .O(gate46inter3));
  inv1  gate431(.a(s_33), .O(gate46inter4));
  nand2 gate432(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate433(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate434(.a(N260), .O(gate46inter7));
  inv1  gate435(.a(N261), .O(gate46inter8));
  nand2 gate436(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate437(.a(s_33), .b(gate46inter3), .O(gate46inter10));
  nor2  gate438(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate439(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate440(.a(gate46inter12), .b(gate46inter1), .O(N305));
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );

  xor2  gate623(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate624(.a(gate49inter0), .b(s_60), .O(gate49inter1));
  and2  gate625(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate626(.a(s_60), .O(gate49inter3));
  inv1  gate627(.a(s_61), .O(gate49inter4));
  nand2 gate628(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate629(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate630(.a(N274), .O(gate49inter7));
  inv1  gate631(.a(N275), .O(gate49inter8));
  nand2 gate632(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate633(.a(s_61), .b(gate49inter3), .O(gate49inter10));
  nor2  gate634(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate635(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate636(.a(gate49inter12), .b(gate49inter1), .O(N314));
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );

  xor2  gate525(.a(N281), .b(N280), .O(gate52inter0));
  nand2 gate526(.a(gate52inter0), .b(s_46), .O(gate52inter1));
  and2  gate527(.a(N281), .b(N280), .O(gate52inter2));
  inv1  gate528(.a(s_46), .O(gate52inter3));
  inv1  gate529(.a(s_47), .O(gate52inter4));
  nand2 gate530(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate531(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate532(.a(N280), .O(gate52inter7));
  inv1  gate533(.a(N281), .O(gate52inter8));
  nand2 gate534(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate535(.a(s_47), .b(gate52inter3), .O(gate52inter10));
  nor2  gate536(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate537(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate538(.a(gate52inter12), .b(gate52inter1), .O(N317));

  xor2  gate357(.a(N283), .b(N282), .O(gate53inter0));
  nand2 gate358(.a(gate53inter0), .b(s_22), .O(gate53inter1));
  and2  gate359(.a(N283), .b(N282), .O(gate53inter2));
  inv1  gate360(.a(s_22), .O(gate53inter3));
  inv1  gate361(.a(s_23), .O(gate53inter4));
  nand2 gate362(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate363(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate364(.a(N282), .O(gate53inter7));
  inv1  gate365(.a(N283), .O(gate53inter8));
  nand2 gate366(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate367(.a(s_23), .b(gate53inter3), .O(gate53inter10));
  nor2  gate368(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate369(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate370(.a(gate53inter12), .b(gate53inter1), .O(N318));
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );

  xor2  gate595(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate596(.a(gate57inter0), .b(s_56), .O(gate57inter1));
  and2  gate597(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate598(.a(s_56), .O(gate57inter3));
  inv1  gate599(.a(s_57), .O(gate57inter4));
  nand2 gate600(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate601(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate602(.a(N290), .O(gate57inter7));
  inv1  gate603(.a(N293), .O(gate57inter8));
  nand2 gate604(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate605(.a(s_57), .b(gate57inter3), .O(gate57inter10));
  nor2  gate606(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate607(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate608(.a(gate57inter12), .b(gate57inter1), .O(N338));
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate497(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate498(.a(gate59inter0), .b(s_42), .O(gate59inter1));
  and2  gate499(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate500(.a(s_42), .O(gate59inter3));
  inv1  gate501(.a(s_43), .O(gate59inter4));
  nand2 gate502(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate503(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate504(.a(N290), .O(gate59inter7));
  inv1  gate505(.a(N296), .O(gate59inter8));
  nand2 gate506(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate507(.a(s_43), .b(gate59inter3), .O(gate59inter10));
  nor2  gate508(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate509(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate510(.a(gate59inter12), .b(gate59inter1), .O(N340));
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );

  xor2  gate259(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate260(.a(gate64inter0), .b(s_8), .O(gate64inter1));
  and2  gate261(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate262(.a(s_8), .O(gate64inter3));
  inv1  gate263(.a(s_9), .O(gate64inter4));
  nand2 gate264(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate265(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate266(.a(N305), .O(gate64inter7));
  inv1  gate267(.a(N311), .O(gate64inter8));
  nand2 gate268(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate269(.a(s_9), .b(gate64inter3), .O(gate64inter10));
  nor2  gate270(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate271(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate272(.a(gate64inter12), .b(gate64inter1), .O(N345));
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );

  xor2  gate315(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate316(.a(gate73inter0), .b(s_16), .O(gate73inter1));
  and2  gate317(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate318(.a(s_16), .O(gate73inter3));
  inv1  gate319(.a(s_17), .O(gate73inter4));
  nand2 gate320(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate321(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate322(.a(N314), .O(gate73inter7));
  inv1  gate323(.a(N346), .O(gate73inter8));
  nand2 gate324(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate325(.a(s_17), .b(gate73inter3), .O(gate73inter10));
  nor2  gate326(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate327(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate328(.a(gate73inter12), .b(gate73inter1), .O(N354));
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate511(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate512(.a(gate176inter0), .b(s_44), .O(gate176inter1));
  and2  gate513(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate514(.a(s_44), .O(gate176inter3));
  inv1  gate515(.a(s_45), .O(gate176inter4));
  nand2 gate516(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate517(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate518(.a(N21), .O(gate176inter7));
  inv1  gate519(.a(N697), .O(gate176inter8));
  nand2 gate520(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate521(.a(s_45), .b(gate176inter3), .O(gate176inter10));
  nor2  gate522(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate523(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate524(.a(gate176inter12), .b(gate176inter1), .O(N729));

  xor2  gate553(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate554(.a(gate177inter0), .b(s_50), .O(gate177inter1));
  and2  gate555(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate556(.a(s_50), .O(gate177inter3));
  inv1  gate557(.a(s_51), .O(gate177inter4));
  nand2 gate558(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate559(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate560(.a(N25), .O(gate177inter7));
  inv1  gate561(.a(N698), .O(gate177inter8));
  nand2 gate562(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate563(.a(s_51), .b(gate177inter3), .O(gate177inter10));
  nor2  gate564(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate565(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate566(.a(gate177inter12), .b(gate177inter1), .O(N730));

  xor2  gate567(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate568(.a(gate178inter0), .b(s_52), .O(gate178inter1));
  and2  gate569(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate570(.a(s_52), .O(gate178inter3));
  inv1  gate571(.a(s_53), .O(gate178inter4));
  nand2 gate572(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate573(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate574(.a(N29), .O(gate178inter7));
  inv1  gate575(.a(N699), .O(gate178inter8));
  nand2 gate576(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate577(.a(s_53), .b(gate178inter3), .O(gate178inter10));
  nor2  gate578(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate579(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate580(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );

  xor2  gate287(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate288(.a(gate182inter0), .b(s_12), .O(gate182inter1));
  and2  gate289(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate290(.a(s_12), .O(gate182inter3));
  inv1  gate291(.a(s_13), .O(gate182inter4));
  nand2 gate292(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate293(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate294(.a(N45), .O(gate182inter7));
  inv1  gate295(.a(N703), .O(gate182inter8));
  nand2 gate296(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate297(.a(s_13), .b(gate182inter3), .O(gate182inter10));
  nor2  gate298(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate299(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate300(.a(gate182inter12), .b(gate182inter1), .O(N735));
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );

  xor2  gate413(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate414(.a(gate191inter0), .b(s_30), .O(gate191inter1));
  and2  gate415(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate416(.a(s_30), .O(gate191inter3));
  inv1  gate417(.a(s_31), .O(gate191inter4));
  nand2 gate418(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate419(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate420(.a(N81), .O(gate191inter7));
  inv1  gate421(.a(N712), .O(gate191inter8));
  nand2 gate422(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate423(.a(s_31), .b(gate191inter3), .O(gate191inter10));
  nor2  gate424(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate425(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate426(.a(gate191inter12), .b(gate191inter1), .O(N744));

  xor2  gate203(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate204(.a(gate192inter0), .b(s_0), .O(gate192inter1));
  and2  gate205(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate206(.a(s_0), .O(gate192inter3));
  inv1  gate207(.a(s_1), .O(gate192inter4));
  nand2 gate208(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate209(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate210(.a(N85), .O(gate192inter7));
  inv1  gate211(.a(N713), .O(gate192inter8));
  nand2 gate212(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate213(.a(s_1), .b(gate192inter3), .O(gate192inter10));
  nor2  gate214(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate215(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate216(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );

  xor2  gate245(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate246(.a(gate195inter0), .b(s_6), .O(gate195inter1));
  and2  gate247(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate248(.a(s_6), .O(gate195inter3));
  inv1  gate249(.a(s_7), .O(gate195inter4));
  nand2 gate250(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate251(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate252(.a(N97), .O(gate195inter7));
  inv1  gate253(.a(N716), .O(gate195inter8));
  nand2 gate254(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate255(.a(s_7), .b(gate195inter3), .O(gate195inter10));
  nor2  gate256(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate257(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate258(.a(gate195inter12), .b(gate195inter1), .O(N748));
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );

  xor2  gate371(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate372(.a(gate199inter0), .b(s_24), .O(gate199inter1));
  and2  gate373(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate374(.a(s_24), .O(gate199inter3));
  inv1  gate375(.a(s_25), .O(gate199inter4));
  nand2 gate376(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate377(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate378(.a(N113), .O(gate199inter7));
  inv1  gate379(.a(N720), .O(gate199inter8));
  nand2 gate380(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate381(.a(s_25), .b(gate199inter3), .O(gate199inter10));
  nor2  gate382(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate383(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate384(.a(gate199inter12), .b(gate199inter1), .O(N752));
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate483(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate484(.a(gate201inter0), .b(s_40), .O(gate201inter1));
  and2  gate485(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate486(.a(s_40), .O(gate201inter3));
  inv1  gate487(.a(s_41), .O(gate201inter4));
  nand2 gate488(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate489(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate490(.a(N121), .O(gate201inter7));
  inv1  gate491(.a(N722), .O(gate201inter8));
  nand2 gate492(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate493(.a(s_41), .b(gate201inter3), .O(gate201inter10));
  nor2  gate494(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate495(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate496(.a(gate201inter12), .b(gate201inter1), .O(N754));

  xor2  gate217(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate218(.a(gate202inter0), .b(s_2), .O(gate202inter1));
  and2  gate219(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate220(.a(s_2), .O(gate202inter3));
  inv1  gate221(.a(s_3), .O(gate202inter4));
  nand2 gate222(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate223(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate224(.a(N125), .O(gate202inter7));
  inv1  gate225(.a(N723), .O(gate202inter8));
  nand2 gate226(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate227(.a(s_3), .b(gate202inter3), .O(gate202inter10));
  nor2  gate228(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate229(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate230(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule