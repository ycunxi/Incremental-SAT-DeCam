module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate378inter0, gate378inter1, gate378inter2, gate378inter3, gate378inter4, gate378inter5, gate378inter6, gate378inter7, gate378inter8, gate378inter9, gate378inter10, gate378inter11, gate378inter12, gate552inter0, gate552inter1, gate552inter2, gate552inter3, gate552inter4, gate552inter5, gate552inter6, gate552inter7, gate552inter8, gate552inter9, gate552inter10, gate552inter11, gate552inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate650inter0, gate650inter1, gate650inter2, gate650inter3, gate650inter4, gate650inter5, gate650inter6, gate650inter7, gate650inter8, gate650inter9, gate650inter10, gate650inter11, gate650inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate613inter0, gate613inter1, gate613inter2, gate613inter3, gate613inter4, gate613inter5, gate613inter6, gate613inter7, gate613inter8, gate613inter9, gate613inter10, gate613inter11, gate613inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate879inter0, gate879inter1, gate879inter2, gate879inter3, gate879inter4, gate879inter5, gate879inter6, gate879inter7, gate879inter8, gate879inter9, gate879inter10, gate879inter11, gate879inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate338inter0, gate338inter1, gate338inter2, gate338inter3, gate338inter4, gate338inter5, gate338inter6, gate338inter7, gate338inter8, gate338inter9, gate338inter10, gate338inter11, gate338inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate530inter0, gate530inter1, gate530inter2, gate530inter3, gate530inter4, gate530inter5, gate530inter6, gate530inter7, gate530inter8, gate530inter9, gate530inter10, gate530inter11, gate530inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12, gate366inter0, gate366inter1, gate366inter2, gate366inter3, gate366inter4, gate366inter5, gate366inter6, gate366inter7, gate366inter8, gate366inter9, gate366inter10, gate366inter11, gate366inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate758inter0, gate758inter1, gate758inter2, gate758inter3, gate758inter4, gate758inter5, gate758inter6, gate758inter7, gate758inter8, gate758inter9, gate758inter10, gate758inter11, gate758inter12, gate876inter0, gate876inter1, gate876inter2, gate876inter3, gate876inter4, gate876inter5, gate876inter6, gate876inter7, gate876inter8, gate876inter9, gate876inter10, gate876inter11, gate876inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate357inter0, gate357inter1, gate357inter2, gate357inter3, gate357inter4, gate357inter5, gate357inter6, gate357inter7, gate357inter8, gate357inter9, gate357inter10, gate357inter11, gate357inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate769inter0, gate769inter1, gate769inter2, gate769inter3, gate769inter4, gate769inter5, gate769inter6, gate769inter7, gate769inter8, gate769inter9, gate769inter10, gate769inter11, gate769inter12, gate632inter0, gate632inter1, gate632inter2, gate632inter3, gate632inter4, gate632inter5, gate632inter6, gate632inter7, gate632inter8, gate632inter9, gate632inter10, gate632inter11, gate632inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate1357(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate1358(.a(gate96inter0), .b(s_68), .O(gate96inter1));
  and2  gate1359(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate1360(.a(s_68), .O(gate96inter3));
  inv1  gate1361(.a(s_69), .O(gate96inter4));
  nand2 gate1362(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1363(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1364(.a(N326), .O(gate96inter7));
  inv1  gate1365(.a(N277), .O(gate96inter8));
  nand2 gate1366(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1367(.a(s_69), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1368(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1369(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1370(.a(gate96inter12), .b(gate96inter1), .O(N601));
nand2 gate97( .a(N326), .b(N280), .O(N602) );

  xor2  gate1105(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate1106(.a(gate98inter0), .b(s_32), .O(gate98inter1));
  and2  gate1107(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate1108(.a(s_32), .O(gate98inter3));
  inv1  gate1109(.a(s_33), .O(gate98inter4));
  nand2 gate1110(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1111(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1112(.a(N260), .O(gate98inter7));
  inv1  gate1113(.a(N72), .O(gate98inter8));
  nand2 gate1114(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1115(.a(s_33), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1116(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1117(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1118(.a(gate98inter12), .b(gate98inter1), .O(N603));

  xor2  gate1189(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate1190(.a(gate99inter0), .b(s_44), .O(gate99inter1));
  and2  gate1191(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate1192(.a(s_44), .O(gate99inter3));
  inv1  gate1193(.a(s_45), .O(gate99inter4));
  nand2 gate1194(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1195(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1196(.a(N260), .O(gate99inter7));
  inv1  gate1197(.a(N300), .O(gate99inter8));
  nand2 gate1198(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1199(.a(s_45), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1200(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1201(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1202(.a(gate99inter12), .b(gate99inter1), .O(N608));
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );

  xor2  gate1371(.a(N1002), .b(N739), .O(gate243inter0));
  nand2 gate1372(.a(gate243inter0), .b(s_70), .O(gate243inter1));
  and2  gate1373(.a(N1002), .b(N739), .O(gate243inter2));
  inv1  gate1374(.a(s_70), .O(gate243inter3));
  inv1  gate1375(.a(s_71), .O(gate243inter4));
  nand2 gate1376(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1377(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1378(.a(N739), .O(gate243inter7));
  inv1  gate1379(.a(N1002), .O(gate243inter8));
  nand2 gate1380(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1381(.a(s_71), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1382(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1383(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1384(.a(gate243inter12), .b(gate243inter1), .O(N1128));
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );

  xor2  gate1077(.a(N1008), .b(N751), .O(gate247inter0));
  nand2 gate1078(.a(gate247inter0), .b(s_28), .O(gate247inter1));
  and2  gate1079(.a(N1008), .b(N751), .O(gate247inter2));
  inv1  gate1080(.a(s_28), .O(gate247inter3));
  inv1  gate1081(.a(s_29), .O(gate247inter4));
  nand2 gate1082(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1083(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1084(.a(N751), .O(gate247inter7));
  inv1  gate1085(.a(N1008), .O(gate247inter8));
  nand2 gate1086(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1087(.a(s_29), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1088(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1089(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1090(.a(gate247inter12), .b(gate247inter1), .O(N1132));
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );

  xor2  gate1049(.a(N1068), .b(N1067), .O(gate263inter0));
  nand2 gate1050(.a(gate263inter0), .b(s_24), .O(gate263inter1));
  and2  gate1051(.a(N1068), .b(N1067), .O(gate263inter2));
  inv1  gate1052(.a(s_24), .O(gate263inter3));
  inv1  gate1053(.a(s_25), .O(gate263inter4));
  nand2 gate1054(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1055(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1056(.a(N1067), .O(gate263inter7));
  inv1  gate1057(.a(N1068), .O(gate263inter8));
  nand2 gate1058(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1059(.a(s_25), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1060(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1061(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1062(.a(gate263inter12), .b(gate263inter1), .O(N1162));
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );

  xor2  gate1315(.a(N938), .b(N1010), .O(gate271inter0));
  nand2 gate1316(.a(gate271inter0), .b(s_62), .O(gate271inter1));
  and2  gate1317(.a(N938), .b(N1010), .O(gate271inter2));
  inv1  gate1318(.a(s_62), .O(gate271inter3));
  inv1  gate1319(.a(s_63), .O(gate271inter4));
  nand2 gate1320(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1321(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1322(.a(N1010), .O(gate271inter7));
  inv1  gate1323(.a(N938), .O(gate271inter8));
  nand2 gate1324(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1325(.a(s_63), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1326(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1327(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1328(.a(gate271inter12), .b(gate271inter1), .O(N1206));
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );

  xor2  gate1133(.a(N968), .b(N1034), .O(gate286inter0));
  nand2 gate1134(.a(gate286inter0), .b(s_36), .O(gate286inter1));
  and2  gate1135(.a(N968), .b(N1034), .O(gate286inter2));
  inv1  gate1136(.a(s_36), .O(gate286inter3));
  inv1  gate1137(.a(s_37), .O(gate286inter4));
  nand2 gate1138(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1139(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1140(.a(N1034), .O(gate286inter7));
  inv1  gate1141(.a(N968), .O(gate286inter8));
  nand2 gate1142(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1143(.a(s_37), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1144(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1145(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1146(.a(gate286inter12), .b(gate286inter1), .O(N1221));
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );

  xor2  gate881(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate882(.a(gate298inter0), .b(s_0), .O(gate298inter1));
  and2  gate883(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate884(.a(s_0), .O(gate298inter3));
  inv1  gate885(.a(s_1), .O(gate298inter4));
  nand2 gate886(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate887(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate888(.a(N1121), .O(gate298inter7));
  inv1  gate889(.a(N1122), .O(gate298inter8));
  nand2 gate890(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate891(.a(s_1), .b(gate298inter3), .O(gate298inter10));
  nor2  gate892(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate893(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate894(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );

  xor2  gate1063(.a(N1207), .b(N691), .O(gate314inter0));
  nand2 gate1064(.a(gate314inter0), .b(s_26), .O(gate314inter1));
  and2  gate1065(.a(N1207), .b(N691), .O(gate314inter2));
  inv1  gate1066(.a(s_26), .O(gate314inter3));
  inv1  gate1067(.a(s_27), .O(gate314inter4));
  nand2 gate1068(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate1069(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate1070(.a(N691), .O(gate314inter7));
  inv1  gate1071(.a(N1207), .O(gate314inter8));
  nand2 gate1072(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate1073(.a(s_27), .b(gate314inter3), .O(gate314inter10));
  nor2  gate1074(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate1075(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate1076(.a(gate314inter12), .b(gate314inter1), .O(N1310));
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );

  xor2  gate1021(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate1022(.a(gate316inter0), .b(s_20), .O(gate316inter1));
  and2  gate1023(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate1024(.a(s_20), .O(gate316inter3));
  inv1  gate1025(.a(s_21), .O(gate316inter4));
  nand2 gate1026(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate1027(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate1028(.a(N697), .O(gate316inter7));
  inv1  gate1029(.a(N1211), .O(gate316inter8));
  nand2 gate1030(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate1031(.a(s_21), .b(gate316inter3), .O(gate316inter10));
  nor2  gate1032(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate1033(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate1034(.a(gate316inter12), .b(gate316inter1), .O(N1312));
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );

  xor2  gate965(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate966(.a(gate326inter0), .b(s_12), .O(gate326inter1));
  and2  gate967(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate968(.a(s_12), .O(gate326inter3));
  inv1  gate969(.a(s_13), .O(gate326inter4));
  nand2 gate970(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate971(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate972(.a(N733), .O(gate326inter7));
  inv1  gate973(.a(N1241), .O(gate326inter8));
  nand2 gate974(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate975(.a(s_13), .b(gate326inter3), .O(gate326inter10));
  nor2  gate976(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate977(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate978(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );

  xor2  gate1147(.a(N1212), .b(N1312), .O(gate338inter0));
  nand2 gate1148(.a(gate338inter0), .b(s_38), .O(gate338inter1));
  and2  gate1149(.a(N1212), .b(N1312), .O(gate338inter2));
  inv1  gate1150(.a(s_38), .O(gate338inter3));
  inv1  gate1151(.a(s_39), .O(gate338inter4));
  nand2 gate1152(.a(gate338inter4), .b(gate338inter3), .O(gate338inter5));
  nor2  gate1153(.a(gate338inter5), .b(gate338inter2), .O(gate338inter6));
  inv1  gate1154(.a(N1312), .O(gate338inter7));
  inv1  gate1155(.a(N1212), .O(gate338inter8));
  nand2 gate1156(.a(gate338inter8), .b(gate338inter7), .O(gate338inter9));
  nand2 gate1157(.a(s_39), .b(gate338inter3), .O(gate338inter10));
  nor2  gate1158(.a(gate338inter10), .b(gate338inter9), .O(gate338inter11));
  nor2  gate1159(.a(gate338inter11), .b(gate338inter6), .O(gate338inter12));
  nand2 gate1160(.a(gate338inter12), .b(gate338inter1), .O(N1361));
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );

  xor2  gate1343(.a(N1346), .b(N649), .O(gate357inter0));
  nand2 gate1344(.a(gate357inter0), .b(s_66), .O(gate357inter1));
  and2  gate1345(.a(N1346), .b(N649), .O(gate357inter2));
  inv1  gate1346(.a(s_66), .O(gate357inter3));
  inv1  gate1347(.a(s_67), .O(gate357inter4));
  nand2 gate1348(.a(gate357inter4), .b(gate357inter3), .O(gate357inter5));
  nor2  gate1349(.a(gate357inter5), .b(gate357inter2), .O(gate357inter6));
  inv1  gate1350(.a(N649), .O(gate357inter7));
  inv1  gate1351(.a(N1346), .O(gate357inter8));
  nand2 gate1352(.a(gate357inter8), .b(gate357inter7), .O(gate357inter9));
  nand2 gate1353(.a(s_67), .b(gate357inter3), .O(gate357inter10));
  nor2  gate1354(.a(gate357inter10), .b(gate357inter9), .O(gate357inter11));
  nor2  gate1355(.a(gate357inter11), .b(gate357inter6), .O(gate357inter12));
  nand2 gate1356(.a(gate357inter12), .b(gate357inter1), .O(N1412));
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );

  xor2  gate1245(.a(N1148), .b(N1355), .O(gate366inter0));
  nand2 gate1246(.a(gate366inter0), .b(s_52), .O(gate366inter1));
  and2  gate1247(.a(N1148), .b(N1355), .O(gate366inter2));
  inv1  gate1248(.a(s_52), .O(gate366inter3));
  inv1  gate1249(.a(s_53), .O(gate366inter4));
  nand2 gate1250(.a(gate366inter4), .b(gate366inter3), .O(gate366inter5));
  nor2  gate1251(.a(gate366inter5), .b(gate366inter2), .O(gate366inter6));
  inv1  gate1252(.a(N1355), .O(gate366inter7));
  inv1  gate1253(.a(N1148), .O(gate366inter8));
  nand2 gate1254(.a(gate366inter8), .b(gate366inter7), .O(gate366inter9));
  nand2 gate1255(.a(s_53), .b(gate366inter3), .O(gate366inter10));
  nor2  gate1256(.a(gate366inter10), .b(gate366inter9), .O(gate366inter11));
  nor2  gate1257(.a(gate366inter11), .b(gate366inter6), .O(gate366inter12));
  nand2 gate1258(.a(gate366inter12), .b(gate366inter1), .O(N1443));
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );

  xor2  gate909(.a(N1156), .b(N1373), .O(gate378inter0));
  nand2 gate910(.a(gate378inter0), .b(s_4), .O(gate378inter1));
  and2  gate911(.a(N1156), .b(N1373), .O(gate378inter2));
  inv1  gate912(.a(s_4), .O(gate378inter3));
  inv1  gate913(.a(s_5), .O(gate378inter4));
  nand2 gate914(.a(gate378inter4), .b(gate378inter3), .O(gate378inter5));
  nor2  gate915(.a(gate378inter5), .b(gate378inter2), .O(gate378inter6));
  inv1  gate916(.a(N1373), .O(gate378inter7));
  inv1  gate917(.a(N1156), .O(gate378inter8));
  nand2 gate918(.a(gate378inter8), .b(gate378inter7), .O(gate378inter9));
  nand2 gate919(.a(s_5), .b(gate378inter3), .O(gate378inter10));
  nor2  gate920(.a(gate378inter10), .b(gate378inter9), .O(gate378inter11));
  nor2  gate921(.a(gate378inter11), .b(gate378inter6), .O(gate378inter12));
  nand2 gate922(.a(gate378inter12), .b(gate378inter1), .O(N1457));
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );

  xor2  gate1329(.a(N1444), .b(N939), .O(gate396inter0));
  nand2 gate1330(.a(gate396inter0), .b(s_64), .O(gate396inter1));
  and2  gate1331(.a(N1444), .b(N939), .O(gate396inter2));
  inv1  gate1332(.a(s_64), .O(gate396inter3));
  inv1  gate1333(.a(s_65), .O(gate396inter4));
  nand2 gate1334(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1335(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1336(.a(N939), .O(gate396inter7));
  inv1  gate1337(.a(N1444), .O(gate396inter8));
  nand2 gate1338(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1339(.a(s_65), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1340(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1341(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1342(.a(gate396inter12), .b(gate396inter1), .O(N1487));
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );

  xor2  gate993(.a(N1496), .b(N1459), .O(gate419inter0));
  nand2 gate994(.a(gate419inter0), .b(s_16), .O(gate419inter1));
  and2  gate995(.a(N1496), .b(N1459), .O(gate419inter2));
  inv1  gate996(.a(s_16), .O(gate419inter3));
  inv1  gate997(.a(s_17), .O(gate419inter4));
  nand2 gate998(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate999(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1000(.a(N1459), .O(gate419inter7));
  inv1  gate1001(.a(N1496), .O(gate419inter8));
  nand2 gate1002(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1003(.a(s_17), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1004(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1005(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1006(.a(gate419inter12), .b(gate419inter1), .O(N1527));
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate937(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate938(.a(gate421inter0), .b(s_8), .O(gate421inter1));
  and2  gate939(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate940(.a(s_8), .O(gate421inter3));
  inv1  gate941(.a(s_9), .O(gate421inter4));
  nand2 gate942(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate943(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate944(.a(N1462), .O(gate421inter7));
  inv1  gate945(.a(N1498), .O(gate421inter8));
  nand2 gate946(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate947(.a(s_9), .b(gate421inter3), .O(gate421inter10));
  nor2  gate948(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate949(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate950(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );

  xor2  gate1091(.a(N1532), .b(N1481), .O(gate433inter0));
  nand2 gate1092(.a(gate433inter0), .b(s_30), .O(gate433inter1));
  and2  gate1093(.a(N1532), .b(N1481), .O(gate433inter2));
  inv1  gate1094(.a(s_30), .O(gate433inter3));
  inv1  gate1095(.a(s_31), .O(gate433inter4));
  nand2 gate1096(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1097(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1098(.a(N1481), .O(gate433inter7));
  inv1  gate1099(.a(N1532), .O(gate433inter8));
  nand2 gate1100(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1101(.a(s_31), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1102(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1103(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1104(.a(gate433inter12), .b(gate433inter1), .O(N1568));
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );

  xor2  gate1161(.a(N1747), .b(N1710), .O(gate511inter0));
  nand2 gate1162(.a(gate511inter0), .b(s_40), .O(gate511inter1));
  and2  gate1163(.a(N1747), .b(N1710), .O(gate511inter2));
  inv1  gate1164(.a(s_40), .O(gate511inter3));
  inv1  gate1165(.a(s_41), .O(gate511inter4));
  nand2 gate1166(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1167(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1168(.a(N1710), .O(gate511inter7));
  inv1  gate1169(.a(N1747), .O(gate511inter8));
  nand2 gate1170(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1171(.a(s_41), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1172(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1173(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1174(.a(gate511inter12), .b(gate511inter1), .O(N1777));
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );

  xor2  gate1203(.a(N1764), .b(N1792), .O(gate530inter0));
  nand2 gate1204(.a(gate530inter0), .b(s_46), .O(gate530inter1));
  and2  gate1205(.a(N1764), .b(N1792), .O(gate530inter2));
  inv1  gate1206(.a(s_46), .O(gate530inter3));
  inv1  gate1207(.a(s_47), .O(gate530inter4));
  nand2 gate1208(.a(gate530inter4), .b(gate530inter3), .O(gate530inter5));
  nor2  gate1209(.a(gate530inter5), .b(gate530inter2), .O(gate530inter6));
  inv1  gate1210(.a(N1792), .O(gate530inter7));
  inv1  gate1211(.a(N1764), .O(gate530inter8));
  nand2 gate1212(.a(gate530inter8), .b(gate530inter7), .O(gate530inter9));
  nand2 gate1213(.a(s_47), .b(gate530inter3), .O(gate530inter10));
  nor2  gate1214(.a(gate530inter10), .b(gate530inter9), .O(gate530inter11));
  nor2  gate1215(.a(gate530inter11), .b(gate530inter6), .O(gate530inter12));
  nand2 gate1216(.a(gate530inter12), .b(gate530inter1), .O(N1815));
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate951(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate952(.a(gate532inter0), .b(s_10), .O(gate532inter1));
  and2  gate953(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate954(.a(s_10), .O(gate532inter3));
  inv1  gate955(.a(s_11), .O(gate532inter4));
  nand2 gate956(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate957(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate958(.a(N1777), .O(gate532inter7));
  inv1  gate959(.a(N1490), .O(gate532inter8));
  nand2 gate960(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate961(.a(s_11), .b(gate532inter3), .O(gate532inter10));
  nor2  gate962(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate963(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate964(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );

  xor2  gate1217(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate1218(.a(gate547inter0), .b(s_48), .O(gate547inter1));
  and2  gate1219(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate1220(.a(s_48), .O(gate547inter3));
  inv1  gate1221(.a(s_49), .O(gate547inter4));
  nand2 gate1222(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate1223(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate1224(.a(N1815), .O(gate547inter7));
  inv1  gate1225(.a(N1707), .O(gate547inter8));
  nand2 gate1226(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate1227(.a(s_49), .b(gate547inter3), .O(gate547inter10));
  nor2  gate1228(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate1229(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate1230(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );

  xor2  gate923(.a(N1728), .b(N1812), .O(gate552inter0));
  nand2 gate924(.a(gate552inter0), .b(s_6), .O(gate552inter1));
  and2  gate925(.a(N1728), .b(N1812), .O(gate552inter2));
  inv1  gate926(.a(s_6), .O(gate552inter3));
  inv1  gate927(.a(s_7), .O(gate552inter4));
  nand2 gate928(.a(gate552inter4), .b(gate552inter3), .O(gate552inter5));
  nor2  gate929(.a(gate552inter5), .b(gate552inter2), .O(gate552inter6));
  inv1  gate930(.a(N1812), .O(gate552inter7));
  inv1  gate931(.a(N1728), .O(gate552inter8));
  nand2 gate932(.a(gate552inter8), .b(gate552inter7), .O(gate552inter9));
  nand2 gate933(.a(s_7), .b(gate552inter3), .O(gate552inter10));
  nor2  gate934(.a(gate552inter10), .b(gate552inter9), .O(gate552inter11));
  nor2  gate935(.a(gate552inter11), .b(gate552inter6), .O(gate552inter12));
  nand2 gate936(.a(gate552inter12), .b(gate552inter1), .O(N1865));
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );

  xor2  gate1399(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate1400(.a(gate562inter0), .b(s_74), .O(gate562inter1));
  and2  gate1401(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate1402(.a(s_74), .O(gate562inter3));
  inv1  gate1403(.a(s_75), .O(gate562inter4));
  nand2 gate1404(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate1405(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate1406(.a(N1643), .O(gate562inter7));
  inv1  gate1407(.a(N1856), .O(gate562inter8));
  nand2 gate1408(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate1409(.a(s_75), .b(gate562inter3), .O(gate562inter10));
  nor2  gate1410(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate1411(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate1412(.a(gate562inter12), .b(gate562inter1), .O(N1885));
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate1231(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate1232(.a(gate565inter0), .b(s_50), .O(gate565inter1));
  and2  gate1233(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate1234(.a(s_50), .O(gate565inter3));
  inv1  gate1235(.a(s_51), .O(gate565inter4));
  nand2 gate1236(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate1237(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate1238(.a(N1838), .O(gate565inter7));
  inv1  gate1239(.a(N1785), .O(gate565inter8));
  nand2 gate1240(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate1241(.a(s_51), .b(gate565inter3), .O(gate565inter10));
  nor2  gate1242(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate1243(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate1244(.a(gate565inter12), .b(gate565inter1), .O(N1896));
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate979(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate980(.a(gate612inter0), .b(s_14), .O(gate612inter1));
  and2  gate981(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate982(.a(s_14), .O(gate612inter3));
  inv1  gate983(.a(s_15), .O(gate612inter4));
  nand2 gate984(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate985(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate986(.a(N673), .O(gate612inter7));
  inv1  gate987(.a(N1976), .O(gate612inter8));
  nand2 gate988(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate989(.a(s_15), .b(gate612inter3), .O(gate612inter10));
  nor2  gate990(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate991(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate992(.a(gate612inter12), .b(gate612inter1), .O(N2008));

  xor2  gate1035(.a(N1978), .b(N670), .O(gate613inter0));
  nand2 gate1036(.a(gate613inter0), .b(s_22), .O(gate613inter1));
  and2  gate1037(.a(N1978), .b(N670), .O(gate613inter2));
  inv1  gate1038(.a(s_22), .O(gate613inter3));
  inv1  gate1039(.a(s_23), .O(gate613inter4));
  nand2 gate1040(.a(gate613inter4), .b(gate613inter3), .O(gate613inter5));
  nor2  gate1041(.a(gate613inter5), .b(gate613inter2), .O(gate613inter6));
  inv1  gate1042(.a(N670), .O(gate613inter7));
  inv1  gate1043(.a(N1978), .O(gate613inter8));
  nand2 gate1044(.a(gate613inter8), .b(gate613inter7), .O(gate613inter9));
  nand2 gate1045(.a(s_23), .b(gate613inter3), .O(gate613inter10));
  nor2  gate1046(.a(gate613inter10), .b(gate613inter9), .O(gate613inter11));
  nor2  gate1047(.a(gate613inter11), .b(gate613inter6), .O(gate613inter12));
  nand2 gate1048(.a(gate613inter12), .b(gate613inter1), .O(N2009));
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );

  xor2  gate1175(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate1176(.a(gate627inter0), .b(s_42), .O(gate627inter1));
  and2  gate1177(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate1178(.a(s_42), .O(gate627inter3));
  inv1  gate1179(.a(s_43), .O(gate627inter4));
  nand2 gate1180(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate1181(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate1182(.a(N1975), .O(gate627inter7));
  inv1  gate1183(.a(N2008), .O(gate627inter8));
  nand2 gate1184(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate1185(.a(s_43), .b(gate627inter3), .O(gate627inter10));
  nor2  gate1186(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate1187(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate1188(.a(gate627inter12), .b(gate627inter1), .O(N2026));
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );

  xor2  gate1441(.a(N2015), .b(N1571), .O(gate632inter0));
  nand2 gate1442(.a(gate632inter0), .b(s_80), .O(gate632inter1));
  and2  gate1443(.a(N2015), .b(N1571), .O(gate632inter2));
  inv1  gate1444(.a(s_80), .O(gate632inter3));
  inv1  gate1445(.a(s_81), .O(gate632inter4));
  nand2 gate1446(.a(gate632inter4), .b(gate632inter3), .O(gate632inter5));
  nor2  gate1447(.a(gate632inter5), .b(gate632inter2), .O(gate632inter6));
  inv1  gate1448(.a(N1571), .O(gate632inter7));
  inv1  gate1449(.a(N2015), .O(gate632inter8));
  nand2 gate1450(.a(gate632inter8), .b(gate632inter7), .O(gate632inter9));
  nand2 gate1451(.a(s_81), .b(gate632inter3), .O(gate632inter10));
  nor2  gate1452(.a(gate632inter10), .b(gate632inter9), .O(gate632inter11));
  nor2  gate1453(.a(gate632inter11), .b(gate632inter6), .O(gate632inter12));
  nand2 gate1454(.a(gate632inter12), .b(gate632inter1), .O(N2037));

  xor2  gate1385(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate1386(.a(gate633inter0), .b(s_72), .O(gate633inter1));
  and2  gate1387(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate1388(.a(s_72), .O(gate633inter3));
  inv1  gate1389(.a(s_73), .O(gate633inter4));
  nand2 gate1390(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate1391(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate1392(.a(N2020), .O(gate633inter7));
  inv1  gate1393(.a(N2000), .O(gate633inter8));
  nand2 gate1394(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate1395(.a(s_73), .b(gate633inter3), .O(gate633inter10));
  nor2  gate1396(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate1397(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate1398(.a(gate633inter12), .b(gate633inter1), .O(N2038));
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );

  xor2  gate1413(.a(N2003), .b(N2023), .O(gate635inter0));
  nand2 gate1414(.a(gate635inter0), .b(s_76), .O(gate635inter1));
  and2  gate1415(.a(N2003), .b(N2023), .O(gate635inter2));
  inv1  gate1416(.a(s_76), .O(gate635inter3));
  inv1  gate1417(.a(s_77), .O(gate635inter4));
  nand2 gate1418(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate1419(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate1420(.a(N2023), .O(gate635inter7));
  inv1  gate1421(.a(N2003), .O(gate635inter8));
  nand2 gate1422(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate1423(.a(s_77), .b(gate635inter3), .O(gate635inter10));
  nor2  gate1424(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate1425(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate1426(.a(gate635inter12), .b(gate635inter1), .O(N2040));
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );

  xor2  gate1007(.a(N290), .b(N2061), .O(gate650inter0));
  nand2 gate1008(.a(gate650inter0), .b(s_18), .O(gate650inter1));
  and2  gate1009(.a(N290), .b(N2061), .O(gate650inter2));
  inv1  gate1010(.a(s_18), .O(gate650inter3));
  inv1  gate1011(.a(s_19), .O(gate650inter4));
  nand2 gate1012(.a(gate650inter4), .b(gate650inter3), .O(gate650inter5));
  nor2  gate1013(.a(gate650inter5), .b(gate650inter2), .O(gate650inter6));
  inv1  gate1014(.a(N2061), .O(gate650inter7));
  inv1  gate1015(.a(N290), .O(gate650inter8));
  nand2 gate1016(.a(gate650inter8), .b(gate650inter7), .O(gate650inter9));
  nand2 gate1017(.a(s_19), .b(gate650inter3), .O(gate650inter10));
  nor2  gate1018(.a(gate650inter10), .b(gate650inter9), .O(gate650inter11));
  nor2  gate1019(.a(gate650inter11), .b(gate650inter6), .O(gate650inter12));
  nand2 gate1020(.a(gate650inter12), .b(gate650inter1), .O(N2081));
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate1259(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate1260(.a(gate667inter0), .b(s_54), .O(gate667inter1));
  and2  gate1261(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate1262(.a(s_54), .O(gate667inter3));
  inv1  gate1263(.a(s_55), .O(gate667inter4));
  nand2 gate1264(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate1265(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate1266(.a(N2199), .O(gate667inter7));
  inv1  gate1267(.a(N1348), .O(gate667inter8));
  nand2 gate1268(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate1269(.a(s_55), .b(gate667inter3), .O(gate667inter10));
  nor2  gate1270(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate1271(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate1272(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate895(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate896(.a(gate671inter0), .b(s_2), .O(gate671inter1));
  and2  gate897(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate898(.a(s_2), .O(gate671inter3));
  inv1  gate899(.a(s_3), .O(gate671inter4));
  nand2 gate900(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate901(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate902(.a(N2205), .O(gate671inter7));
  inv1  gate903(.a(N913), .O(gate671inter8));
  nand2 gate904(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate905(.a(s_3), .b(gate671inter3), .O(gate671inter10));
  nor2  gate906(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate907(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate908(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );

  xor2  gate1273(.a(N543), .b(N2570), .O(gate758inter0));
  nand2 gate1274(.a(gate758inter0), .b(s_56), .O(gate758inter1));
  and2  gate1275(.a(N543), .b(N2570), .O(gate758inter2));
  inv1  gate1276(.a(s_56), .O(gate758inter3));
  inv1  gate1277(.a(s_57), .O(gate758inter4));
  nand2 gate1278(.a(gate758inter4), .b(gate758inter3), .O(gate758inter5));
  nor2  gate1279(.a(gate758inter5), .b(gate758inter2), .O(gate758inter6));
  inv1  gate1280(.a(N2570), .O(gate758inter7));
  inv1  gate1281(.a(N543), .O(gate758inter8));
  nand2 gate1282(.a(gate758inter8), .b(gate758inter7), .O(gate758inter9));
  nand2 gate1283(.a(s_57), .b(gate758inter3), .O(gate758inter10));
  nor2  gate1284(.a(gate758inter10), .b(gate758inter9), .O(gate758inter11));
  nor2  gate1285(.a(gate758inter11), .b(gate758inter6), .O(gate758inter12));
  nand2 gate1286(.a(gate758inter12), .b(gate758inter1), .O(N2682));
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );

  xor2  gate1427(.a(N538), .b(N2639), .O(gate769inter0));
  nand2 gate1428(.a(gate769inter0), .b(s_78), .O(gate769inter1));
  and2  gate1429(.a(N538), .b(N2639), .O(gate769inter2));
  inv1  gate1430(.a(s_78), .O(gate769inter3));
  inv1  gate1431(.a(s_79), .O(gate769inter4));
  nand2 gate1432(.a(gate769inter4), .b(gate769inter3), .O(gate769inter5));
  nor2  gate1433(.a(gate769inter5), .b(gate769inter2), .O(gate769inter6));
  inv1  gate1434(.a(N2639), .O(gate769inter7));
  inv1  gate1435(.a(N538), .O(gate769inter8));
  nand2 gate1436(.a(gate769inter8), .b(gate769inter7), .O(gate769inter9));
  nand2 gate1437(.a(s_79), .b(gate769inter3), .O(gate769inter10));
  nor2  gate1438(.a(gate769inter10), .b(gate769inter9), .O(gate769inter11));
  nor2  gate1439(.a(gate769inter11), .b(gate769inter6), .O(gate769inter12));
  nand2 gate1440(.a(gate769inter12), .b(gate769inter1), .O(N2724));
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );

  xor2  gate1301(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1302(.a(gate856inter0), .b(s_60), .O(gate856inter1));
  and2  gate1303(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1304(.a(s_60), .O(gate856inter3));
  inv1  gate1305(.a(s_61), .O(gate856inter4));
  nand2 gate1306(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1307(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1308(.a(N2843), .O(gate856inter7));
  inv1  gate1309(.a(N886), .O(gate856inter8));
  nand2 gate1310(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1311(.a(s_61), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1312(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1313(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1314(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );

  xor2  gate1287(.a(N1461), .b(N2883), .O(gate876inter0));
  nand2 gate1288(.a(gate876inter0), .b(s_58), .O(gate876inter1));
  and2  gate1289(.a(N1461), .b(N2883), .O(gate876inter2));
  inv1  gate1290(.a(s_58), .O(gate876inter3));
  inv1  gate1291(.a(s_59), .O(gate876inter4));
  nand2 gate1292(.a(gate876inter4), .b(gate876inter3), .O(gate876inter5));
  nor2  gate1293(.a(gate876inter5), .b(gate876inter2), .O(gate876inter6));
  inv1  gate1294(.a(N2883), .O(gate876inter7));
  inv1  gate1295(.a(N1461), .O(gate876inter8));
  nand2 gate1296(.a(gate876inter8), .b(gate876inter7), .O(gate876inter9));
  nand2 gate1297(.a(s_59), .b(gate876inter3), .O(gate876inter10));
  nor2  gate1298(.a(gate876inter10), .b(gate876inter9), .O(gate876inter11));
  nor2  gate1299(.a(gate876inter11), .b(gate876inter6), .O(gate876inter12));
  nand2 gate1300(.a(gate876inter12), .b(gate876inter1), .O(N2895));
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );

  xor2  gate1119(.a(N2897), .b(N2895), .O(gate879inter0));
  nand2 gate1120(.a(gate879inter0), .b(s_34), .O(gate879inter1));
  and2  gate1121(.a(N2897), .b(N2895), .O(gate879inter2));
  inv1  gate1122(.a(s_34), .O(gate879inter3));
  inv1  gate1123(.a(s_35), .O(gate879inter4));
  nand2 gate1124(.a(gate879inter4), .b(gate879inter3), .O(gate879inter5));
  nor2  gate1125(.a(gate879inter5), .b(gate879inter2), .O(gate879inter6));
  inv1  gate1126(.a(N2895), .O(gate879inter7));
  inv1  gate1127(.a(N2897), .O(gate879inter8));
  nand2 gate1128(.a(gate879inter8), .b(gate879inter7), .O(gate879inter9));
  nand2 gate1129(.a(s_35), .b(gate879inter3), .O(gate879inter10));
  nor2  gate1130(.a(gate879inter10), .b(gate879inter9), .O(gate879inter11));
  nor2  gate1131(.a(gate879inter11), .b(gate879inter6), .O(gate879inter12));
  nand2 gate1132(.a(gate879inter12), .b(gate879inter1), .O(N2898));
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule