module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate329(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate330(.a(gate3inter0), .b(s_18), .O(gate3inter1));
  and2  gate331(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate332(.a(s_18), .O(gate3inter3));
  inv1  gate333(.a(s_19), .O(gate3inter4));
  nand2 gate334(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate335(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate336(.a(N17), .O(gate3inter7));
  inv1  gate337(.a(N21), .O(gate3inter8));
  nand2 gate338(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate339(.a(s_19), .b(gate3inter3), .O(gate3inter10));
  nor2  gate340(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate341(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate342(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );

  xor2  gate553(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate554(.a(gate5inter0), .b(s_50), .O(gate5inter1));
  and2  gate555(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate556(.a(s_50), .O(gate5inter3));
  inv1  gate557(.a(s_51), .O(gate5inter4));
  nand2 gate558(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate559(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate560(.a(N33), .O(gate5inter7));
  inv1  gate561(.a(N37), .O(gate5inter8));
  nand2 gate562(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate563(.a(s_51), .b(gate5inter3), .O(gate5inter10));
  nor2  gate564(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate565(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate566(.a(gate5inter12), .b(gate5inter1), .O(N254));
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );

  xor2  gate217(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate218(.a(gate13inter0), .b(s_2), .O(gate13inter1));
  and2  gate219(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate220(.a(s_2), .O(gate13inter3));
  inv1  gate221(.a(s_3), .O(gate13inter4));
  nand2 gate222(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate223(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate224(.a(N97), .O(gate13inter7));
  inv1  gate225(.a(N101), .O(gate13inter8));
  nand2 gate226(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate227(.a(s_3), .b(gate13inter3), .O(gate13inter10));
  nor2  gate228(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate229(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate230(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );

  xor2  gate301(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate302(.a(gate16inter0), .b(s_14), .O(gate16inter1));
  and2  gate303(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate304(.a(s_14), .O(gate16inter3));
  inv1  gate305(.a(s_15), .O(gate16inter4));
  nand2 gate306(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate307(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate308(.a(N121), .O(gate16inter7));
  inv1  gate309(.a(N125), .O(gate16inter8));
  nand2 gate310(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate311(.a(s_15), .b(gate16inter3), .O(gate16inter10));
  nor2  gate312(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate313(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate314(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );

  xor2  gate427(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate428(.a(gate26inter0), .b(s_32), .O(gate26inter1));
  and2  gate429(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate430(.a(s_32), .O(gate26inter3));
  inv1  gate431(.a(s_33), .O(gate26inter4));
  nand2 gate432(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate433(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate434(.a(N33), .O(gate26inter7));
  inv1  gate435(.a(N49), .O(gate26inter8));
  nand2 gate436(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate437(.a(s_33), .b(gate26inter3), .O(gate26inter10));
  nor2  gate438(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate439(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate440(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate343(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate344(.a(gate30inter0), .b(s_20), .O(gate30inter1));
  and2  gate345(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate346(.a(s_20), .O(gate30inter3));
  inv1  gate347(.a(s_21), .O(gate30inter4));
  nand2 gate348(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate349(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate350(.a(N41), .O(gate30inter7));
  inv1  gate351(.a(N57), .O(gate30inter8));
  nand2 gate352(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate353(.a(s_21), .b(gate30inter3), .O(gate30inter10));
  nor2  gate354(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate355(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate356(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );

  xor2  gate525(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate526(.a(gate32inter0), .b(s_46), .O(gate32inter1));
  and2  gate527(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate528(.a(s_46), .O(gate32inter3));
  inv1  gate529(.a(s_47), .O(gate32inter4));
  nand2 gate530(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate531(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate532(.a(N45), .O(gate32inter7));
  inv1  gate533(.a(N61), .O(gate32inter8));
  nand2 gate534(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate535(.a(s_47), .b(gate32inter3), .O(gate32inter10));
  nor2  gate536(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate537(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate538(.a(gate32inter12), .b(gate32inter1), .O(N281));
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate441(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate442(.a(gate42inter0), .b(s_34), .O(gate42inter1));
  and2  gate443(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate444(.a(s_34), .O(gate42inter3));
  inv1  gate445(.a(s_35), .O(gate42inter4));
  nand2 gate446(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate447(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate448(.a(N252), .O(gate42inter7));
  inv1  gate449(.a(N253), .O(gate42inter8));
  nand2 gate450(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate451(.a(s_35), .b(gate42inter3), .O(gate42inter10));
  nor2  gate452(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate453(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate454(.a(gate42inter12), .b(gate42inter1), .O(N293));
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate273(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate274(.a(gate47inter0), .b(s_10), .O(gate47inter1));
  and2  gate275(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate276(.a(s_10), .O(gate47inter3));
  inv1  gate277(.a(s_11), .O(gate47inter4));
  nand2 gate278(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate279(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate280(.a(N262), .O(gate47inter7));
  inv1  gate281(.a(N263), .O(gate47inter8));
  nand2 gate282(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate283(.a(s_11), .b(gate47inter3), .O(gate47inter10));
  nor2  gate284(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate285(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate286(.a(gate47inter12), .b(gate47inter1), .O(N308));

  xor2  gate371(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate372(.a(gate48inter0), .b(s_24), .O(gate48inter1));
  and2  gate373(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate374(.a(s_24), .O(gate48inter3));
  inv1  gate375(.a(s_25), .O(gate48inter4));
  nand2 gate376(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate377(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate378(.a(N264), .O(gate48inter7));
  inv1  gate379(.a(N265), .O(gate48inter8));
  nand2 gate380(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate381(.a(s_25), .b(gate48inter3), .O(gate48inter10));
  nor2  gate382(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate383(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate384(.a(gate48inter12), .b(gate48inter1), .O(N311));
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate567(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate568(.a(gate59inter0), .b(s_52), .O(gate59inter1));
  and2  gate569(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate570(.a(s_52), .O(gate59inter3));
  inv1  gate571(.a(s_53), .O(gate59inter4));
  nand2 gate572(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate573(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate574(.a(N290), .O(gate59inter7));
  inv1  gate575(.a(N296), .O(gate59inter8));
  nand2 gate576(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate577(.a(s_53), .b(gate59inter3), .O(gate59inter10));
  nor2  gate578(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate579(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate580(.a(gate59inter12), .b(gate59inter1), .O(N340));

  xor2  gate455(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate456(.a(gate60inter0), .b(s_36), .O(gate60inter1));
  and2  gate457(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate458(.a(s_36), .O(gate60inter3));
  inv1  gate459(.a(s_37), .O(gate60inter4));
  nand2 gate460(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate461(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate462(.a(N293), .O(gate60inter7));
  inv1  gate463(.a(N299), .O(gate60inter8));
  nand2 gate464(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate465(.a(s_37), .b(gate60inter3), .O(gate60inter10));
  nor2  gate466(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate467(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate468(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate581(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate582(.a(gate62inter0), .b(s_54), .O(gate62inter1));
  and2  gate583(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate584(.a(s_54), .O(gate62inter3));
  inv1  gate585(.a(s_55), .O(gate62inter4));
  nand2 gate586(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate587(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate588(.a(N308), .O(gate62inter7));
  inv1  gate589(.a(N311), .O(gate62inter8));
  nand2 gate590(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate591(.a(s_55), .b(gate62inter3), .O(gate62inter10));
  nor2  gate592(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate593(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate594(.a(gate62inter12), .b(gate62inter1), .O(N343));

  xor2  gate469(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate470(.a(gate63inter0), .b(s_38), .O(gate63inter1));
  and2  gate471(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate472(.a(s_38), .O(gate63inter3));
  inv1  gate473(.a(s_39), .O(gate63inter4));
  nand2 gate474(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate475(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate476(.a(N302), .O(gate63inter7));
  inv1  gate477(.a(N308), .O(gate63inter8));
  nand2 gate478(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate479(.a(s_39), .b(gate63inter3), .O(gate63inter10));
  nor2  gate480(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate481(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate482(.a(gate63inter12), .b(gate63inter1), .O(N344));
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate609(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate610(.a(gate65inter0), .b(s_58), .O(gate65inter1));
  and2  gate611(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate612(.a(s_58), .O(gate65inter3));
  inv1  gate613(.a(s_59), .O(gate65inter4));
  nand2 gate614(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate615(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate616(.a(N266), .O(gate65inter7));
  inv1  gate617(.a(N342), .O(gate65inter8));
  nand2 gate618(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate619(.a(s_59), .b(gate65inter3), .O(gate65inter10));
  nor2  gate620(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate621(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate622(.a(gate65inter12), .b(gate65inter1), .O(N346));
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate385(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate386(.a(gate70inter0), .b(s_26), .O(gate70inter1));
  and2  gate387(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate388(.a(s_26), .O(gate70inter3));
  inv1  gate389(.a(s_27), .O(gate70inter4));
  nand2 gate390(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate391(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate392(.a(N271), .O(gate70inter7));
  inv1  gate393(.a(N339), .O(gate70inter8));
  nand2 gate394(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate395(.a(s_27), .b(gate70inter3), .O(gate70inter10));
  nor2  gate396(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate397(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate398(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );

  xor2  gate259(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate260(.a(gate76inter0), .b(s_8), .O(gate76inter1));
  and2  gate261(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate262(.a(s_8), .O(gate76inter3));
  inv1  gate263(.a(s_9), .O(gate76inter4));
  nand2 gate264(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate265(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate266(.a(N317), .O(gate76inter7));
  inv1  gate267(.a(N349), .O(gate76inter8));
  nand2 gate268(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate269(.a(s_9), .b(gate76inter3), .O(gate76inter10));
  nor2  gate270(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate271(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate272(.a(gate76inter12), .b(gate76inter1), .O(N393));
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate511(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate512(.a(gate172inter0), .b(s_44), .O(gate172inter1));
  and2  gate513(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate514(.a(s_44), .O(gate172inter3));
  inv1  gate515(.a(s_45), .O(gate172inter4));
  nand2 gate516(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate517(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate518(.a(N5), .O(gate172inter7));
  inv1  gate519(.a(N693), .O(gate172inter8));
  nand2 gate520(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate521(.a(s_45), .b(gate172inter3), .O(gate172inter10));
  nor2  gate522(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate523(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate524(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );

  xor2  gate287(.a(N696), .b(N17), .O(gate175inter0));
  nand2 gate288(.a(gate175inter0), .b(s_12), .O(gate175inter1));
  and2  gate289(.a(N696), .b(N17), .O(gate175inter2));
  inv1  gate290(.a(s_12), .O(gate175inter3));
  inv1  gate291(.a(s_13), .O(gate175inter4));
  nand2 gate292(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate293(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate294(.a(N17), .O(gate175inter7));
  inv1  gate295(.a(N696), .O(gate175inter8));
  nand2 gate296(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate297(.a(s_13), .b(gate175inter3), .O(gate175inter10));
  nor2  gate298(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate299(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate300(.a(gate175inter12), .b(gate175inter1), .O(N728));
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );

  xor2  gate539(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate540(.a(gate179inter0), .b(s_48), .O(gate179inter1));
  and2  gate541(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate542(.a(s_48), .O(gate179inter3));
  inv1  gate543(.a(s_49), .O(gate179inter4));
  nand2 gate544(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate545(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate546(.a(N33), .O(gate179inter7));
  inv1  gate547(.a(N700), .O(gate179inter8));
  nand2 gate548(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate549(.a(s_49), .b(gate179inter3), .O(gate179inter10));
  nor2  gate550(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate551(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate552(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );

  xor2  gate595(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate596(.a(gate181inter0), .b(s_56), .O(gate181inter1));
  and2  gate597(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate598(.a(s_56), .O(gate181inter3));
  inv1  gate599(.a(s_57), .O(gate181inter4));
  nand2 gate600(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate601(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate602(.a(N41), .O(gate181inter7));
  inv1  gate603(.a(N702), .O(gate181inter8));
  nand2 gate604(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate605(.a(s_57), .b(gate181inter3), .O(gate181inter10));
  nor2  gate606(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate607(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate608(.a(gate181inter12), .b(gate181inter1), .O(N734));
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );

  xor2  gate245(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate246(.a(gate184inter0), .b(s_6), .O(gate184inter1));
  and2  gate247(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate248(.a(s_6), .O(gate184inter3));
  inv1  gate249(.a(s_7), .O(gate184inter4));
  nand2 gate250(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate251(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate252(.a(N53), .O(gate184inter7));
  inv1  gate253(.a(N705), .O(gate184inter8));
  nand2 gate254(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate255(.a(s_7), .b(gate184inter3), .O(gate184inter10));
  nor2  gate256(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate257(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate258(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate357(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate358(.a(gate186inter0), .b(s_22), .O(gate186inter1));
  and2  gate359(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate360(.a(s_22), .O(gate186inter3));
  inv1  gate361(.a(s_23), .O(gate186inter4));
  nand2 gate362(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate363(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate364(.a(N61), .O(gate186inter7));
  inv1  gate365(.a(N707), .O(gate186inter8));
  nand2 gate366(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate367(.a(s_23), .b(gate186inter3), .O(gate186inter10));
  nor2  gate368(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate369(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate370(.a(gate186inter12), .b(gate186inter1), .O(N739));

  xor2  gate203(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate204(.a(gate187inter0), .b(s_0), .O(gate187inter1));
  and2  gate205(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate206(.a(s_0), .O(gate187inter3));
  inv1  gate207(.a(s_1), .O(gate187inter4));
  nand2 gate208(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate209(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate210(.a(N65), .O(gate187inter7));
  inv1  gate211(.a(N708), .O(gate187inter8));
  nand2 gate212(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate213(.a(s_1), .b(gate187inter3), .O(gate187inter10));
  nor2  gate214(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate215(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate216(.a(gate187inter12), .b(gate187inter1), .O(N740));
xor2 gate188( .a(N69), .b(N709), .O(N741) );

  xor2  gate413(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate414(.a(gate189inter0), .b(s_30), .O(gate189inter1));
  and2  gate415(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate416(.a(s_30), .O(gate189inter3));
  inv1  gate417(.a(s_31), .O(gate189inter4));
  nand2 gate418(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate419(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate420(.a(N73), .O(gate189inter7));
  inv1  gate421(.a(N710), .O(gate189inter8));
  nand2 gate422(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate423(.a(s_31), .b(gate189inter3), .O(gate189inter10));
  nor2  gate424(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate425(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate426(.a(gate189inter12), .b(gate189inter1), .O(N742));
xor2 gate190( .a(N77), .b(N711), .O(N743) );

  xor2  gate623(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate624(.a(gate191inter0), .b(s_60), .O(gate191inter1));
  and2  gate625(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate626(.a(s_60), .O(gate191inter3));
  inv1  gate627(.a(s_61), .O(gate191inter4));
  nand2 gate628(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate629(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate630(.a(N81), .O(gate191inter7));
  inv1  gate631(.a(N712), .O(gate191inter8));
  nand2 gate632(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate633(.a(s_61), .b(gate191inter3), .O(gate191inter10));
  nor2  gate634(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate635(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate636(.a(gate191inter12), .b(gate191inter1), .O(N744));

  xor2  gate497(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate498(.a(gate192inter0), .b(s_42), .O(gate192inter1));
  and2  gate499(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate500(.a(s_42), .O(gate192inter3));
  inv1  gate501(.a(s_43), .O(gate192inter4));
  nand2 gate502(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate503(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate504(.a(N85), .O(gate192inter7));
  inv1  gate505(.a(N713), .O(gate192inter8));
  nand2 gate506(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate507(.a(s_43), .b(gate192inter3), .O(gate192inter10));
  nor2  gate508(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate509(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate510(.a(gate192inter12), .b(gate192inter1), .O(N745));

  xor2  gate231(.a(N714), .b(N89), .O(gate193inter0));
  nand2 gate232(.a(gate193inter0), .b(s_4), .O(gate193inter1));
  and2  gate233(.a(N714), .b(N89), .O(gate193inter2));
  inv1  gate234(.a(s_4), .O(gate193inter3));
  inv1  gate235(.a(s_5), .O(gate193inter4));
  nand2 gate236(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate237(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate238(.a(N89), .O(gate193inter7));
  inv1  gate239(.a(N714), .O(gate193inter8));
  nand2 gate240(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate241(.a(s_5), .b(gate193inter3), .O(gate193inter10));
  nor2  gate242(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate243(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate244(.a(gate193inter12), .b(gate193inter1), .O(N746));
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );

  xor2  gate315(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate316(.a(gate196inter0), .b(s_16), .O(gate196inter1));
  and2  gate317(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate318(.a(s_16), .O(gate196inter3));
  inv1  gate319(.a(s_17), .O(gate196inter4));
  nand2 gate320(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate321(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate322(.a(N101), .O(gate196inter7));
  inv1  gate323(.a(N717), .O(gate196inter8));
  nand2 gate324(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate325(.a(s_17), .b(gate196inter3), .O(gate196inter10));
  nor2  gate326(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate327(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate328(.a(gate196inter12), .b(gate196inter1), .O(N749));
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );

  xor2  gate483(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate484(.a(gate199inter0), .b(s_40), .O(gate199inter1));
  and2  gate485(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate486(.a(s_40), .O(gate199inter3));
  inv1  gate487(.a(s_41), .O(gate199inter4));
  nand2 gate488(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate489(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate490(.a(N113), .O(gate199inter7));
  inv1  gate491(.a(N720), .O(gate199inter8));
  nand2 gate492(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate493(.a(s_41), .b(gate199inter3), .O(gate199inter10));
  nor2  gate494(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate495(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate496(.a(gate199inter12), .b(gate199inter1), .O(N752));
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );

  xor2  gate399(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate400(.a(gate202inter0), .b(s_28), .O(gate202inter1));
  and2  gate401(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate402(.a(s_28), .O(gate202inter3));
  inv1  gate403(.a(s_29), .O(gate202inter4));
  nand2 gate404(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate405(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate406(.a(N125), .O(gate202inter7));
  inv1  gate407(.a(N723), .O(gate202inter8));
  nand2 gate408(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate409(.a(s_29), .b(gate202inter3), .O(gate202inter10));
  nor2  gate410(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate411(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate412(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule