module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2787(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2788(.a(gate14inter0), .b(s_320), .O(gate14inter1));
  and2  gate2789(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2790(.a(s_320), .O(gate14inter3));
  inv1  gate2791(.a(s_321), .O(gate14inter4));
  nand2 gate2792(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2793(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2794(.a(G11), .O(gate14inter7));
  inv1  gate2795(.a(G12), .O(gate14inter8));
  nand2 gate2796(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2797(.a(s_321), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2798(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2799(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2800(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1107(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1108(.a(gate15inter0), .b(s_80), .O(gate15inter1));
  and2  gate1109(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1110(.a(s_80), .O(gate15inter3));
  inv1  gate1111(.a(s_81), .O(gate15inter4));
  nand2 gate1112(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1113(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1114(.a(G13), .O(gate15inter7));
  inv1  gate1115(.a(G14), .O(gate15inter8));
  nand2 gate1116(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1117(.a(s_81), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1118(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1119(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1120(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate659(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate660(.a(gate16inter0), .b(s_16), .O(gate16inter1));
  and2  gate661(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate662(.a(s_16), .O(gate16inter3));
  inv1  gate663(.a(s_17), .O(gate16inter4));
  nand2 gate664(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate665(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate666(.a(G15), .O(gate16inter7));
  inv1  gate667(.a(G16), .O(gate16inter8));
  nand2 gate668(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate669(.a(s_17), .b(gate16inter3), .O(gate16inter10));
  nor2  gate670(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate671(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate672(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2899(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2900(.a(gate17inter0), .b(s_336), .O(gate17inter1));
  and2  gate2901(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2902(.a(s_336), .O(gate17inter3));
  inv1  gate2903(.a(s_337), .O(gate17inter4));
  nand2 gate2904(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2905(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2906(.a(G17), .O(gate17inter7));
  inv1  gate2907(.a(G18), .O(gate17inter8));
  nand2 gate2908(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2909(.a(s_337), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2910(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2911(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2912(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2185(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2186(.a(gate27inter0), .b(s_234), .O(gate27inter1));
  and2  gate2187(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2188(.a(s_234), .O(gate27inter3));
  inv1  gate2189(.a(s_235), .O(gate27inter4));
  nand2 gate2190(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2191(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2192(.a(G2), .O(gate27inter7));
  inv1  gate2193(.a(G6), .O(gate27inter8));
  nand2 gate2194(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2195(.a(s_235), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2196(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2197(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2198(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1653(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1654(.a(gate28inter0), .b(s_158), .O(gate28inter1));
  and2  gate1655(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1656(.a(s_158), .O(gate28inter3));
  inv1  gate1657(.a(s_159), .O(gate28inter4));
  nand2 gate1658(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1659(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1660(.a(G10), .O(gate28inter7));
  inv1  gate1661(.a(G14), .O(gate28inter8));
  nand2 gate1662(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1663(.a(s_159), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1664(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1665(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1666(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate799(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate800(.a(gate29inter0), .b(s_36), .O(gate29inter1));
  and2  gate801(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate802(.a(s_36), .O(gate29inter3));
  inv1  gate803(.a(s_37), .O(gate29inter4));
  nand2 gate804(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate805(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate806(.a(G3), .O(gate29inter7));
  inv1  gate807(.a(G7), .O(gate29inter8));
  nand2 gate808(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate809(.a(s_37), .b(gate29inter3), .O(gate29inter10));
  nor2  gate810(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate811(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate812(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1933(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1934(.a(gate30inter0), .b(s_198), .O(gate30inter1));
  and2  gate1935(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1936(.a(s_198), .O(gate30inter3));
  inv1  gate1937(.a(s_199), .O(gate30inter4));
  nand2 gate1938(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1939(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1940(.a(G11), .O(gate30inter7));
  inv1  gate1941(.a(G15), .O(gate30inter8));
  nand2 gate1942(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1943(.a(s_199), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1944(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1945(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1946(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1135(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1136(.a(gate33inter0), .b(s_84), .O(gate33inter1));
  and2  gate1137(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1138(.a(s_84), .O(gate33inter3));
  inv1  gate1139(.a(s_85), .O(gate33inter4));
  nand2 gate1140(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1141(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1142(.a(G17), .O(gate33inter7));
  inv1  gate1143(.a(G21), .O(gate33inter8));
  nand2 gate1144(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1145(.a(s_85), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1146(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1147(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1148(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate995(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate996(.a(gate34inter0), .b(s_64), .O(gate34inter1));
  and2  gate997(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate998(.a(s_64), .O(gate34inter3));
  inv1  gate999(.a(s_65), .O(gate34inter4));
  nand2 gate1000(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1001(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1002(.a(G25), .O(gate34inter7));
  inv1  gate1003(.a(G29), .O(gate34inter8));
  nand2 gate1004(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1005(.a(s_65), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1006(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1007(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1008(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2549(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2550(.a(gate36inter0), .b(s_286), .O(gate36inter1));
  and2  gate2551(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2552(.a(s_286), .O(gate36inter3));
  inv1  gate2553(.a(s_287), .O(gate36inter4));
  nand2 gate2554(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2555(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2556(.a(G26), .O(gate36inter7));
  inv1  gate2557(.a(G30), .O(gate36inter8));
  nand2 gate2558(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2559(.a(s_287), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2560(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2561(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2562(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate2087(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2088(.a(gate37inter0), .b(s_220), .O(gate37inter1));
  and2  gate2089(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2090(.a(s_220), .O(gate37inter3));
  inv1  gate2091(.a(s_221), .O(gate37inter4));
  nand2 gate2092(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2093(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2094(.a(G19), .O(gate37inter7));
  inv1  gate2095(.a(G23), .O(gate37inter8));
  nand2 gate2096(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2097(.a(s_221), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2098(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2099(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2100(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2465(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2466(.a(gate39inter0), .b(s_274), .O(gate39inter1));
  and2  gate2467(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2468(.a(s_274), .O(gate39inter3));
  inv1  gate2469(.a(s_275), .O(gate39inter4));
  nand2 gate2470(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2471(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2472(.a(G20), .O(gate39inter7));
  inv1  gate2473(.a(G24), .O(gate39inter8));
  nand2 gate2474(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2475(.a(s_275), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2476(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2477(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2478(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1415(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1416(.a(gate41inter0), .b(s_124), .O(gate41inter1));
  and2  gate1417(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1418(.a(s_124), .O(gate41inter3));
  inv1  gate1419(.a(s_125), .O(gate41inter4));
  nand2 gate1420(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1421(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1422(.a(G1), .O(gate41inter7));
  inv1  gate1423(.a(G266), .O(gate41inter8));
  nand2 gate1424(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1425(.a(s_125), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1426(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1427(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1428(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2619(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2620(.a(gate42inter0), .b(s_296), .O(gate42inter1));
  and2  gate2621(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2622(.a(s_296), .O(gate42inter3));
  inv1  gate2623(.a(s_297), .O(gate42inter4));
  nand2 gate2624(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2625(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2626(.a(G2), .O(gate42inter7));
  inv1  gate2627(.a(G266), .O(gate42inter8));
  nand2 gate2628(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2629(.a(s_297), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2630(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2631(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2632(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate2003(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2004(.a(gate45inter0), .b(s_208), .O(gate45inter1));
  and2  gate2005(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2006(.a(s_208), .O(gate45inter3));
  inv1  gate2007(.a(s_209), .O(gate45inter4));
  nand2 gate2008(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2009(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2010(.a(G5), .O(gate45inter7));
  inv1  gate2011(.a(G272), .O(gate45inter8));
  nand2 gate2012(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2013(.a(s_209), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2014(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2015(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2016(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1065(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1066(.a(gate46inter0), .b(s_74), .O(gate46inter1));
  and2  gate1067(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1068(.a(s_74), .O(gate46inter3));
  inv1  gate1069(.a(s_75), .O(gate46inter4));
  nand2 gate1070(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1071(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1072(.a(G6), .O(gate46inter7));
  inv1  gate1073(.a(G272), .O(gate46inter8));
  nand2 gate1074(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1075(.a(s_75), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1076(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1077(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1078(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1401(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1402(.a(gate47inter0), .b(s_122), .O(gate47inter1));
  and2  gate1403(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1404(.a(s_122), .O(gate47inter3));
  inv1  gate1405(.a(s_123), .O(gate47inter4));
  nand2 gate1406(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1407(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1408(.a(G7), .O(gate47inter7));
  inv1  gate1409(.a(G275), .O(gate47inter8));
  nand2 gate1410(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1411(.a(s_123), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1412(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1413(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1414(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1233(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1234(.a(gate48inter0), .b(s_98), .O(gate48inter1));
  and2  gate1235(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1236(.a(s_98), .O(gate48inter3));
  inv1  gate1237(.a(s_99), .O(gate48inter4));
  nand2 gate1238(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1239(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1240(.a(G8), .O(gate48inter7));
  inv1  gate1241(.a(G275), .O(gate48inter8));
  nand2 gate1242(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1243(.a(s_99), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1244(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1245(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1246(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2297(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2298(.a(gate54inter0), .b(s_250), .O(gate54inter1));
  and2  gate2299(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2300(.a(s_250), .O(gate54inter3));
  inv1  gate2301(.a(s_251), .O(gate54inter4));
  nand2 gate2302(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2303(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2304(.a(G14), .O(gate54inter7));
  inv1  gate2305(.a(G284), .O(gate54inter8));
  nand2 gate2306(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2307(.a(s_251), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2308(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2309(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2310(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1331(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1332(.a(gate55inter0), .b(s_112), .O(gate55inter1));
  and2  gate1333(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1334(.a(s_112), .O(gate55inter3));
  inv1  gate1335(.a(s_113), .O(gate55inter4));
  nand2 gate1336(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1337(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1338(.a(G15), .O(gate55inter7));
  inv1  gate1339(.a(G287), .O(gate55inter8));
  nand2 gate1340(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1341(.a(s_113), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1342(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1343(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1344(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1303(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1304(.a(gate56inter0), .b(s_108), .O(gate56inter1));
  and2  gate1305(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1306(.a(s_108), .O(gate56inter3));
  inv1  gate1307(.a(s_109), .O(gate56inter4));
  nand2 gate1308(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1309(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1310(.a(G16), .O(gate56inter7));
  inv1  gate1311(.a(G287), .O(gate56inter8));
  nand2 gate1312(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1313(.a(s_109), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1314(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1315(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1316(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate631(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate632(.a(gate59inter0), .b(s_12), .O(gate59inter1));
  and2  gate633(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate634(.a(s_12), .O(gate59inter3));
  inv1  gate635(.a(s_13), .O(gate59inter4));
  nand2 gate636(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate637(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate638(.a(G19), .O(gate59inter7));
  inv1  gate639(.a(G293), .O(gate59inter8));
  nand2 gate640(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate641(.a(s_13), .b(gate59inter3), .O(gate59inter10));
  nor2  gate642(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate643(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate644(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1737(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1738(.a(gate60inter0), .b(s_170), .O(gate60inter1));
  and2  gate1739(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1740(.a(s_170), .O(gate60inter3));
  inv1  gate1741(.a(s_171), .O(gate60inter4));
  nand2 gate1742(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1743(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1744(.a(G20), .O(gate60inter7));
  inv1  gate1745(.a(G293), .O(gate60inter8));
  nand2 gate1746(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1747(.a(s_171), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1748(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1749(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1750(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1499(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1500(.a(gate64inter0), .b(s_136), .O(gate64inter1));
  and2  gate1501(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1502(.a(s_136), .O(gate64inter3));
  inv1  gate1503(.a(s_137), .O(gate64inter4));
  nand2 gate1504(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1505(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1506(.a(G24), .O(gate64inter7));
  inv1  gate1507(.a(G299), .O(gate64inter8));
  nand2 gate1508(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1509(.a(s_137), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1510(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1511(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1512(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate729(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate730(.a(gate68inter0), .b(s_26), .O(gate68inter1));
  and2  gate731(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate732(.a(s_26), .O(gate68inter3));
  inv1  gate733(.a(s_27), .O(gate68inter4));
  nand2 gate734(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate735(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate736(.a(G28), .O(gate68inter7));
  inv1  gate737(.a(G305), .O(gate68inter8));
  nand2 gate738(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate739(.a(s_27), .b(gate68inter3), .O(gate68inter10));
  nor2  gate740(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate741(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate742(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate715(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate716(.a(gate69inter0), .b(s_24), .O(gate69inter1));
  and2  gate717(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate718(.a(s_24), .O(gate69inter3));
  inv1  gate719(.a(s_25), .O(gate69inter4));
  nand2 gate720(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate721(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate722(.a(G29), .O(gate69inter7));
  inv1  gate723(.a(G308), .O(gate69inter8));
  nand2 gate724(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate725(.a(s_25), .b(gate69inter3), .O(gate69inter10));
  nor2  gate726(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate727(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate728(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2703(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2704(.a(gate70inter0), .b(s_308), .O(gate70inter1));
  and2  gate2705(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2706(.a(s_308), .O(gate70inter3));
  inv1  gate2707(.a(s_309), .O(gate70inter4));
  nand2 gate2708(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2709(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2710(.a(G30), .O(gate70inter7));
  inv1  gate2711(.a(G308), .O(gate70inter8));
  nand2 gate2712(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2713(.a(s_309), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2714(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2715(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2716(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate2339(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2340(.a(gate71inter0), .b(s_256), .O(gate71inter1));
  and2  gate2341(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2342(.a(s_256), .O(gate71inter3));
  inv1  gate2343(.a(s_257), .O(gate71inter4));
  nand2 gate2344(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2345(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2346(.a(G31), .O(gate71inter7));
  inv1  gate2347(.a(G311), .O(gate71inter8));
  nand2 gate2348(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2349(.a(s_257), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2350(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2351(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2352(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2101(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2102(.a(gate72inter0), .b(s_222), .O(gate72inter1));
  and2  gate2103(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2104(.a(s_222), .O(gate72inter3));
  inv1  gate2105(.a(s_223), .O(gate72inter4));
  nand2 gate2106(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2107(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2108(.a(G32), .O(gate72inter7));
  inv1  gate2109(.a(G311), .O(gate72inter8));
  nand2 gate2110(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2111(.a(s_223), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2112(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2113(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2114(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate2773(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2774(.a(gate73inter0), .b(s_318), .O(gate73inter1));
  and2  gate2775(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2776(.a(s_318), .O(gate73inter3));
  inv1  gate2777(.a(s_319), .O(gate73inter4));
  nand2 gate2778(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2779(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2780(.a(G1), .O(gate73inter7));
  inv1  gate2781(.a(G314), .O(gate73inter8));
  nand2 gate2782(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2783(.a(s_319), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2784(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2785(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2786(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate771(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate772(.a(gate75inter0), .b(s_32), .O(gate75inter1));
  and2  gate773(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate774(.a(s_32), .O(gate75inter3));
  inv1  gate775(.a(s_33), .O(gate75inter4));
  nand2 gate776(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate777(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate778(.a(G9), .O(gate75inter7));
  inv1  gate779(.a(G317), .O(gate75inter8));
  nand2 gate780(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate781(.a(s_33), .b(gate75inter3), .O(gate75inter10));
  nor2  gate782(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate783(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate784(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2157(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2158(.a(gate79inter0), .b(s_230), .O(gate79inter1));
  and2  gate2159(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2160(.a(s_230), .O(gate79inter3));
  inv1  gate2161(.a(s_231), .O(gate79inter4));
  nand2 gate2162(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2163(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2164(.a(G10), .O(gate79inter7));
  inv1  gate2165(.a(G323), .O(gate79inter8));
  nand2 gate2166(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2167(.a(s_231), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2168(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2169(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2170(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2633(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2634(.a(gate84inter0), .b(s_298), .O(gate84inter1));
  and2  gate2635(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2636(.a(s_298), .O(gate84inter3));
  inv1  gate2637(.a(s_299), .O(gate84inter4));
  nand2 gate2638(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2639(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2640(.a(G15), .O(gate84inter7));
  inv1  gate2641(.a(G329), .O(gate84inter8));
  nand2 gate2642(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2643(.a(s_299), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2644(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2645(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2646(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate981(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate982(.a(gate85inter0), .b(s_62), .O(gate85inter1));
  and2  gate983(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate984(.a(s_62), .O(gate85inter3));
  inv1  gate985(.a(s_63), .O(gate85inter4));
  nand2 gate986(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate987(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate988(.a(G4), .O(gate85inter7));
  inv1  gate989(.a(G332), .O(gate85inter8));
  nand2 gate990(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate991(.a(s_63), .b(gate85inter3), .O(gate85inter10));
  nor2  gate992(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate993(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate994(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1667(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1668(.a(gate86inter0), .b(s_160), .O(gate86inter1));
  and2  gate1669(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1670(.a(s_160), .O(gate86inter3));
  inv1  gate1671(.a(s_161), .O(gate86inter4));
  nand2 gate1672(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1673(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1674(.a(G8), .O(gate86inter7));
  inv1  gate1675(.a(G332), .O(gate86inter8));
  nand2 gate1676(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1677(.a(s_161), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1678(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1679(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1680(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1821(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1822(.a(gate90inter0), .b(s_182), .O(gate90inter1));
  and2  gate1823(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1824(.a(s_182), .O(gate90inter3));
  inv1  gate1825(.a(s_183), .O(gate90inter4));
  nand2 gate1826(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1827(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1828(.a(G21), .O(gate90inter7));
  inv1  gate1829(.a(G338), .O(gate90inter8));
  nand2 gate1830(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1831(.a(s_183), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1832(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1833(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1834(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1625(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1626(.a(gate93inter0), .b(s_154), .O(gate93inter1));
  and2  gate1627(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1628(.a(s_154), .O(gate93inter3));
  inv1  gate1629(.a(s_155), .O(gate93inter4));
  nand2 gate1630(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1631(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1632(.a(G18), .O(gate93inter7));
  inv1  gate1633(.a(G344), .O(gate93inter8));
  nand2 gate1634(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1635(.a(s_155), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1636(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1637(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1638(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1891(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1892(.a(gate94inter0), .b(s_192), .O(gate94inter1));
  and2  gate1893(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1894(.a(s_192), .O(gate94inter3));
  inv1  gate1895(.a(s_193), .O(gate94inter4));
  nand2 gate1896(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1897(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1898(.a(G22), .O(gate94inter7));
  inv1  gate1899(.a(G344), .O(gate94inter8));
  nand2 gate1900(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1901(.a(s_193), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1902(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1903(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1904(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate2801(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2802(.a(gate95inter0), .b(s_322), .O(gate95inter1));
  and2  gate2803(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2804(.a(s_322), .O(gate95inter3));
  inv1  gate2805(.a(s_323), .O(gate95inter4));
  nand2 gate2806(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2807(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2808(.a(G26), .O(gate95inter7));
  inv1  gate2809(.a(G347), .O(gate95inter8));
  nand2 gate2810(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2811(.a(s_323), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2812(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2813(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2814(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2381(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2382(.a(gate98inter0), .b(s_262), .O(gate98inter1));
  and2  gate2383(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2384(.a(s_262), .O(gate98inter3));
  inv1  gate2385(.a(s_263), .O(gate98inter4));
  nand2 gate2386(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2387(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2388(.a(G23), .O(gate98inter7));
  inv1  gate2389(.a(G350), .O(gate98inter8));
  nand2 gate2390(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2391(.a(s_263), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2392(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2393(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2394(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2059(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2060(.a(gate100inter0), .b(s_216), .O(gate100inter1));
  and2  gate2061(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2062(.a(s_216), .O(gate100inter3));
  inv1  gate2063(.a(s_217), .O(gate100inter4));
  nand2 gate2064(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2065(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2066(.a(G31), .O(gate100inter7));
  inv1  gate2067(.a(G353), .O(gate100inter8));
  nand2 gate2068(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2069(.a(s_217), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2070(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2071(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2072(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate603(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate604(.a(gate101inter0), .b(s_8), .O(gate101inter1));
  and2  gate605(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate606(.a(s_8), .O(gate101inter3));
  inv1  gate607(.a(s_9), .O(gate101inter4));
  nand2 gate608(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate609(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate610(.a(G20), .O(gate101inter7));
  inv1  gate611(.a(G356), .O(gate101inter8));
  nand2 gate612(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate613(.a(s_9), .b(gate101inter3), .O(gate101inter10));
  nor2  gate614(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate615(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate616(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2591(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2592(.a(gate102inter0), .b(s_292), .O(gate102inter1));
  and2  gate2593(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2594(.a(s_292), .O(gate102inter3));
  inv1  gate2595(.a(s_293), .O(gate102inter4));
  nand2 gate2596(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2597(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2598(.a(G24), .O(gate102inter7));
  inv1  gate2599(.a(G356), .O(gate102inter8));
  nand2 gate2600(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2601(.a(s_293), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2602(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2603(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2604(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate785(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate786(.a(gate106inter0), .b(s_34), .O(gate106inter1));
  and2  gate787(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate788(.a(s_34), .O(gate106inter3));
  inv1  gate789(.a(s_35), .O(gate106inter4));
  nand2 gate790(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate791(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate792(.a(G364), .O(gate106inter7));
  inv1  gate793(.a(G365), .O(gate106inter8));
  nand2 gate794(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate795(.a(s_35), .b(gate106inter3), .O(gate106inter10));
  nor2  gate796(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate797(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate798(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2507(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2508(.a(gate108inter0), .b(s_280), .O(gate108inter1));
  and2  gate2509(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2510(.a(s_280), .O(gate108inter3));
  inv1  gate2511(.a(s_281), .O(gate108inter4));
  nand2 gate2512(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2513(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2514(.a(G368), .O(gate108inter7));
  inv1  gate2515(.a(G369), .O(gate108inter8));
  nand2 gate2516(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2517(.a(s_281), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2518(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2519(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2520(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2815(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2816(.a(gate110inter0), .b(s_324), .O(gate110inter1));
  and2  gate2817(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2818(.a(s_324), .O(gate110inter3));
  inv1  gate2819(.a(s_325), .O(gate110inter4));
  nand2 gate2820(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2821(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2822(.a(G372), .O(gate110inter7));
  inv1  gate2823(.a(G373), .O(gate110inter8));
  nand2 gate2824(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2825(.a(s_325), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2826(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2827(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2828(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2717(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2718(.a(gate111inter0), .b(s_310), .O(gate111inter1));
  and2  gate2719(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2720(.a(s_310), .O(gate111inter3));
  inv1  gate2721(.a(s_311), .O(gate111inter4));
  nand2 gate2722(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2723(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2724(.a(G374), .O(gate111inter7));
  inv1  gate2725(.a(G375), .O(gate111inter8));
  nand2 gate2726(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2727(.a(s_311), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2728(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2729(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2730(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1723(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1724(.a(gate113inter0), .b(s_168), .O(gate113inter1));
  and2  gate1725(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1726(.a(s_168), .O(gate113inter3));
  inv1  gate1727(.a(s_169), .O(gate113inter4));
  nand2 gate1728(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1729(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1730(.a(G378), .O(gate113inter7));
  inv1  gate1731(.a(G379), .O(gate113inter8));
  nand2 gate1732(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1733(.a(s_169), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1734(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1735(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1736(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1121(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1122(.a(gate119inter0), .b(s_82), .O(gate119inter1));
  and2  gate1123(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1124(.a(s_82), .O(gate119inter3));
  inv1  gate1125(.a(s_83), .O(gate119inter4));
  nand2 gate1126(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1127(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1128(.a(G390), .O(gate119inter7));
  inv1  gate1129(.a(G391), .O(gate119inter8));
  nand2 gate1130(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1131(.a(s_83), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1132(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1133(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1134(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1793(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1794(.a(gate121inter0), .b(s_178), .O(gate121inter1));
  and2  gate1795(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1796(.a(s_178), .O(gate121inter3));
  inv1  gate1797(.a(s_179), .O(gate121inter4));
  nand2 gate1798(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1799(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1800(.a(G394), .O(gate121inter7));
  inv1  gate1801(.a(G395), .O(gate121inter8));
  nand2 gate1802(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1803(.a(s_179), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1804(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1805(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1806(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate869(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate870(.a(gate122inter0), .b(s_46), .O(gate122inter1));
  and2  gate871(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate872(.a(s_46), .O(gate122inter3));
  inv1  gate873(.a(s_47), .O(gate122inter4));
  nand2 gate874(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate875(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate876(.a(G396), .O(gate122inter7));
  inv1  gate877(.a(G397), .O(gate122inter8));
  nand2 gate878(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate879(.a(s_47), .b(gate122inter3), .O(gate122inter10));
  nor2  gate880(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate881(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate882(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2675(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2676(.a(gate125inter0), .b(s_304), .O(gate125inter1));
  and2  gate2677(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2678(.a(s_304), .O(gate125inter3));
  inv1  gate2679(.a(s_305), .O(gate125inter4));
  nand2 gate2680(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2681(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2682(.a(G402), .O(gate125inter7));
  inv1  gate2683(.a(G403), .O(gate125inter8));
  nand2 gate2684(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2685(.a(s_305), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2686(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2687(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2688(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1527(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1528(.a(gate128inter0), .b(s_140), .O(gate128inter1));
  and2  gate1529(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1530(.a(s_140), .O(gate128inter3));
  inv1  gate1531(.a(s_141), .O(gate128inter4));
  nand2 gate1532(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1533(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1534(.a(G408), .O(gate128inter7));
  inv1  gate1535(.a(G409), .O(gate128inter8));
  nand2 gate1536(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1537(.a(s_141), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1538(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1539(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1540(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1569(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1570(.a(gate131inter0), .b(s_146), .O(gate131inter1));
  and2  gate1571(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1572(.a(s_146), .O(gate131inter3));
  inv1  gate1573(.a(s_147), .O(gate131inter4));
  nand2 gate1574(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1575(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1576(.a(G414), .O(gate131inter7));
  inv1  gate1577(.a(G415), .O(gate131inter8));
  nand2 gate1578(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1579(.a(s_147), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1580(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1581(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1582(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate855(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate856(.a(gate132inter0), .b(s_44), .O(gate132inter1));
  and2  gate857(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate858(.a(s_44), .O(gate132inter3));
  inv1  gate859(.a(s_45), .O(gate132inter4));
  nand2 gate860(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate861(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate862(.a(G416), .O(gate132inter7));
  inv1  gate863(.a(G417), .O(gate132inter8));
  nand2 gate864(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate865(.a(s_45), .b(gate132inter3), .O(gate132inter10));
  nor2  gate866(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate867(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate868(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1163(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1164(.a(gate136inter0), .b(s_88), .O(gate136inter1));
  and2  gate1165(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1166(.a(s_88), .O(gate136inter3));
  inv1  gate1167(.a(s_89), .O(gate136inter4));
  nand2 gate1168(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1169(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1170(.a(G424), .O(gate136inter7));
  inv1  gate1171(.a(G425), .O(gate136inter8));
  nand2 gate1172(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1173(.a(s_89), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1174(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1175(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1176(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1093(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1094(.a(gate138inter0), .b(s_78), .O(gate138inter1));
  and2  gate1095(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1096(.a(s_78), .O(gate138inter3));
  inv1  gate1097(.a(s_79), .O(gate138inter4));
  nand2 gate1098(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1099(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1100(.a(G432), .O(gate138inter7));
  inv1  gate1101(.a(G435), .O(gate138inter8));
  nand2 gate1102(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1103(.a(s_79), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1104(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1105(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1106(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1471(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1472(.a(gate140inter0), .b(s_132), .O(gate140inter1));
  and2  gate1473(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1474(.a(s_132), .O(gate140inter3));
  inv1  gate1475(.a(s_133), .O(gate140inter4));
  nand2 gate1476(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1477(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1478(.a(G444), .O(gate140inter7));
  inv1  gate1479(.a(G447), .O(gate140inter8));
  nand2 gate1480(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1481(.a(s_133), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1482(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1483(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1484(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1177(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1178(.a(gate145inter0), .b(s_90), .O(gate145inter1));
  and2  gate1179(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1180(.a(s_90), .O(gate145inter3));
  inv1  gate1181(.a(s_91), .O(gate145inter4));
  nand2 gate1182(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1183(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1184(.a(G474), .O(gate145inter7));
  inv1  gate1185(.a(G477), .O(gate145inter8));
  nand2 gate1186(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1187(.a(s_91), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1188(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1189(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1190(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1275(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1276(.a(gate146inter0), .b(s_104), .O(gate146inter1));
  and2  gate1277(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1278(.a(s_104), .O(gate146inter3));
  inv1  gate1279(.a(s_105), .O(gate146inter4));
  nand2 gate1280(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1281(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1282(.a(G480), .O(gate146inter7));
  inv1  gate1283(.a(G483), .O(gate146inter8));
  nand2 gate1284(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1285(.a(s_105), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1286(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1287(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1288(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate897(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate898(.a(gate148inter0), .b(s_50), .O(gate148inter1));
  and2  gate899(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate900(.a(s_50), .O(gate148inter3));
  inv1  gate901(.a(s_51), .O(gate148inter4));
  nand2 gate902(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate903(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate904(.a(G492), .O(gate148inter7));
  inv1  gate905(.a(G495), .O(gate148inter8));
  nand2 gate906(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate907(.a(s_51), .b(gate148inter3), .O(gate148inter10));
  nor2  gate908(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate909(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate910(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate1023(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1024(.a(gate149inter0), .b(s_68), .O(gate149inter1));
  and2  gate1025(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1026(.a(s_68), .O(gate149inter3));
  inv1  gate1027(.a(s_69), .O(gate149inter4));
  nand2 gate1028(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1029(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1030(.a(G498), .O(gate149inter7));
  inv1  gate1031(.a(G501), .O(gate149inter8));
  nand2 gate1032(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1033(.a(s_69), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1034(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1035(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1036(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2395(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2396(.a(gate151inter0), .b(s_264), .O(gate151inter1));
  and2  gate2397(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2398(.a(s_264), .O(gate151inter3));
  inv1  gate2399(.a(s_265), .O(gate151inter4));
  nand2 gate2400(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2401(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2402(.a(G510), .O(gate151inter7));
  inv1  gate2403(.a(G513), .O(gate151inter8));
  nand2 gate2404(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2405(.a(s_265), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2406(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2407(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2408(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate645(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate646(.a(gate154inter0), .b(s_14), .O(gate154inter1));
  and2  gate647(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate648(.a(s_14), .O(gate154inter3));
  inv1  gate649(.a(s_15), .O(gate154inter4));
  nand2 gate650(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate651(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate652(.a(G429), .O(gate154inter7));
  inv1  gate653(.a(G522), .O(gate154inter8));
  nand2 gate654(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate655(.a(s_15), .b(gate154inter3), .O(gate154inter10));
  nor2  gate656(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate657(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate658(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1219(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1220(.a(gate156inter0), .b(s_96), .O(gate156inter1));
  and2  gate1221(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1222(.a(s_96), .O(gate156inter3));
  inv1  gate1223(.a(s_97), .O(gate156inter4));
  nand2 gate1224(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1225(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1226(.a(G435), .O(gate156inter7));
  inv1  gate1227(.a(G525), .O(gate156inter8));
  nand2 gate1228(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1229(.a(s_97), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1230(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1231(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1232(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2283(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2284(.a(gate159inter0), .b(s_248), .O(gate159inter1));
  and2  gate2285(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2286(.a(s_248), .O(gate159inter3));
  inv1  gate2287(.a(s_249), .O(gate159inter4));
  nand2 gate2288(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2289(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2290(.a(G444), .O(gate159inter7));
  inv1  gate2291(.a(G531), .O(gate159inter8));
  nand2 gate2292(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2293(.a(s_249), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2294(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2295(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2296(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2437(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2438(.a(gate161inter0), .b(s_270), .O(gate161inter1));
  and2  gate2439(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2440(.a(s_270), .O(gate161inter3));
  inv1  gate2441(.a(s_271), .O(gate161inter4));
  nand2 gate2442(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2443(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2444(.a(G450), .O(gate161inter7));
  inv1  gate2445(.a(G534), .O(gate161inter8));
  nand2 gate2446(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2447(.a(s_271), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2448(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2449(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2450(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate2031(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2032(.a(gate162inter0), .b(s_212), .O(gate162inter1));
  and2  gate2033(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2034(.a(s_212), .O(gate162inter3));
  inv1  gate2035(.a(s_213), .O(gate162inter4));
  nand2 gate2036(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2037(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2038(.a(G453), .O(gate162inter7));
  inv1  gate2039(.a(G534), .O(gate162inter8));
  nand2 gate2040(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2041(.a(s_213), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2042(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2043(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2044(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1485(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1486(.a(gate164inter0), .b(s_134), .O(gate164inter1));
  and2  gate1487(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1488(.a(s_134), .O(gate164inter3));
  inv1  gate1489(.a(s_135), .O(gate164inter4));
  nand2 gate1490(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1491(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1492(.a(G459), .O(gate164inter7));
  inv1  gate1493(.a(G537), .O(gate164inter8));
  nand2 gate1494(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1495(.a(s_135), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1496(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1497(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1498(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate1905(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1906(.a(gate165inter0), .b(s_194), .O(gate165inter1));
  and2  gate1907(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1908(.a(s_194), .O(gate165inter3));
  inv1  gate1909(.a(s_195), .O(gate165inter4));
  nand2 gate1910(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1911(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1912(.a(G462), .O(gate165inter7));
  inv1  gate1913(.a(G540), .O(gate165inter8));
  nand2 gate1914(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1915(.a(s_195), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1916(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1917(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1918(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate827(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate828(.a(gate166inter0), .b(s_40), .O(gate166inter1));
  and2  gate829(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate830(.a(s_40), .O(gate166inter3));
  inv1  gate831(.a(s_41), .O(gate166inter4));
  nand2 gate832(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate833(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate834(.a(G465), .O(gate166inter7));
  inv1  gate835(.a(G540), .O(gate166inter8));
  nand2 gate836(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate837(.a(s_41), .b(gate166inter3), .O(gate166inter10));
  nor2  gate838(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate839(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate840(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1205(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1206(.a(gate168inter0), .b(s_94), .O(gate168inter1));
  and2  gate1207(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1208(.a(s_94), .O(gate168inter3));
  inv1  gate1209(.a(s_95), .O(gate168inter4));
  nand2 gate1210(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1211(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1212(.a(G471), .O(gate168inter7));
  inv1  gate1213(.a(G543), .O(gate168inter8));
  nand2 gate1214(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1215(.a(s_95), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1216(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1217(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1218(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2885(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2886(.a(gate169inter0), .b(s_334), .O(gate169inter1));
  and2  gate2887(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2888(.a(s_334), .O(gate169inter3));
  inv1  gate2889(.a(s_335), .O(gate169inter4));
  nand2 gate2890(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2891(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2892(.a(G474), .O(gate169inter7));
  inv1  gate2893(.a(G546), .O(gate169inter8));
  nand2 gate2894(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2895(.a(s_335), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2896(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2897(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2898(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate841(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate842(.a(gate172inter0), .b(s_42), .O(gate172inter1));
  and2  gate843(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate844(.a(s_42), .O(gate172inter3));
  inv1  gate845(.a(s_43), .O(gate172inter4));
  nand2 gate846(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate847(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate848(.a(G483), .O(gate172inter7));
  inv1  gate849(.a(G549), .O(gate172inter8));
  nand2 gate850(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate851(.a(s_43), .b(gate172inter3), .O(gate172inter10));
  nor2  gate852(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate853(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate854(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1457(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1458(.a(gate173inter0), .b(s_130), .O(gate173inter1));
  and2  gate1459(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1460(.a(s_130), .O(gate173inter3));
  inv1  gate1461(.a(s_131), .O(gate173inter4));
  nand2 gate1462(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1463(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1464(.a(G486), .O(gate173inter7));
  inv1  gate1465(.a(G552), .O(gate173inter8));
  nand2 gate1466(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1467(.a(s_131), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1468(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1469(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1470(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2017(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2018(.a(gate174inter0), .b(s_210), .O(gate174inter1));
  and2  gate2019(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2020(.a(s_210), .O(gate174inter3));
  inv1  gate2021(.a(s_211), .O(gate174inter4));
  nand2 gate2022(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2023(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2024(.a(G489), .O(gate174inter7));
  inv1  gate2025(.a(G552), .O(gate174inter8));
  nand2 gate2026(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2027(.a(s_211), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2028(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2029(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2030(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2745(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2746(.a(gate175inter0), .b(s_314), .O(gate175inter1));
  and2  gate2747(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2748(.a(s_314), .O(gate175inter3));
  inv1  gate2749(.a(s_315), .O(gate175inter4));
  nand2 gate2750(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2751(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2752(.a(G492), .O(gate175inter7));
  inv1  gate2753(.a(G555), .O(gate175inter8));
  nand2 gate2754(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2755(.a(s_315), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2756(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2757(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2758(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate911(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate912(.a(gate176inter0), .b(s_52), .O(gate176inter1));
  and2  gate913(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate914(.a(s_52), .O(gate176inter3));
  inv1  gate915(.a(s_53), .O(gate176inter4));
  nand2 gate916(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate917(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate918(.a(G495), .O(gate176inter7));
  inv1  gate919(.a(G555), .O(gate176inter8));
  nand2 gate920(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate921(.a(s_53), .b(gate176inter3), .O(gate176inter10));
  nor2  gate922(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate923(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate924(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2647(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2648(.a(gate179inter0), .b(s_300), .O(gate179inter1));
  and2  gate2649(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2650(.a(s_300), .O(gate179inter3));
  inv1  gate2651(.a(s_301), .O(gate179inter4));
  nand2 gate2652(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2653(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2654(.a(G504), .O(gate179inter7));
  inv1  gate2655(.a(G561), .O(gate179inter8));
  nand2 gate2656(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2657(.a(s_301), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2658(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2659(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2660(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate2927(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2928(.a(gate180inter0), .b(s_340), .O(gate180inter1));
  and2  gate2929(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2930(.a(s_340), .O(gate180inter3));
  inv1  gate2931(.a(s_341), .O(gate180inter4));
  nand2 gate2932(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2933(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2934(.a(G507), .O(gate180inter7));
  inv1  gate2935(.a(G561), .O(gate180inter8));
  nand2 gate2936(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2937(.a(s_341), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2938(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2939(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2940(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1751(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1752(.a(gate181inter0), .b(s_172), .O(gate181inter1));
  and2  gate1753(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1754(.a(s_172), .O(gate181inter3));
  inv1  gate1755(.a(s_173), .O(gate181inter4));
  nand2 gate1756(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1757(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1758(.a(G510), .O(gate181inter7));
  inv1  gate1759(.a(G564), .O(gate181inter8));
  nand2 gate1760(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1761(.a(s_173), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1762(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1763(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1764(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1345(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1346(.a(gate182inter0), .b(s_114), .O(gate182inter1));
  and2  gate1347(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1348(.a(s_114), .O(gate182inter3));
  inv1  gate1349(.a(s_115), .O(gate182inter4));
  nand2 gate1350(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1351(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1352(.a(G513), .O(gate182inter7));
  inv1  gate1353(.a(G564), .O(gate182inter8));
  nand2 gate1354(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1355(.a(s_115), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1356(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1357(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1358(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1919(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1920(.a(gate186inter0), .b(s_196), .O(gate186inter1));
  and2  gate1921(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1922(.a(s_196), .O(gate186inter3));
  inv1  gate1923(.a(s_197), .O(gate186inter4));
  nand2 gate1924(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1925(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1926(.a(G572), .O(gate186inter7));
  inv1  gate1927(.a(G573), .O(gate186inter8));
  nand2 gate1928(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1929(.a(s_197), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1930(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1931(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1932(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1051(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1052(.a(gate187inter0), .b(s_72), .O(gate187inter1));
  and2  gate1053(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1054(.a(s_72), .O(gate187inter3));
  inv1  gate1055(.a(s_73), .O(gate187inter4));
  nand2 gate1056(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1057(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1058(.a(G574), .O(gate187inter7));
  inv1  gate1059(.a(G575), .O(gate187inter8));
  nand2 gate1060(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1061(.a(s_73), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1062(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1063(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1064(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2521(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2522(.a(gate189inter0), .b(s_282), .O(gate189inter1));
  and2  gate2523(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2524(.a(s_282), .O(gate189inter3));
  inv1  gate2525(.a(s_283), .O(gate189inter4));
  nand2 gate2526(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2527(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2528(.a(G578), .O(gate189inter7));
  inv1  gate2529(.a(G579), .O(gate189inter8));
  nand2 gate2530(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2531(.a(s_283), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2532(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2533(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2534(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1849(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1850(.a(gate195inter0), .b(s_186), .O(gate195inter1));
  and2  gate1851(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1852(.a(s_186), .O(gate195inter3));
  inv1  gate1853(.a(s_187), .O(gate195inter4));
  nand2 gate1854(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1855(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1856(.a(G590), .O(gate195inter7));
  inv1  gate1857(.a(G591), .O(gate195inter8));
  nand2 gate1858(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1859(.a(s_187), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1860(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1861(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1862(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2451(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2452(.a(gate197inter0), .b(s_272), .O(gate197inter1));
  and2  gate2453(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2454(.a(s_272), .O(gate197inter3));
  inv1  gate2455(.a(s_273), .O(gate197inter4));
  nand2 gate2456(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2457(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2458(.a(G594), .O(gate197inter7));
  inv1  gate2459(.a(G595), .O(gate197inter8));
  nand2 gate2460(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2461(.a(s_273), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2462(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2463(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2464(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1541(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1542(.a(gate199inter0), .b(s_142), .O(gate199inter1));
  and2  gate1543(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1544(.a(s_142), .O(gate199inter3));
  inv1  gate1545(.a(s_143), .O(gate199inter4));
  nand2 gate1546(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1547(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1548(.a(G598), .O(gate199inter7));
  inv1  gate1549(.a(G599), .O(gate199inter8));
  nand2 gate1550(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1551(.a(s_143), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1552(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1553(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1554(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1149(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1150(.a(gate200inter0), .b(s_86), .O(gate200inter1));
  and2  gate1151(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1152(.a(s_86), .O(gate200inter3));
  inv1  gate1153(.a(s_87), .O(gate200inter4));
  nand2 gate1154(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1155(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1156(.a(G600), .O(gate200inter7));
  inv1  gate1157(.a(G601), .O(gate200inter8));
  nand2 gate1158(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1159(.a(s_87), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1160(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1161(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1162(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1947(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1948(.a(gate201inter0), .b(s_200), .O(gate201inter1));
  and2  gate1949(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1950(.a(s_200), .O(gate201inter3));
  inv1  gate1951(.a(s_201), .O(gate201inter4));
  nand2 gate1952(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1953(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1954(.a(G602), .O(gate201inter7));
  inv1  gate1955(.a(G607), .O(gate201inter8));
  nand2 gate1956(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1957(.a(s_201), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1958(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1959(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1960(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate561(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate562(.a(gate202inter0), .b(s_2), .O(gate202inter1));
  and2  gate563(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate564(.a(s_2), .O(gate202inter3));
  inv1  gate565(.a(s_3), .O(gate202inter4));
  nand2 gate566(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate567(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate568(.a(G612), .O(gate202inter7));
  inv1  gate569(.a(G617), .O(gate202inter8));
  nand2 gate570(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate571(.a(s_3), .b(gate202inter3), .O(gate202inter10));
  nor2  gate572(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate573(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate574(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2535(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2536(.a(gate205inter0), .b(s_284), .O(gate205inter1));
  and2  gate2537(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2538(.a(s_284), .O(gate205inter3));
  inv1  gate2539(.a(s_285), .O(gate205inter4));
  nand2 gate2540(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2541(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2542(.a(G622), .O(gate205inter7));
  inv1  gate2543(.a(G627), .O(gate205inter8));
  nand2 gate2544(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2545(.a(s_285), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2546(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2547(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2548(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2353(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2354(.a(gate211inter0), .b(s_258), .O(gate211inter1));
  and2  gate2355(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2356(.a(s_258), .O(gate211inter3));
  inv1  gate2357(.a(s_259), .O(gate211inter4));
  nand2 gate2358(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2359(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2360(.a(G612), .O(gate211inter7));
  inv1  gate2361(.a(G669), .O(gate211inter8));
  nand2 gate2362(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2363(.a(s_259), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2364(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2365(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2366(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2227(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2228(.a(gate212inter0), .b(s_240), .O(gate212inter1));
  and2  gate2229(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2230(.a(s_240), .O(gate212inter3));
  inv1  gate2231(.a(s_241), .O(gate212inter4));
  nand2 gate2232(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2233(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2234(.a(G617), .O(gate212inter7));
  inv1  gate2235(.a(G669), .O(gate212inter8));
  nand2 gate2236(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2237(.a(s_241), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2238(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2239(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2240(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1639(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1640(.a(gate214inter0), .b(s_156), .O(gate214inter1));
  and2  gate1641(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1642(.a(s_156), .O(gate214inter3));
  inv1  gate1643(.a(s_157), .O(gate214inter4));
  nand2 gate1644(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1645(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1646(.a(G612), .O(gate214inter7));
  inv1  gate1647(.a(G672), .O(gate214inter8));
  nand2 gate1648(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1649(.a(s_157), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1650(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1651(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1652(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1009(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1010(.a(gate215inter0), .b(s_66), .O(gate215inter1));
  and2  gate1011(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1012(.a(s_66), .O(gate215inter3));
  inv1  gate1013(.a(s_67), .O(gate215inter4));
  nand2 gate1014(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1015(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1016(.a(G607), .O(gate215inter7));
  inv1  gate1017(.a(G675), .O(gate215inter8));
  nand2 gate1018(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1019(.a(s_67), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1020(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1021(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1022(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1807(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1808(.a(gate219inter0), .b(s_180), .O(gate219inter1));
  and2  gate1809(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1810(.a(s_180), .O(gate219inter3));
  inv1  gate1811(.a(s_181), .O(gate219inter4));
  nand2 gate1812(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1813(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1814(.a(G632), .O(gate219inter7));
  inv1  gate1815(.a(G681), .O(gate219inter8));
  nand2 gate1816(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1817(.a(s_181), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1818(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1819(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1820(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2199(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2200(.a(gate222inter0), .b(s_236), .O(gate222inter1));
  and2  gate2201(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2202(.a(s_236), .O(gate222inter3));
  inv1  gate2203(.a(s_237), .O(gate222inter4));
  nand2 gate2204(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2205(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2206(.a(G632), .O(gate222inter7));
  inv1  gate2207(.a(G684), .O(gate222inter8));
  nand2 gate2208(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2209(.a(s_237), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2210(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2211(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2212(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2759(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2760(.a(gate224inter0), .b(s_316), .O(gate224inter1));
  and2  gate2761(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2762(.a(s_316), .O(gate224inter3));
  inv1  gate2763(.a(s_317), .O(gate224inter4));
  nand2 gate2764(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2765(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2766(.a(G637), .O(gate224inter7));
  inv1  gate2767(.a(G687), .O(gate224inter8));
  nand2 gate2768(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2769(.a(s_317), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2770(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2771(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2772(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate939(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate940(.a(gate227inter0), .b(s_56), .O(gate227inter1));
  and2  gate941(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate942(.a(s_56), .O(gate227inter3));
  inv1  gate943(.a(s_57), .O(gate227inter4));
  nand2 gate944(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate945(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate946(.a(G694), .O(gate227inter7));
  inv1  gate947(.a(G695), .O(gate227inter8));
  nand2 gate948(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate949(.a(s_57), .b(gate227inter3), .O(gate227inter10));
  nor2  gate950(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate951(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate952(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2115(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2116(.a(gate232inter0), .b(s_224), .O(gate232inter1));
  and2  gate2117(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2118(.a(s_224), .O(gate232inter3));
  inv1  gate2119(.a(s_225), .O(gate232inter4));
  nand2 gate2120(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2121(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2122(.a(G704), .O(gate232inter7));
  inv1  gate2123(.a(G705), .O(gate232inter8));
  nand2 gate2124(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2125(.a(s_225), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2126(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2127(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2128(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate743(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate744(.a(gate235inter0), .b(s_28), .O(gate235inter1));
  and2  gate745(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate746(.a(s_28), .O(gate235inter3));
  inv1  gate747(.a(s_29), .O(gate235inter4));
  nand2 gate748(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate749(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate750(.a(G248), .O(gate235inter7));
  inv1  gate751(.a(G724), .O(gate235inter8));
  nand2 gate752(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate753(.a(s_29), .b(gate235inter3), .O(gate235inter10));
  nor2  gate754(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate755(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate756(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2423(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2424(.a(gate236inter0), .b(s_268), .O(gate236inter1));
  and2  gate2425(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2426(.a(s_268), .O(gate236inter3));
  inv1  gate2427(.a(s_269), .O(gate236inter4));
  nand2 gate2428(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2429(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2430(.a(G251), .O(gate236inter7));
  inv1  gate2431(.a(G727), .O(gate236inter8));
  nand2 gate2432(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2433(.a(s_269), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2434(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2435(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2436(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate2255(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2256(.a(gate237inter0), .b(s_244), .O(gate237inter1));
  and2  gate2257(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2258(.a(s_244), .O(gate237inter3));
  inv1  gate2259(.a(s_245), .O(gate237inter4));
  nand2 gate2260(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2261(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2262(.a(G254), .O(gate237inter7));
  inv1  gate2263(.a(G706), .O(gate237inter8));
  nand2 gate2264(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2265(.a(s_245), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2266(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2267(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2268(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1597(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1598(.a(gate243inter0), .b(s_150), .O(gate243inter1));
  and2  gate1599(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1600(.a(s_150), .O(gate243inter3));
  inv1  gate1601(.a(s_151), .O(gate243inter4));
  nand2 gate1602(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1603(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1604(.a(G245), .O(gate243inter7));
  inv1  gate1605(.a(G733), .O(gate243inter8));
  nand2 gate1606(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1607(.a(s_151), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1608(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1609(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1610(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate953(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate954(.a(gate246inter0), .b(s_58), .O(gate246inter1));
  and2  gate955(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate956(.a(s_58), .O(gate246inter3));
  inv1  gate957(.a(s_59), .O(gate246inter4));
  nand2 gate958(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate959(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate960(.a(G724), .O(gate246inter7));
  inv1  gate961(.a(G736), .O(gate246inter8));
  nand2 gate962(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate963(.a(s_59), .b(gate246inter3), .O(gate246inter10));
  nor2  gate964(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate965(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate966(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate575(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate576(.a(gate248inter0), .b(s_4), .O(gate248inter1));
  and2  gate577(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate578(.a(s_4), .O(gate248inter3));
  inv1  gate579(.a(s_5), .O(gate248inter4));
  nand2 gate580(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate581(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate582(.a(G727), .O(gate248inter7));
  inv1  gate583(.a(G739), .O(gate248inter8));
  nand2 gate584(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate585(.a(s_5), .b(gate248inter3), .O(gate248inter10));
  nor2  gate586(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate587(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate588(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1583(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1584(.a(gate253inter0), .b(s_148), .O(gate253inter1));
  and2  gate1585(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1586(.a(s_148), .O(gate253inter3));
  inv1  gate1587(.a(s_149), .O(gate253inter4));
  nand2 gate1588(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1589(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1590(.a(G260), .O(gate253inter7));
  inv1  gate1591(.a(G748), .O(gate253inter8));
  nand2 gate1592(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1593(.a(s_149), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1594(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1595(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1596(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate757(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate758(.a(gate254inter0), .b(s_30), .O(gate254inter1));
  and2  gate759(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate760(.a(s_30), .O(gate254inter3));
  inv1  gate761(.a(s_31), .O(gate254inter4));
  nand2 gate762(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate763(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate764(.a(G712), .O(gate254inter7));
  inv1  gate765(.a(G748), .O(gate254inter8));
  nand2 gate766(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate767(.a(s_31), .b(gate254inter3), .O(gate254inter10));
  nor2  gate768(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate769(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate770(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate617(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate618(.a(gate258inter0), .b(s_10), .O(gate258inter1));
  and2  gate619(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate620(.a(s_10), .O(gate258inter3));
  inv1  gate621(.a(s_11), .O(gate258inter4));
  nand2 gate622(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate623(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate624(.a(G756), .O(gate258inter7));
  inv1  gate625(.a(G757), .O(gate258inter8));
  nand2 gate626(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate627(.a(s_11), .b(gate258inter3), .O(gate258inter10));
  nor2  gate628(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate629(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate630(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2367(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2368(.a(gate262inter0), .b(s_260), .O(gate262inter1));
  and2  gate2369(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2370(.a(s_260), .O(gate262inter3));
  inv1  gate2371(.a(s_261), .O(gate262inter4));
  nand2 gate2372(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2373(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2374(.a(G764), .O(gate262inter7));
  inv1  gate2375(.a(G765), .O(gate262inter8));
  nand2 gate2376(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2377(.a(s_261), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2378(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2379(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2380(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2073(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2074(.a(gate263inter0), .b(s_218), .O(gate263inter1));
  and2  gate2075(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2076(.a(s_218), .O(gate263inter3));
  inv1  gate2077(.a(s_219), .O(gate263inter4));
  nand2 gate2078(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2079(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2080(.a(G766), .O(gate263inter7));
  inv1  gate2081(.a(G767), .O(gate263inter8));
  nand2 gate2082(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2083(.a(s_219), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2084(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2085(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2086(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate547(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate548(.a(gate264inter0), .b(s_0), .O(gate264inter1));
  and2  gate549(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate550(.a(s_0), .O(gate264inter3));
  inv1  gate551(.a(s_1), .O(gate264inter4));
  nand2 gate552(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate553(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate554(.a(G768), .O(gate264inter7));
  inv1  gate555(.a(G769), .O(gate264inter8));
  nand2 gate556(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate557(.a(s_1), .b(gate264inter3), .O(gate264inter10));
  nor2  gate558(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate559(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate560(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2171(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2172(.a(gate267inter0), .b(s_232), .O(gate267inter1));
  and2  gate2173(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2174(.a(s_232), .O(gate267inter3));
  inv1  gate2175(.a(s_233), .O(gate267inter4));
  nand2 gate2176(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2177(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2178(.a(G648), .O(gate267inter7));
  inv1  gate2179(.a(G776), .O(gate267inter8));
  nand2 gate2180(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2181(.a(s_233), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2182(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2183(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2184(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1555(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1556(.a(gate268inter0), .b(s_144), .O(gate268inter1));
  and2  gate1557(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1558(.a(s_144), .O(gate268inter3));
  inv1  gate1559(.a(s_145), .O(gate268inter4));
  nand2 gate1560(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1561(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1562(.a(G651), .O(gate268inter7));
  inv1  gate1563(.a(G779), .O(gate268inter8));
  nand2 gate1564(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1565(.a(s_145), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1566(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1567(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1568(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1709(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1710(.a(gate270inter0), .b(s_166), .O(gate270inter1));
  and2  gate1711(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1712(.a(s_166), .O(gate270inter3));
  inv1  gate1713(.a(s_167), .O(gate270inter4));
  nand2 gate1714(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1715(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1716(.a(G657), .O(gate270inter7));
  inv1  gate1717(.a(G785), .O(gate270inter8));
  nand2 gate1718(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1719(.a(s_167), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1720(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1721(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1722(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate925(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate926(.a(gate272inter0), .b(s_54), .O(gate272inter1));
  and2  gate927(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate928(.a(s_54), .O(gate272inter3));
  inv1  gate929(.a(s_55), .O(gate272inter4));
  nand2 gate930(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate931(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate932(.a(G663), .O(gate272inter7));
  inv1  gate933(.a(G791), .O(gate272inter8));
  nand2 gate934(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate935(.a(s_55), .b(gate272inter3), .O(gate272inter10));
  nor2  gate936(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate937(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate938(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1373(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1374(.a(gate274inter0), .b(s_118), .O(gate274inter1));
  and2  gate1375(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1376(.a(s_118), .O(gate274inter3));
  inv1  gate1377(.a(s_119), .O(gate274inter4));
  nand2 gate1378(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1379(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1380(.a(G770), .O(gate274inter7));
  inv1  gate1381(.a(G794), .O(gate274inter8));
  nand2 gate1382(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1383(.a(s_119), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1384(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1385(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1386(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1443(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1444(.a(gate277inter0), .b(s_128), .O(gate277inter1));
  and2  gate1445(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1446(.a(s_128), .O(gate277inter3));
  inv1  gate1447(.a(s_129), .O(gate277inter4));
  nand2 gate1448(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1449(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1450(.a(G648), .O(gate277inter7));
  inv1  gate1451(.a(G800), .O(gate277inter8));
  nand2 gate1452(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1453(.a(s_129), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1454(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1455(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1456(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2143(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2144(.a(gate279inter0), .b(s_228), .O(gate279inter1));
  and2  gate2145(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2146(.a(s_228), .O(gate279inter3));
  inv1  gate2147(.a(s_229), .O(gate279inter4));
  nand2 gate2148(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2149(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2150(.a(G651), .O(gate279inter7));
  inv1  gate2151(.a(G803), .O(gate279inter8));
  nand2 gate2152(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2153(.a(s_229), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2154(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2155(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2156(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate589(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate590(.a(gate281inter0), .b(s_6), .O(gate281inter1));
  and2  gate591(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate592(.a(s_6), .O(gate281inter3));
  inv1  gate593(.a(s_7), .O(gate281inter4));
  nand2 gate594(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate595(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate596(.a(G654), .O(gate281inter7));
  inv1  gate597(.a(G806), .O(gate281inter8));
  nand2 gate598(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate599(.a(s_7), .b(gate281inter3), .O(gate281inter10));
  nor2  gate600(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate601(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate602(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2493(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2494(.a(gate285inter0), .b(s_278), .O(gate285inter1));
  and2  gate2495(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2496(.a(s_278), .O(gate285inter3));
  inv1  gate2497(.a(s_279), .O(gate285inter4));
  nand2 gate2498(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2499(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2500(.a(G660), .O(gate285inter7));
  inv1  gate2501(.a(G812), .O(gate285inter8));
  nand2 gate2502(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2503(.a(s_279), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2504(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2505(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2506(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate967(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate968(.a(gate286inter0), .b(s_60), .O(gate286inter1));
  and2  gate969(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate970(.a(s_60), .O(gate286inter3));
  inv1  gate971(.a(s_61), .O(gate286inter4));
  nand2 gate972(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate973(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate974(.a(G788), .O(gate286inter7));
  inv1  gate975(.a(G812), .O(gate286inter8));
  nand2 gate976(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate977(.a(s_61), .b(gate286inter3), .O(gate286inter10));
  nor2  gate978(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate979(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate980(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2577(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2578(.a(gate287inter0), .b(s_290), .O(gate287inter1));
  and2  gate2579(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2580(.a(s_290), .O(gate287inter3));
  inv1  gate2581(.a(s_291), .O(gate287inter4));
  nand2 gate2582(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2583(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2584(.a(G663), .O(gate287inter7));
  inv1  gate2585(.a(G815), .O(gate287inter8));
  nand2 gate2586(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2587(.a(s_291), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2588(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2589(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2590(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1765(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1766(.a(gate289inter0), .b(s_174), .O(gate289inter1));
  and2  gate1767(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1768(.a(s_174), .O(gate289inter3));
  inv1  gate1769(.a(s_175), .O(gate289inter4));
  nand2 gate1770(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1771(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1772(.a(G818), .O(gate289inter7));
  inv1  gate1773(.a(G819), .O(gate289inter8));
  nand2 gate1774(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1775(.a(s_175), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1776(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1777(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1778(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1989(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1990(.a(gate292inter0), .b(s_206), .O(gate292inter1));
  and2  gate1991(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1992(.a(s_206), .O(gate292inter3));
  inv1  gate1993(.a(s_207), .O(gate292inter4));
  nand2 gate1994(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1995(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1996(.a(G824), .O(gate292inter7));
  inv1  gate1997(.a(G825), .O(gate292inter8));
  nand2 gate1998(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1999(.a(s_207), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2000(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2001(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2002(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1961(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1962(.a(gate395inter0), .b(s_202), .O(gate395inter1));
  and2  gate1963(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1964(.a(s_202), .O(gate395inter3));
  inv1  gate1965(.a(s_203), .O(gate395inter4));
  nand2 gate1966(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1967(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1968(.a(G9), .O(gate395inter7));
  inv1  gate1969(.a(G1060), .O(gate395inter8));
  nand2 gate1970(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1971(.a(s_203), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1972(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1973(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1974(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate2479(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2480(.a(gate399inter0), .b(s_276), .O(gate399inter1));
  and2  gate2481(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2482(.a(s_276), .O(gate399inter3));
  inv1  gate2483(.a(s_277), .O(gate399inter4));
  nand2 gate2484(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2485(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2486(.a(G13), .O(gate399inter7));
  inv1  gate2487(.a(G1072), .O(gate399inter8));
  nand2 gate2488(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2489(.a(s_277), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2490(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2491(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2492(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2605(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2606(.a(gate404inter0), .b(s_294), .O(gate404inter1));
  and2  gate2607(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2608(.a(s_294), .O(gate404inter3));
  inv1  gate2609(.a(s_295), .O(gate404inter4));
  nand2 gate2610(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2611(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2612(.a(G18), .O(gate404inter7));
  inv1  gate2613(.a(G1087), .O(gate404inter8));
  nand2 gate2614(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2615(.a(s_295), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2616(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2617(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2618(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate2857(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2858(.a(gate405inter0), .b(s_330), .O(gate405inter1));
  and2  gate2859(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2860(.a(s_330), .O(gate405inter3));
  inv1  gate2861(.a(s_331), .O(gate405inter4));
  nand2 gate2862(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2863(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2864(.a(G19), .O(gate405inter7));
  inv1  gate2865(.a(G1090), .O(gate405inter8));
  nand2 gate2866(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2867(.a(s_331), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2868(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2869(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2870(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2689(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2690(.a(gate411inter0), .b(s_306), .O(gate411inter1));
  and2  gate2691(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2692(.a(s_306), .O(gate411inter3));
  inv1  gate2693(.a(s_307), .O(gate411inter4));
  nand2 gate2694(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2695(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2696(.a(G25), .O(gate411inter7));
  inv1  gate2697(.a(G1108), .O(gate411inter8));
  nand2 gate2698(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2699(.a(s_307), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2700(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2701(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2702(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2213(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2214(.a(gate412inter0), .b(s_238), .O(gate412inter1));
  and2  gate2215(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2216(.a(s_238), .O(gate412inter3));
  inv1  gate2217(.a(s_239), .O(gate412inter4));
  nand2 gate2218(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2219(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2220(.a(G26), .O(gate412inter7));
  inv1  gate2221(.a(G1111), .O(gate412inter8));
  nand2 gate2222(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2223(.a(s_239), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2224(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2225(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2226(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate813(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate814(.a(gate413inter0), .b(s_38), .O(gate413inter1));
  and2  gate815(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate816(.a(s_38), .O(gate413inter3));
  inv1  gate817(.a(s_39), .O(gate413inter4));
  nand2 gate818(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate819(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate820(.a(G27), .O(gate413inter7));
  inv1  gate821(.a(G1114), .O(gate413inter8));
  nand2 gate822(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate823(.a(s_39), .b(gate413inter3), .O(gate413inter10));
  nor2  gate824(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate825(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate826(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2045(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2046(.a(gate418inter0), .b(s_214), .O(gate418inter1));
  and2  gate2047(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2048(.a(s_214), .O(gate418inter3));
  inv1  gate2049(.a(s_215), .O(gate418inter4));
  nand2 gate2050(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2051(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2052(.a(G32), .O(gate418inter7));
  inv1  gate2053(.a(G1129), .O(gate418inter8));
  nand2 gate2054(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2055(.a(s_215), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2056(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2057(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2058(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1079(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1080(.a(gate421inter0), .b(s_76), .O(gate421inter1));
  and2  gate1081(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1082(.a(s_76), .O(gate421inter3));
  inv1  gate1083(.a(s_77), .O(gate421inter4));
  nand2 gate1084(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1085(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1086(.a(G2), .O(gate421inter7));
  inv1  gate1087(.a(G1135), .O(gate421inter8));
  nand2 gate1088(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1089(.a(s_77), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1090(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1091(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1092(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1513(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1514(.a(gate424inter0), .b(s_138), .O(gate424inter1));
  and2  gate1515(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1516(.a(s_138), .O(gate424inter3));
  inv1  gate1517(.a(s_139), .O(gate424inter4));
  nand2 gate1518(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1519(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1520(.a(G1042), .O(gate424inter7));
  inv1  gate1521(.a(G1138), .O(gate424inter8));
  nand2 gate1522(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1523(.a(s_139), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1524(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1525(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1526(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate673(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate674(.a(gate431inter0), .b(s_18), .O(gate431inter1));
  and2  gate675(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate676(.a(s_18), .O(gate431inter3));
  inv1  gate677(.a(s_19), .O(gate431inter4));
  nand2 gate678(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate679(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate680(.a(G7), .O(gate431inter7));
  inv1  gate681(.a(G1150), .O(gate431inter8));
  nand2 gate682(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate683(.a(s_19), .b(gate431inter3), .O(gate431inter10));
  nor2  gate684(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate685(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate686(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1779(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1780(.a(gate432inter0), .b(s_176), .O(gate432inter1));
  and2  gate1781(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1782(.a(s_176), .O(gate432inter3));
  inv1  gate1783(.a(s_177), .O(gate432inter4));
  nand2 gate1784(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1785(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1786(.a(G1054), .O(gate432inter7));
  inv1  gate1787(.a(G1150), .O(gate432inter8));
  nand2 gate1788(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1789(.a(s_177), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1790(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1791(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1792(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2311(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2312(.a(gate433inter0), .b(s_252), .O(gate433inter1));
  and2  gate2313(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2314(.a(s_252), .O(gate433inter3));
  inv1  gate2315(.a(s_253), .O(gate433inter4));
  nand2 gate2316(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2317(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2318(.a(G8), .O(gate433inter7));
  inv1  gate2319(.a(G1153), .O(gate433inter8));
  nand2 gate2320(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2321(.a(s_253), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2322(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2323(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2324(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate2563(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2564(.a(gate434inter0), .b(s_288), .O(gate434inter1));
  and2  gate2565(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2566(.a(s_288), .O(gate434inter3));
  inv1  gate2567(.a(s_289), .O(gate434inter4));
  nand2 gate2568(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2569(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2570(.a(G1057), .O(gate434inter7));
  inv1  gate2571(.a(G1153), .O(gate434inter8));
  nand2 gate2572(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2573(.a(s_289), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2574(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2575(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2576(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2241(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2242(.a(gate438inter0), .b(s_242), .O(gate438inter1));
  and2  gate2243(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2244(.a(s_242), .O(gate438inter3));
  inv1  gate2245(.a(s_243), .O(gate438inter4));
  nand2 gate2246(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2247(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2248(.a(G1063), .O(gate438inter7));
  inv1  gate2249(.a(G1159), .O(gate438inter8));
  nand2 gate2250(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2251(.a(s_243), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2252(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2253(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2254(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate687(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate688(.a(gate439inter0), .b(s_20), .O(gate439inter1));
  and2  gate689(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate690(.a(s_20), .O(gate439inter3));
  inv1  gate691(.a(s_21), .O(gate439inter4));
  nand2 gate692(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate693(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate694(.a(G11), .O(gate439inter7));
  inv1  gate695(.a(G1162), .O(gate439inter8));
  nand2 gate696(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate697(.a(s_21), .b(gate439inter3), .O(gate439inter10));
  nor2  gate698(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate699(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate700(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1611(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1612(.a(gate440inter0), .b(s_152), .O(gate440inter1));
  and2  gate1613(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1614(.a(s_152), .O(gate440inter3));
  inv1  gate1615(.a(s_153), .O(gate440inter4));
  nand2 gate1616(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1617(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1618(.a(G1066), .O(gate440inter7));
  inv1  gate1619(.a(G1162), .O(gate440inter8));
  nand2 gate1620(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1621(.a(s_153), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1622(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1623(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1624(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1835(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1836(.a(gate445inter0), .b(s_184), .O(gate445inter1));
  and2  gate1837(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1838(.a(s_184), .O(gate445inter3));
  inv1  gate1839(.a(s_185), .O(gate445inter4));
  nand2 gate1840(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1841(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1842(.a(G14), .O(gate445inter7));
  inv1  gate1843(.a(G1171), .O(gate445inter8));
  nand2 gate1844(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1845(.a(s_185), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1846(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1847(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1848(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1863(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1864(.a(gate449inter0), .b(s_188), .O(gate449inter1));
  and2  gate1865(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1866(.a(s_188), .O(gate449inter3));
  inv1  gate1867(.a(s_189), .O(gate449inter4));
  nand2 gate1868(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1869(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1870(.a(G16), .O(gate449inter7));
  inv1  gate1871(.a(G1177), .O(gate449inter8));
  nand2 gate1872(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1873(.a(s_189), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1874(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1875(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1876(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1247(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1248(.a(gate450inter0), .b(s_100), .O(gate450inter1));
  and2  gate1249(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1250(.a(s_100), .O(gate450inter3));
  inv1  gate1251(.a(s_101), .O(gate450inter4));
  nand2 gate1252(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1253(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1254(.a(G1081), .O(gate450inter7));
  inv1  gate1255(.a(G1177), .O(gate450inter8));
  nand2 gate1256(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1257(.a(s_101), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1258(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1259(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1260(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1387(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1388(.a(gate453inter0), .b(s_120), .O(gate453inter1));
  and2  gate1389(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1390(.a(s_120), .O(gate453inter3));
  inv1  gate1391(.a(s_121), .O(gate453inter4));
  nand2 gate1392(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1393(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1394(.a(G18), .O(gate453inter7));
  inv1  gate1395(.a(G1183), .O(gate453inter8));
  nand2 gate1396(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1397(.a(s_121), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1398(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1399(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1400(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1877(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1878(.a(gate457inter0), .b(s_190), .O(gate457inter1));
  and2  gate1879(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1880(.a(s_190), .O(gate457inter3));
  inv1  gate1881(.a(s_191), .O(gate457inter4));
  nand2 gate1882(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1883(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1884(.a(G20), .O(gate457inter7));
  inv1  gate1885(.a(G1189), .O(gate457inter8));
  nand2 gate1886(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1887(.a(s_191), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1888(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1889(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1890(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1975(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1976(.a(gate458inter0), .b(s_204), .O(gate458inter1));
  and2  gate1977(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1978(.a(s_204), .O(gate458inter3));
  inv1  gate1979(.a(s_205), .O(gate458inter4));
  nand2 gate1980(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1981(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1982(.a(G1093), .O(gate458inter7));
  inv1  gate1983(.a(G1189), .O(gate458inter8));
  nand2 gate1984(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1985(.a(s_205), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1986(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1987(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1988(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1289(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1290(.a(gate459inter0), .b(s_106), .O(gate459inter1));
  and2  gate1291(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1292(.a(s_106), .O(gate459inter3));
  inv1  gate1293(.a(s_107), .O(gate459inter4));
  nand2 gate1294(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1295(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1296(.a(G21), .O(gate459inter7));
  inv1  gate1297(.a(G1192), .O(gate459inter8));
  nand2 gate1298(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1299(.a(s_107), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1300(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1301(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1302(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2913(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2914(.a(gate461inter0), .b(s_338), .O(gate461inter1));
  and2  gate2915(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2916(.a(s_338), .O(gate461inter3));
  inv1  gate2917(.a(s_339), .O(gate461inter4));
  nand2 gate2918(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2919(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2920(.a(G22), .O(gate461inter7));
  inv1  gate2921(.a(G1195), .O(gate461inter8));
  nand2 gate2922(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2923(.a(s_339), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2924(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2925(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2926(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1359(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1360(.a(gate466inter0), .b(s_116), .O(gate466inter1));
  and2  gate1361(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1362(.a(s_116), .O(gate466inter3));
  inv1  gate1363(.a(s_117), .O(gate466inter4));
  nand2 gate1364(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1365(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1366(.a(G1105), .O(gate466inter7));
  inv1  gate1367(.a(G1201), .O(gate466inter8));
  nand2 gate1368(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1369(.a(s_117), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1370(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1371(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1372(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate2829(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2830(.a(gate468inter0), .b(s_326), .O(gate468inter1));
  and2  gate2831(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2832(.a(s_326), .O(gate468inter3));
  inv1  gate2833(.a(s_327), .O(gate468inter4));
  nand2 gate2834(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2835(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2836(.a(G1108), .O(gate468inter7));
  inv1  gate2837(.a(G1204), .O(gate468inter8));
  nand2 gate2838(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2839(.a(s_327), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2840(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2841(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2842(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2129(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2130(.a(gate471inter0), .b(s_226), .O(gate471inter1));
  and2  gate2131(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2132(.a(s_226), .O(gate471inter3));
  inv1  gate2133(.a(s_227), .O(gate471inter4));
  nand2 gate2134(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2135(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2136(.a(G27), .O(gate471inter7));
  inv1  gate2137(.a(G1210), .O(gate471inter8));
  nand2 gate2138(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2139(.a(s_227), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2140(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2141(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2142(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate883(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate884(.a(gate472inter0), .b(s_48), .O(gate472inter1));
  and2  gate885(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate886(.a(s_48), .O(gate472inter3));
  inv1  gate887(.a(s_49), .O(gate472inter4));
  nand2 gate888(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate889(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate890(.a(G1114), .O(gate472inter7));
  inv1  gate891(.a(G1210), .O(gate472inter8));
  nand2 gate892(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate893(.a(s_49), .b(gate472inter3), .O(gate472inter10));
  nor2  gate894(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate895(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate896(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2661(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2662(.a(gate474inter0), .b(s_302), .O(gate474inter1));
  and2  gate2663(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2664(.a(s_302), .O(gate474inter3));
  inv1  gate2665(.a(s_303), .O(gate474inter4));
  nand2 gate2666(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2667(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2668(.a(G1117), .O(gate474inter7));
  inv1  gate2669(.a(G1213), .O(gate474inter8));
  nand2 gate2670(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2671(.a(s_303), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2672(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2673(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2674(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate2731(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2732(.a(gate475inter0), .b(s_312), .O(gate475inter1));
  and2  gate2733(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2734(.a(s_312), .O(gate475inter3));
  inv1  gate2735(.a(s_313), .O(gate475inter4));
  nand2 gate2736(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2737(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2738(.a(G29), .O(gate475inter7));
  inv1  gate2739(.a(G1216), .O(gate475inter8));
  nand2 gate2740(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2741(.a(s_313), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2742(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2743(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2744(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2325(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2326(.a(gate476inter0), .b(s_254), .O(gate476inter1));
  and2  gate2327(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2328(.a(s_254), .O(gate476inter3));
  inv1  gate2329(.a(s_255), .O(gate476inter4));
  nand2 gate2330(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2331(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2332(.a(G1120), .O(gate476inter7));
  inv1  gate2333(.a(G1216), .O(gate476inter8));
  nand2 gate2334(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2335(.a(s_255), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2336(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2337(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2338(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate2409(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2410(.a(gate477inter0), .b(s_266), .O(gate477inter1));
  and2  gate2411(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2412(.a(s_266), .O(gate477inter3));
  inv1  gate2413(.a(s_267), .O(gate477inter4));
  nand2 gate2414(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2415(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2416(.a(G30), .O(gate477inter7));
  inv1  gate2417(.a(G1219), .O(gate477inter8));
  nand2 gate2418(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2419(.a(s_267), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2420(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2421(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2422(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate701(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate702(.a(gate481inter0), .b(s_22), .O(gate481inter1));
  and2  gate703(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate704(.a(s_22), .O(gate481inter3));
  inv1  gate705(.a(s_23), .O(gate481inter4));
  nand2 gate706(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate707(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate708(.a(G32), .O(gate481inter7));
  inv1  gate709(.a(G1225), .O(gate481inter8));
  nand2 gate710(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate711(.a(s_23), .b(gate481inter3), .O(gate481inter10));
  nor2  gate712(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate713(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate714(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1317(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1318(.a(gate485inter0), .b(s_110), .O(gate485inter1));
  and2  gate1319(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1320(.a(s_110), .O(gate485inter3));
  inv1  gate1321(.a(s_111), .O(gate485inter4));
  nand2 gate1322(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1323(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1324(.a(G1232), .O(gate485inter7));
  inv1  gate1325(.a(G1233), .O(gate485inter8));
  nand2 gate1326(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1327(.a(s_111), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1328(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1329(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1330(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1191(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1192(.a(gate486inter0), .b(s_92), .O(gate486inter1));
  and2  gate1193(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1194(.a(s_92), .O(gate486inter3));
  inv1  gate1195(.a(s_93), .O(gate486inter4));
  nand2 gate1196(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1197(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1198(.a(G1234), .O(gate486inter7));
  inv1  gate1199(.a(G1235), .O(gate486inter8));
  nand2 gate1200(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1201(.a(s_93), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1202(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1203(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1204(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2843(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2844(.a(gate487inter0), .b(s_328), .O(gate487inter1));
  and2  gate2845(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2846(.a(s_328), .O(gate487inter3));
  inv1  gate2847(.a(s_329), .O(gate487inter4));
  nand2 gate2848(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2849(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2850(.a(G1236), .O(gate487inter7));
  inv1  gate2851(.a(G1237), .O(gate487inter8));
  nand2 gate2852(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2853(.a(s_329), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2854(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2855(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2856(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1429(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1430(.a(gate488inter0), .b(s_126), .O(gate488inter1));
  and2  gate1431(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1432(.a(s_126), .O(gate488inter3));
  inv1  gate1433(.a(s_127), .O(gate488inter4));
  nand2 gate1434(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1435(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1436(.a(G1238), .O(gate488inter7));
  inv1  gate1437(.a(G1239), .O(gate488inter8));
  nand2 gate1438(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1439(.a(s_127), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1440(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1441(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1442(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2871(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2872(.a(gate490inter0), .b(s_332), .O(gate490inter1));
  and2  gate2873(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2874(.a(s_332), .O(gate490inter3));
  inv1  gate2875(.a(s_333), .O(gate490inter4));
  nand2 gate2876(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2877(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2878(.a(G1242), .O(gate490inter7));
  inv1  gate2879(.a(G1243), .O(gate490inter8));
  nand2 gate2880(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2881(.a(s_333), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2882(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2883(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2884(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1261(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1262(.a(gate494inter0), .b(s_102), .O(gate494inter1));
  and2  gate1263(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1264(.a(s_102), .O(gate494inter3));
  inv1  gate1265(.a(s_103), .O(gate494inter4));
  nand2 gate1266(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1267(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1268(.a(G1250), .O(gate494inter7));
  inv1  gate1269(.a(G1251), .O(gate494inter8));
  nand2 gate1270(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1271(.a(s_103), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1272(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1273(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1274(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1695(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1696(.a(gate497inter0), .b(s_164), .O(gate497inter1));
  and2  gate1697(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1698(.a(s_164), .O(gate497inter3));
  inv1  gate1699(.a(s_165), .O(gate497inter4));
  nand2 gate1700(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1701(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1702(.a(G1256), .O(gate497inter7));
  inv1  gate1703(.a(G1257), .O(gate497inter8));
  nand2 gate1704(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1705(.a(s_165), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1706(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1707(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1708(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2269(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2270(.a(gate500inter0), .b(s_246), .O(gate500inter1));
  and2  gate2271(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2272(.a(s_246), .O(gate500inter3));
  inv1  gate2273(.a(s_247), .O(gate500inter4));
  nand2 gate2274(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2275(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2276(.a(G1262), .O(gate500inter7));
  inv1  gate2277(.a(G1263), .O(gate500inter8));
  nand2 gate2278(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2279(.a(s_247), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2280(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2281(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2282(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1037(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1038(.a(gate503inter0), .b(s_70), .O(gate503inter1));
  and2  gate1039(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1040(.a(s_70), .O(gate503inter3));
  inv1  gate1041(.a(s_71), .O(gate503inter4));
  nand2 gate1042(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1043(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1044(.a(G1268), .O(gate503inter7));
  inv1  gate1045(.a(G1269), .O(gate503inter8));
  nand2 gate1046(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1047(.a(s_71), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1048(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1049(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1050(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1681(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1682(.a(gate509inter0), .b(s_162), .O(gate509inter1));
  and2  gate1683(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1684(.a(s_162), .O(gate509inter3));
  inv1  gate1685(.a(s_163), .O(gate509inter4));
  nand2 gate1686(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1687(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1688(.a(G1280), .O(gate509inter7));
  inv1  gate1689(.a(G1281), .O(gate509inter8));
  nand2 gate1690(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1691(.a(s_163), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1692(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1693(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1694(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule