module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate767inter0, gate767inter1, gate767inter2, gate767inter3, gate767inter4, gate767inter5, gate767inter6, gate767inter7, gate767inter8, gate767inter9, gate767inter10, gate767inter11, gate767inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate750inter0, gate750inter1, gate750inter2, gate750inter3, gate750inter4, gate750inter5, gate750inter6, gate750inter7, gate750inter8, gate750inter9, gate750inter10, gate750inter11, gate750inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate866inter0, gate866inter1, gate866inter2, gate866inter3, gate866inter4, gate866inter5, gate866inter6, gate866inter7, gate866inter8, gate866inter9, gate866inter10, gate866inter11, gate866inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate797inter0, gate797inter1, gate797inter2, gate797inter3, gate797inter4, gate797inter5, gate797inter6, gate797inter7, gate797inter8, gate797inter9, gate797inter10, gate797inter11, gate797inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate545inter0, gate545inter1, gate545inter2, gate545inter3, gate545inter4, gate545inter5, gate545inter6, gate545inter7, gate545inter8, gate545inter9, gate545inter10, gate545inter11, gate545inter12, gate583inter0, gate583inter1, gate583inter2, gate583inter3, gate583inter4, gate583inter5, gate583inter6, gate583inter7, gate583inter8, gate583inter9, gate583inter10, gate583inter11, gate583inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate814inter0, gate814inter1, gate814inter2, gate814inter3, gate814inter4, gate814inter5, gate814inter6, gate814inter7, gate814inter8, gate814inter9, gate814inter10, gate814inter11, gate814inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate587inter0, gate587inter1, gate587inter2, gate587inter3, gate587inter4, gate587inter5, gate587inter6, gate587inter7, gate587inter8, gate587inter9, gate587inter10, gate587inter11, gate587inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate631inter0, gate631inter1, gate631inter2, gate631inter3, gate631inter4, gate631inter5, gate631inter6, gate631inter7, gate631inter8, gate631inter9, gate631inter10, gate631inter11, gate631inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate758inter0, gate758inter1, gate758inter2, gate758inter3, gate758inter4, gate758inter5, gate758inter6, gate758inter7, gate758inter8, gate758inter9, gate758inter10, gate758inter11, gate758inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate315inter0, gate315inter1, gate315inter2, gate315inter3, gate315inter4, gate315inter5, gate315inter6, gate315inter7, gate315inter8, gate315inter9, gate315inter10, gate315inter11, gate315inter12, gate834inter0, gate834inter1, gate834inter2, gate834inter3, gate834inter4, gate834inter5, gate834inter6, gate834inter7, gate834inter8, gate834inter9, gate834inter10, gate834inter11, gate834inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate303inter0, gate303inter1, gate303inter2, gate303inter3, gate303inter4, gate303inter5, gate303inter6, gate303inter7, gate303inter8, gate303inter9, gate303inter10, gate303inter11, gate303inter12, gate867inter0, gate867inter1, gate867inter2, gate867inter3, gate867inter4, gate867inter5, gate867inter6, gate867inter7, gate867inter8, gate867inter9, gate867inter10, gate867inter11, gate867inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate368inter0, gate368inter1, gate368inter2, gate368inter3, gate368inter4, gate368inter5, gate368inter6, gate368inter7, gate368inter8, gate368inter9, gate368inter10, gate368inter11, gate368inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate643inter0, gate643inter1, gate643inter2, gate643inter3, gate643inter4, gate643inter5, gate643inter6, gate643inter7, gate643inter8, gate643inter9, gate643inter10, gate643inter11, gate643inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate349inter0, gate349inter1, gate349inter2, gate349inter3, gate349inter4, gate349inter5, gate349inter6, gate349inter7, gate349inter8, gate349inter9, gate349inter10, gate349inter11, gate349inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate786inter0, gate786inter1, gate786inter2, gate786inter3, gate786inter4, gate786inter5, gate786inter6, gate786inter7, gate786inter8, gate786inter9, gate786inter10, gate786inter11, gate786inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate370inter0, gate370inter1, gate370inter2, gate370inter3, gate370inter4, gate370inter5, gate370inter6, gate370inter7, gate370inter8, gate370inter9, gate370inter10, gate370inter11, gate370inter12, gate804inter0, gate804inter1, gate804inter2, gate804inter3, gate804inter4, gate804inter5, gate804inter6, gate804inter7, gate804inter8, gate804inter9, gate804inter10, gate804inter11, gate804inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate363inter0, gate363inter1, gate363inter2, gate363inter3, gate363inter4, gate363inter5, gate363inter6, gate363inter7, gate363inter8, gate363inter9, gate363inter10, gate363inter11, gate363inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate552inter0, gate552inter1, gate552inter2, gate552inter3, gate552inter4, gate552inter5, gate552inter6, gate552inter7, gate552inter8, gate552inter9, gate552inter10, gate552inter11, gate552inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate771inter0, gate771inter1, gate771inter2, gate771inter3, gate771inter4, gate771inter5, gate771inter6, gate771inter7, gate771inter8, gate771inter9, gate771inter10, gate771inter11, gate771inter12, gate685inter0, gate685inter1, gate685inter2, gate685inter3, gate685inter4, gate685inter5, gate685inter6, gate685inter7, gate685inter8, gate685inter9, gate685inter10, gate685inter11, gate685inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate680inter0, gate680inter1, gate680inter2, gate680inter3, gate680inter4, gate680inter5, gate680inter6, gate680inter7, gate680inter8, gate680inter9, gate680inter10, gate680inter11, gate680inter12, gate842inter0, gate842inter1, gate842inter2, gate842inter3, gate842inter4, gate842inter5, gate842inter6, gate842inter7, gate842inter8, gate842inter9, gate842inter10, gate842inter11, gate842inter12, gate779inter0, gate779inter1, gate779inter2, gate779inter3, gate779inter4, gate779inter5, gate779inter6, gate779inter7, gate779inter8, gate779inter9, gate779inter10, gate779inter11, gate779inter12, gate542inter0, gate542inter1, gate542inter2, gate542inter3, gate542inter4, gate542inter5, gate542inter6, gate542inter7, gate542inter8, gate542inter9, gate542inter10, gate542inter11, gate542inter12, gate800inter0, gate800inter1, gate800inter2, gate800inter3, gate800inter4, gate800inter5, gate800inter6, gate800inter7, gate800inter8, gate800inter9, gate800inter10, gate800inter11, gate800inter12, gate818inter0, gate818inter1, gate818inter2, gate818inter3, gate818inter4, gate818inter5, gate818inter6, gate818inter7, gate818inter8, gate818inter9, gate818inter10, gate818inter11, gate818inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate642inter0, gate642inter1, gate642inter2, gate642inter3, gate642inter4, gate642inter5, gate642inter6, gate642inter7, gate642inter8, gate642inter9, gate642inter10, gate642inter11, gate642inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate807inter0, gate807inter1, gate807inter2, gate807inter3, gate807inter4, gate807inter5, gate807inter6, gate807inter7, gate807inter8, gate807inter9, gate807inter10, gate807inter11, gate807inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate879inter0, gate879inter1, gate879inter2, gate879inter3, gate879inter4, gate879inter5, gate879inter6, gate879inter7, gate879inter8, gate879inter9, gate879inter10, gate879inter11, gate879inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate855inter0, gate855inter1, gate855inter2, gate855inter3, gate855inter4, gate855inter5, gate855inter6, gate855inter7, gate855inter8, gate855inter9, gate855inter10, gate855inter11, gate855inter12, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12, gate339inter0, gate339inter1, gate339inter2, gate339inter3, gate339inter4, gate339inter5, gate339inter6, gate339inter7, gate339inter8, gate339inter9, gate339inter10, gate339inter11, gate339inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate798inter0, gate798inter1, gate798inter2, gate798inter3, gate798inter4, gate798inter5, gate798inter6, gate798inter7, gate798inter8, gate798inter9, gate798inter10, gate798inter11, gate798inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate765inter0, gate765inter1, gate765inter2, gate765inter3, gate765inter4, gate765inter5, gate765inter6, gate765inter7, gate765inter8, gate765inter9, gate765inter10, gate765inter11, gate765inter12, gate864inter0, gate864inter1, gate864inter2, gate864inter3, gate864inter4, gate864inter5, gate864inter6, gate864inter7, gate864inter8, gate864inter9, gate864inter10, gate864inter11, gate864inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate550inter0, gate550inter1, gate550inter2, gate550inter3, gate550inter4, gate550inter5, gate550inter6, gate550inter7, gate550inter8, gate550inter9, gate550inter10, gate550inter11, gate550inter12;



inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );

  xor2  gate1609(.a(N280), .b(N326), .O(gate97inter0));
  nand2 gate1610(.a(gate97inter0), .b(s_104), .O(gate97inter1));
  and2  gate1611(.a(N280), .b(N326), .O(gate97inter2));
  inv1  gate1612(.a(s_104), .O(gate97inter3));
  inv1  gate1613(.a(s_105), .O(gate97inter4));
  nand2 gate1614(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1615(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1616(.a(N326), .O(gate97inter7));
  inv1  gate1617(.a(N280), .O(gate97inter8));
  nand2 gate1618(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1619(.a(s_105), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1620(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1621(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1622(.a(gate97inter12), .b(gate97inter1), .O(N602));
nand2 gate98( .a(N260), .b(N72), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );

  xor2  gate2057(.a(N612), .b(N49), .O(gate162inter0));
  nand2 gate2058(.a(gate162inter0), .b(s_168), .O(gate162inter1));
  and2  gate2059(.a(N612), .b(N49), .O(gate162inter2));
  inv1  gate2060(.a(s_168), .O(gate162inter3));
  inv1  gate2061(.a(s_169), .O(gate162inter4));
  nand2 gate2062(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2063(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2064(.a(N49), .O(gate162inter7));
  inv1  gate2065(.a(N612), .O(gate162inter8));
  nand2 gate2066(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2067(.a(s_169), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2068(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2069(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2070(.a(gate162inter12), .b(gate162inter1), .O(N907));
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );

  xor2  gate1049(.a(N890), .b(N625), .O(gate235inter0));
  nand2 gate1050(.a(gate235inter0), .b(s_24), .O(gate235inter1));
  and2  gate1051(.a(N890), .b(N625), .O(gate235inter2));
  inv1  gate1052(.a(s_24), .O(gate235inter3));
  inv1  gate1053(.a(s_25), .O(gate235inter4));
  nand2 gate1054(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1055(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1056(.a(N625), .O(gate235inter7));
  inv1  gate1057(.a(N890), .O(gate235inter8));
  nand2 gate1058(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1059(.a(s_25), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1060(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1061(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1062(.a(gate235inter12), .b(gate235inter1), .O(N1063));

  xor2  gate1021(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate1022(.a(gate236inter0), .b(s_20), .O(gate236inter1));
  and2  gate1023(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate1024(.a(s_20), .O(gate236inter3));
  inv1  gate1025(.a(s_21), .O(gate236inter4));
  nand2 gate1026(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1027(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1028(.a(N622), .O(gate236inter7));
  inv1  gate1029(.a(N891), .O(gate236inter8));
  nand2 gate1030(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1031(.a(s_21), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1032(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1033(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1034(.a(gate236inter12), .b(gate236inter1), .O(N1064));
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );

  xor2  gate1511(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate1512(.a(gate245inter0), .b(s_90), .O(gate245inter1));
  and2  gate1513(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate1514(.a(s_90), .O(gate245inter3));
  inv1  gate1515(.a(s_91), .O(gate245inter4));
  nand2 gate1516(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1517(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1518(.a(N745), .O(gate245inter7));
  inv1  gate1519(.a(N1005), .O(gate245inter8));
  nand2 gate1520(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1521(.a(s_91), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1522(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1523(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1524(.a(gate245inter12), .b(gate245inter1), .O(N1130));
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );

  xor2  gate1077(.a(N923), .b(N922), .O(gate269inter0));
  nand2 gate1078(.a(gate269inter0), .b(s_28), .O(gate269inter1));
  and2  gate1079(.a(N923), .b(N922), .O(gate269inter2));
  inv1  gate1080(.a(s_28), .O(gate269inter3));
  inv1  gate1081(.a(s_29), .O(gate269inter4));
  nand2 gate1082(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1083(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1084(.a(N922), .O(gate269inter7));
  inv1  gate1085(.a(N923), .O(gate269inter8));
  nand2 gate1086(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1087(.a(s_29), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1088(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1089(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1090(.a(gate269inter12), .b(gate269inter1), .O(N1188));
inv1 gate270( .a(N1010), .O(N1205) );

  xor2  gate1413(.a(N938), .b(N1010), .O(gate271inter0));
  nand2 gate1414(.a(gate271inter0), .b(s_76), .O(gate271inter1));
  and2  gate1415(.a(N938), .b(N1010), .O(gate271inter2));
  inv1  gate1416(.a(s_76), .O(gate271inter3));
  inv1  gate1417(.a(s_77), .O(gate271inter4));
  nand2 gate1418(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1419(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1420(.a(N1010), .O(gate271inter7));
  inv1  gate1421(.a(N938), .O(gate271inter8));
  nand2 gate1422(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1423(.a(s_77), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1424(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1425(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1426(.a(gate271inter12), .b(gate271inter1), .O(N1206));
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate1133(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate1134(.a(gate277inter0), .b(s_36), .O(gate277inter1));
  and2  gate1135(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate1136(.a(s_36), .O(gate277inter3));
  inv1  gate1137(.a(s_37), .O(gate277inter4));
  nand2 gate1138(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1139(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1140(.a(N1019), .O(gate277inter7));
  inv1  gate1141(.a(N950), .O(gate277inter8));
  nand2 gate1142(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1143(.a(s_37), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1144(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1145(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1146(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );

  xor2  gate1553(.a(N984), .b(N981), .O(gate296inter0));
  nand2 gate1554(.a(gate296inter0), .b(s_96), .O(gate296inter1));
  and2  gate1555(.a(N984), .b(N981), .O(gate296inter2));
  inv1  gate1556(.a(s_96), .O(gate296inter3));
  inv1  gate1557(.a(s_97), .O(gate296inter4));
  nand2 gate1558(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1559(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1560(.a(N981), .O(gate296inter7));
  inv1  gate1561(.a(N984), .O(gate296inter8));
  nand2 gate1562(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1563(.a(s_97), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1564(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1565(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1566(.a(gate296inter12), .b(gate296inter1), .O(N1231));
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );

  xor2  gate1301(.a(N1001), .b(N1049), .O(gate303inter0));
  nand2 gate1302(.a(gate303inter0), .b(s_60), .O(gate303inter1));
  and2  gate1303(.a(N1001), .b(N1049), .O(gate303inter2));
  inv1  gate1304(.a(s_60), .O(gate303inter3));
  inv1  gate1305(.a(s_61), .O(gate303inter4));
  nand2 gate1306(.a(gate303inter4), .b(gate303inter3), .O(gate303inter5));
  nor2  gate1307(.a(gate303inter5), .b(gate303inter2), .O(gate303inter6));
  inv1  gate1308(.a(N1049), .O(gate303inter7));
  inv1  gate1309(.a(N1001), .O(gate303inter8));
  nand2 gate1310(.a(gate303inter8), .b(gate303inter7), .O(gate303inter9));
  nand2 gate1311(.a(s_61), .b(gate303inter3), .O(gate303inter10));
  nor2  gate1312(.a(gate303inter10), .b(gate303inter9), .O(gate303inter11));
  nor2  gate1313(.a(gate303inter11), .b(gate303inter6), .O(gate303inter12));
  nand2 gate1314(.a(gate303inter12), .b(gate303inter1), .O(N1242));
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate1847(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate1848(.a(gate312inter0), .b(s_138), .O(gate312inter1));
  and2  gate1849(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate1850(.a(s_138), .O(gate312inter3));
  inv1  gate1851(.a(s_139), .O(gate312inter4));
  nand2 gate1852(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate1853(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate1854(.a(N631), .O(gate312inter7));
  inv1  gate1855(.a(N1159), .O(gate312inter8));
  nand2 gate1856(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate1857(.a(s_139), .b(gate312inter3), .O(gate312inter10));
  nor2  gate1858(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate1859(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate1860(.a(gate312inter12), .b(gate312inter1), .O(N1267));

  xor2  gate951(.a(N1205), .b(N688), .O(gate313inter0));
  nand2 gate952(.a(gate313inter0), .b(s_10), .O(gate313inter1));
  and2  gate953(.a(N1205), .b(N688), .O(gate313inter2));
  inv1  gate954(.a(s_10), .O(gate313inter3));
  inv1  gate955(.a(s_11), .O(gate313inter4));
  nand2 gate956(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate957(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate958(.a(N688), .O(gate313inter7));
  inv1  gate959(.a(N1205), .O(gate313inter8));
  nand2 gate960(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate961(.a(s_11), .b(gate313inter3), .O(gate313inter10));
  nor2  gate962(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate963(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate964(.a(gate313inter12), .b(gate313inter1), .O(N1309));
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );

  xor2  gate1231(.a(N1209), .b(N694), .O(gate315inter0));
  nand2 gate1232(.a(gate315inter0), .b(s_50), .O(gate315inter1));
  and2  gate1233(.a(N1209), .b(N694), .O(gate315inter2));
  inv1  gate1234(.a(s_50), .O(gate315inter3));
  inv1  gate1235(.a(s_51), .O(gate315inter4));
  nand2 gate1236(.a(gate315inter4), .b(gate315inter3), .O(gate315inter5));
  nor2  gate1237(.a(gate315inter5), .b(gate315inter2), .O(gate315inter6));
  inv1  gate1238(.a(N694), .O(gate315inter7));
  inv1  gate1239(.a(N1209), .O(gate315inter8));
  nand2 gate1240(.a(gate315inter8), .b(gate315inter7), .O(gate315inter9));
  nand2 gate1241(.a(s_51), .b(gate315inter3), .O(gate315inter10));
  nor2  gate1242(.a(gate315inter10), .b(gate315inter9), .O(gate315inter11));
  nor2  gate1243(.a(gate315inter11), .b(gate315inter6), .O(gate315inter12));
  nand2 gate1244(.a(gate315inter12), .b(gate315inter1), .O(N1311));

  xor2  gate1329(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate1330(.a(gate316inter0), .b(s_64), .O(gate316inter1));
  and2  gate1331(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate1332(.a(s_64), .O(gate316inter3));
  inv1  gate1333(.a(s_65), .O(gate316inter4));
  nand2 gate1334(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate1335(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate1336(.a(N697), .O(gate316inter7));
  inv1  gate1337(.a(N1211), .O(gate316inter8));
  nand2 gate1338(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate1339(.a(s_65), .b(gate316inter3), .O(gate316inter10));
  nor2  gate1340(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate1341(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate1342(.a(gate316inter12), .b(gate316inter1), .O(N1312));
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );

  xor2  gate1567(.a(N1160), .b(N1267), .O(gate328inter0));
  nand2 gate1568(.a(gate328inter0), .b(s_98), .O(gate328inter1));
  and2  gate1569(.a(N1160), .b(N1267), .O(gate328inter2));
  inv1  gate1570(.a(s_98), .O(gate328inter3));
  inv1  gate1571(.a(s_99), .O(gate328inter4));
  nand2 gate1572(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate1573(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate1574(.a(N1267), .O(gate328inter7));
  inv1  gate1575(.a(N1160), .O(gate328inter8));
  nand2 gate1576(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate1577(.a(s_99), .b(gate328inter3), .O(gate328inter10));
  nor2  gate1578(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate1579(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate1580(.a(gate328inter12), .b(gate328inter1), .O(N1344));
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );

  xor2  gate1959(.a(N1214), .b(N1313), .O(gate339inter0));
  nand2 gate1960(.a(gate339inter0), .b(s_154), .O(gate339inter1));
  and2  gate1961(.a(N1214), .b(N1313), .O(gate339inter2));
  inv1  gate1962(.a(s_154), .O(gate339inter3));
  inv1  gate1963(.a(s_155), .O(gate339inter4));
  nand2 gate1964(.a(gate339inter4), .b(gate339inter3), .O(gate339inter5));
  nor2  gate1965(.a(gate339inter5), .b(gate339inter2), .O(gate339inter6));
  inv1  gate1966(.a(N1313), .O(gate339inter7));
  inv1  gate1967(.a(N1214), .O(gate339inter8));
  nand2 gate1968(.a(gate339inter8), .b(gate339inter7), .O(gate339inter9));
  nand2 gate1969(.a(s_155), .b(gate339inter3), .O(gate339inter10));
  nor2  gate1970(.a(gate339inter10), .b(gate339inter9), .O(gate339inter11));
  nor2  gate1971(.a(gate339inter11), .b(gate339inter6), .O(gate339inter12));
  nand2 gate1972(.a(gate339inter12), .b(gate339inter1), .O(N1364));
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );

  xor2  gate1259(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate1260(.a(gate342inter0), .b(s_54), .O(gate342inter1));
  and2  gate1261(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate1262(.a(s_54), .O(gate342inter3));
  inv1  gate1263(.a(s_55), .O(gate342inter4));
  nand2 gate1264(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate1265(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate1266(.a(N1316), .O(gate342inter7));
  inv1  gate1267(.a(N1224), .O(gate342inter8));
  nand2 gate1268(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate1269(.a(s_55), .b(gate342inter3), .O(gate342inter10));
  nor2  gate1270(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate1271(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate1272(.a(gate342inter12), .b(gate342inter1), .O(N1373));
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );

  xor2  gate1399(.a(N993), .b(N1235), .O(gate349inter0));
  nand2 gate1400(.a(gate349inter0), .b(s_74), .O(gate349inter1));
  and2  gate1401(.a(N993), .b(N1235), .O(gate349inter2));
  inv1  gate1402(.a(s_74), .O(gate349inter3));
  inv1  gate1403(.a(s_75), .O(gate349inter4));
  nand2 gate1404(.a(gate349inter4), .b(gate349inter3), .O(gate349inter5));
  nor2  gate1405(.a(gate349inter5), .b(gate349inter2), .O(gate349inter6));
  inv1  gate1406(.a(N1235), .O(gate349inter7));
  inv1  gate1407(.a(N993), .O(gate349inter8));
  nand2 gate1408(.a(gate349inter8), .b(gate349inter7), .O(gate349inter9));
  nand2 gate1409(.a(s_75), .b(gate349inter3), .O(gate349inter10));
  nor2  gate1410(.a(gate349inter10), .b(gate349inter9), .O(gate349inter11));
  nor2  gate1411(.a(gate349inter11), .b(gate349inter6), .O(gate349inter12));
  nand2 gate1412(.a(gate349inter12), .b(gate349inter1), .O(N1389));
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );

  xor2  gate1973(.a(N1388), .b(N637), .O(gate362inter0));
  nand2 gate1974(.a(gate362inter0), .b(s_156), .O(gate362inter1));
  and2  gate1975(.a(N1388), .b(N637), .O(gate362inter2));
  inv1  gate1976(.a(s_156), .O(gate362inter3));
  inv1  gate1977(.a(s_157), .O(gate362inter4));
  nand2 gate1978(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate1979(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate1980(.a(N637), .O(gate362inter7));
  inv1  gate1981(.a(N1388), .O(gate362inter8));
  nand2 gate1982(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate1983(.a(s_157), .b(gate362inter3), .O(gate362inter10));
  nor2  gate1984(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate1985(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate1986(.a(gate362inter12), .b(gate362inter1), .O(N1434));

  xor2  gate1595(.a(N1396), .b(N640), .O(gate363inter0));
  nand2 gate1596(.a(gate363inter0), .b(s_102), .O(gate363inter1));
  and2  gate1597(.a(N1396), .b(N640), .O(gate363inter2));
  inv1  gate1598(.a(s_102), .O(gate363inter3));
  inv1  gate1599(.a(s_103), .O(gate363inter4));
  nand2 gate1600(.a(gate363inter4), .b(gate363inter3), .O(gate363inter5));
  nor2  gate1601(.a(gate363inter5), .b(gate363inter2), .O(gate363inter6));
  inv1  gate1602(.a(N640), .O(gate363inter7));
  inv1  gate1603(.a(N1396), .O(gate363inter8));
  nand2 gate1604(.a(gate363inter8), .b(gate363inter7), .O(gate363inter9));
  nand2 gate1605(.a(s_103), .b(gate363inter3), .O(gate363inter10));
  nor2  gate1606(.a(gate363inter10), .b(gate363inter9), .O(gate363inter11));
  nor2  gate1607(.a(gate363inter11), .b(gate363inter6), .O(gate363inter12));
  nand2 gate1608(.a(gate363inter12), .b(gate363inter1), .O(N1438));

  xor2  gate1791(.a(N1398), .b(N646), .O(gate364inter0));
  nand2 gate1792(.a(gate364inter0), .b(s_130), .O(gate364inter1));
  and2  gate1793(.a(N1398), .b(N646), .O(gate364inter2));
  inv1  gate1794(.a(s_130), .O(gate364inter3));
  inv1  gate1795(.a(s_131), .O(gate364inter4));
  nand2 gate1796(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate1797(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate1798(.a(N646), .O(gate364inter7));
  inv1  gate1799(.a(N1398), .O(gate364inter8));
  nand2 gate1800(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate1801(.a(s_131), .b(gate364inter3), .O(gate364inter10));
  nor2  gate1802(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate1803(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate1804(.a(gate364inter12), .b(gate364inter1), .O(N1439));
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );

  xor2  gate1343(.a(N1149), .b(N1352), .O(gate368inter0));
  nand2 gate1344(.a(gate368inter0), .b(s_66), .O(gate368inter1));
  and2  gate1345(.a(N1149), .b(N1352), .O(gate368inter2));
  inv1  gate1346(.a(s_66), .O(gate368inter3));
  inv1  gate1347(.a(s_67), .O(gate368inter4));
  nand2 gate1348(.a(gate368inter4), .b(gate368inter3), .O(gate368inter5));
  nor2  gate1349(.a(gate368inter5), .b(gate368inter2), .O(gate368inter6));
  inv1  gate1350(.a(N1352), .O(gate368inter7));
  inv1  gate1351(.a(N1149), .O(gate368inter8));
  nand2 gate1352(.a(gate368inter8), .b(gate368inter7), .O(gate368inter9));
  nand2 gate1353(.a(s_67), .b(gate368inter3), .O(gate368inter10));
  nor2  gate1354(.a(gate368inter10), .b(gate368inter9), .O(gate368inter11));
  nor2  gate1355(.a(gate368inter11), .b(gate368inter6), .O(gate368inter12));
  nand2 gate1356(.a(gate368inter12), .b(gate368inter1), .O(N1445));
inv1 gate369( .a(N1352), .O(N1446) );

  xor2  gate1525(.a(N1151), .b(N1358), .O(gate370inter0));
  nand2 gate1526(.a(gate370inter0), .b(s_92), .O(gate370inter1));
  and2  gate1527(.a(N1151), .b(N1358), .O(gate370inter2));
  inv1  gate1528(.a(s_92), .O(gate370inter3));
  inv1  gate1529(.a(s_93), .O(gate370inter4));
  nand2 gate1530(.a(gate370inter4), .b(gate370inter3), .O(gate370inter5));
  nor2  gate1531(.a(gate370inter5), .b(gate370inter2), .O(gate370inter6));
  inv1  gate1532(.a(N1358), .O(gate370inter7));
  inv1  gate1533(.a(N1151), .O(gate370inter8));
  nand2 gate1534(.a(gate370inter8), .b(gate370inter7), .O(gate370inter9));
  nand2 gate1535(.a(s_93), .b(gate370inter3), .O(gate370inter10));
  nor2  gate1536(.a(gate370inter10), .b(gate370inter9), .O(gate370inter11));
  nor2  gate1537(.a(gate370inter11), .b(gate370inter6), .O(gate370inter12));
  nand2 gate1538(.a(gate370inter12), .b(gate370inter1), .O(N1447));
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );

  xor2  gate1385(.a(N1240), .b(N1390), .O(gate392inter0));
  nand2 gate1386(.a(gate392inter0), .b(s_72), .O(gate392inter1));
  and2  gate1387(.a(N1240), .b(N1390), .O(gate392inter2));
  inv1  gate1388(.a(s_72), .O(gate392inter3));
  inv1  gate1389(.a(s_73), .O(gate392inter4));
  nand2 gate1390(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1391(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1392(.a(N1390), .O(gate392inter7));
  inv1  gate1393(.a(N1240), .O(gate392inter8));
  nand2 gate1394(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1395(.a(s_73), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1396(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1397(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1398(.a(gate392inter12), .b(gate392inter1), .O(N1476));
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );

  xor2  gate1637(.a(N1493), .b(N1453), .O(gate416inter0));
  nand2 gate1638(.a(gate416inter0), .b(s_108), .O(gate416inter1));
  and2  gate1639(.a(N1493), .b(N1453), .O(gate416inter2));
  inv1  gate1640(.a(s_108), .O(gate416inter3));
  inv1  gate1641(.a(s_109), .O(gate416inter4));
  nand2 gate1642(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1643(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1644(.a(N1453), .O(gate416inter7));
  inv1  gate1645(.a(N1493), .O(gate416inter8));
  nand2 gate1646(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1647(.a(s_109), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1648(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1649(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1650(.a(gate416inter12), .b(gate416inter1), .O(N1521));
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );

  xor2  gate1105(.a(N1500), .b(N1469), .O(gate426inter0));
  nand2 gate1106(.a(gate426inter0), .b(s_32), .O(gate426inter1));
  and2  gate1107(.a(N1500), .b(N1469), .O(gate426inter2));
  inv1  gate1108(.a(s_32), .O(gate426inter3));
  inv1  gate1109(.a(s_33), .O(gate426inter4));
  nand2 gate1110(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1111(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1112(.a(N1469), .O(gate426inter7));
  inv1  gate1113(.a(N1500), .O(gate426inter8));
  nand2 gate1114(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1115(.a(s_33), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1116(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1117(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1118(.a(gate426inter12), .b(gate426inter1), .O(N1537));
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );

  xor2  gate2015(.a(N1531), .b(N1484), .O(gate432inter0));
  nand2 gate2016(.a(gate432inter0), .b(s_162), .O(gate432inter1));
  and2  gate2017(.a(N1531), .b(N1484), .O(gate432inter2));
  inv1  gate2018(.a(s_162), .O(gate432inter3));
  inv1  gate2019(.a(s_163), .O(gate432inter4));
  nand2 gate2020(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2021(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2022(.a(N1484), .O(gate432inter7));
  inv1  gate2023(.a(N1531), .O(gate432inter8));
  nand2 gate2024(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2025(.a(s_163), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2026(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2027(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2028(.a(gate432inter12), .b(gate432inter1), .O(N1567));
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );

  xor2  gate1175(.a(N1530), .b(N1540), .O(gate440inter0));
  nand2 gate1176(.a(gate440inter0), .b(s_42), .O(gate440inter1));
  and2  gate1177(.a(N1530), .b(N1540), .O(gate440inter2));
  inv1  gate1178(.a(s_42), .O(gate440inter3));
  inv1  gate1179(.a(s_43), .O(gate440inter4));
  nand2 gate1180(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1181(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1182(.a(N1540), .O(gate440inter7));
  inv1  gate1183(.a(N1530), .O(gate440inter8));
  nand2 gate1184(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1185(.a(s_43), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1186(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1187(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1188(.a(gate440inter12), .b(gate440inter1), .O(N1594));
inv1 gate441( .a(N1540), .O(N1595) );

  xor2  gate1287(.a(N1568), .b(N1567), .O(gate442inter0));
  nand2 gate1288(.a(gate442inter0), .b(s_58), .O(gate442inter1));
  and2  gate1289(.a(N1568), .b(N1567), .O(gate442inter2));
  inv1  gate1290(.a(s_58), .O(gate442inter3));
  inv1  gate1291(.a(s_59), .O(gate442inter4));
  nand2 gate1292(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1293(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1294(.a(N1567), .O(gate442inter7));
  inv1  gate1295(.a(N1568), .O(gate442inter8));
  nand2 gate1296(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1297(.a(s_59), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1298(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1299(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1300(.a(gate442inter12), .b(gate442inter1), .O(N1596));
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );

  xor2  gate1483(.a(N1595), .b(N1478), .O(gate452inter0));
  nand2 gate1484(.a(gate452inter0), .b(s_86), .O(gate452inter1));
  and2  gate1485(.a(N1595), .b(N1478), .O(gate452inter2));
  inv1  gate1486(.a(s_86), .O(gate452inter3));
  inv1  gate1487(.a(s_87), .O(gate452inter4));
  nand2 gate1488(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1489(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1490(.a(N1478), .O(gate452inter7));
  inv1  gate1491(.a(N1595), .O(gate452inter8));
  nand2 gate1492(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1493(.a(s_87), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1494(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1495(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1496(.a(gate452inter12), .b(gate452inter1), .O(N1636));
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );

  xor2  gate1441(.a(N893), .b(N1596), .O(gate462inter0));
  nand2 gate1442(.a(gate462inter0), .b(s_80), .O(gate462inter1));
  and2  gate1443(.a(N893), .b(N1596), .O(gate462inter2));
  inv1  gate1444(.a(s_80), .O(gate462inter3));
  inv1  gate1445(.a(s_81), .O(gate462inter4));
  nand2 gate1446(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1447(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1448(.a(N1596), .O(gate462inter7));
  inv1  gate1449(.a(N893), .O(gate462inter8));
  nand2 gate1450(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1451(.a(s_81), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1452(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1453(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1454(.a(gate462inter12), .b(gate462inter1), .O(N1671));
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );

  xor2  gate2001(.a(N1681), .b(N1031), .O(gate483inter0));
  nand2 gate2002(.a(gate483inter0), .b(s_160), .O(gate483inter1));
  and2  gate2003(.a(N1681), .b(N1031), .O(gate483inter2));
  inv1  gate2004(.a(s_160), .O(gate483inter3));
  inv1  gate2005(.a(s_161), .O(gate483inter4));
  nand2 gate2006(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2007(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2008(.a(N1031), .O(gate483inter7));
  inv1  gate2009(.a(N1681), .O(gate483inter8));
  nand2 gate2010(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2011(.a(s_161), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2012(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2013(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2014(.a(gate483inter12), .b(gate483inter1), .O(N1713));
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );

  xor2  gate1819(.a(N1709), .b(N1600), .O(gate497inter0));
  nand2 gate1820(.a(gate497inter0), .b(s_134), .O(gate497inter1));
  and2  gate1821(.a(N1709), .b(N1600), .O(gate497inter2));
  inv1  gate1822(.a(s_134), .O(gate497inter3));
  inv1  gate1823(.a(s_135), .O(gate497inter4));
  nand2 gate1824(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1825(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1826(.a(N1600), .O(gate497inter7));
  inv1  gate1827(.a(N1709), .O(gate497inter8));
  nand2 gate1828(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1829(.a(s_135), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1830(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1831(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1832(.a(gate497inter12), .b(gate497inter1), .O(N1746));
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );

  xor2  gate1777(.a(N1721), .b(N1537), .O(gate501inter0));
  nand2 gate1778(.a(gate501inter0), .b(s_128), .O(gate501inter1));
  and2  gate1779(.a(N1721), .b(N1537), .O(gate501inter2));
  inv1  gate1780(.a(s_128), .O(gate501inter3));
  inv1  gate1781(.a(s_129), .O(gate501inter4));
  nand2 gate1782(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1783(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1784(.a(N1537), .O(gate501inter7));
  inv1  gate1785(.a(N1721), .O(gate501inter8));
  nand2 gate1786(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1787(.a(s_129), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1788(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1789(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1790(.a(gate501inter12), .b(gate501inter1), .O(N1759));
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );

  xor2  gate1147(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate1148(.a(gate508inter0), .b(s_38), .O(gate508inter1));
  and2  gate1149(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate1150(.a(s_38), .O(gate508inter3));
  inv1  gate1151(.a(s_39), .O(gate508inter4));
  nand2 gate1152(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1153(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1154(.a(N1723), .O(gate508inter7));
  inv1  gate1155(.a(N1413), .O(gate508inter8));
  nand2 gate1156(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1157(.a(s_39), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1158(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1159(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1160(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate923(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate924(.a(gate513inter0), .b(s_6), .O(gate513inter1));
  and2  gate925(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate926(.a(s_6), .O(gate513inter3));
  inv1  gate927(.a(s_7), .O(gate513inter4));
  nand2 gate928(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate929(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate930(.a(N1731), .O(gate513inter7));
  inv1  gate931(.a(N1682), .O(gate513inter8));
  nand2 gate932(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate933(.a(s_7), .b(gate513inter3), .O(gate513inter10));
  nor2  gate934(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate935(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate936(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );

  xor2  gate1035(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate1036(.a(gate520inter0), .b(s_22), .O(gate520inter1));
  and2  gate1037(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate1038(.a(s_22), .O(gate520inter3));
  inv1  gate1039(.a(s_23), .O(gate520inter4));
  nand2 gate1040(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate1041(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate1042(.a(N1751), .O(gate520inter7));
  inv1  gate1043(.a(N1155), .O(gate520inter8));
  nand2 gate1044(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate1045(.a(s_23), .b(gate520inter3), .O(gate520inter10));
  nor2  gate1046(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate1047(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate1048(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate1063(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate1064(.a(gate522inter0), .b(s_26), .O(gate522inter1));
  and2  gate1065(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate1066(.a(s_26), .O(gate522inter3));
  inv1  gate1067(.a(s_27), .O(gate522inter4));
  nand2 gate1068(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate1069(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate1070(.a(N1740), .O(gate522inter7));
  inv1  gate1071(.a(N1769), .O(gate522inter8));
  nand2 gate1072(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate1073(.a(s_27), .b(gate522inter3), .O(gate522inter10));
  nor2  gate1074(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate1075(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate1076(.a(gate522inter12), .b(gate522inter1), .O(N1798));
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );

  xor2  gate1735(.a(N1787), .b(N1810), .O(gate542inter0));
  nand2 gate1736(.a(gate542inter0), .b(s_122), .O(gate542inter1));
  and2  gate1737(.a(N1787), .b(N1810), .O(gate542inter2));
  inv1  gate1738(.a(s_122), .O(gate542inter3));
  inv1  gate1739(.a(s_123), .O(gate542inter4));
  nand2 gate1740(.a(gate542inter4), .b(gate542inter3), .O(gate542inter5));
  nor2  gate1741(.a(gate542inter5), .b(gate542inter2), .O(gate542inter6));
  inv1  gate1742(.a(N1810), .O(gate542inter7));
  inv1  gate1743(.a(N1787), .O(gate542inter8));
  nand2 gate1744(.a(gate542inter8), .b(gate542inter7), .O(gate542inter9));
  nand2 gate1745(.a(s_123), .b(gate542inter3), .O(gate542inter10));
  nor2  gate1746(.a(gate542inter10), .b(gate542inter9), .O(gate542inter11));
  nor2  gate1747(.a(gate542inter11), .b(gate542inter6), .O(gate542inter12));
  nand2 gate1748(.a(gate542inter12), .b(gate542inter1), .O(N1841));
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );

  xor2  gate993(.a(N1825), .b(N1795), .O(gate545inter0));
  nand2 gate994(.a(gate545inter0), .b(s_16), .O(gate545inter1));
  and2  gate995(.a(N1825), .b(N1795), .O(gate545inter2));
  inv1  gate996(.a(s_16), .O(gate545inter3));
  inv1  gate997(.a(s_17), .O(gate545inter4));
  nand2 gate998(.a(gate545inter4), .b(gate545inter3), .O(gate545inter5));
  nor2  gate999(.a(gate545inter5), .b(gate545inter2), .O(gate545inter6));
  inv1  gate1000(.a(N1795), .O(gate545inter7));
  inv1  gate1001(.a(N1825), .O(gate545inter8));
  nand2 gate1002(.a(gate545inter8), .b(gate545inter7), .O(gate545inter9));
  nand2 gate1003(.a(s_17), .b(gate545inter3), .O(gate545inter10));
  nor2  gate1004(.a(gate545inter10), .b(gate545inter9), .O(gate545inter11));
  nor2  gate1005(.a(gate545inter11), .b(gate545inter6), .O(gate545inter12));
  nand2 gate1006(.a(gate545inter12), .b(gate545inter1), .O(N1850));

  xor2  gate1469(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate1470(.a(gate546inter0), .b(s_84), .O(gate546inter1));
  and2  gate1471(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate1472(.a(s_84), .O(gate546inter3));
  inv1  gate1473(.a(s_85), .O(gate546inter4));
  nand2 gate1474(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate1475(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate1476(.a(N1319), .O(gate546inter7));
  inv1  gate1477(.a(N1827), .O(gate546inter8));
  nand2 gate1478(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate1479(.a(s_85), .b(gate546inter3), .O(gate546inter10));
  nor2  gate1480(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate1481(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate1482(.a(gate546inter12), .b(gate546inter1), .O(N1852));

  xor2  gate1805(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate1806(.a(gate547inter0), .b(s_132), .O(gate547inter1));
  and2  gate1807(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate1808(.a(s_132), .O(gate547inter3));
  inv1  gate1809(.a(s_133), .O(gate547inter4));
  nand2 gate1810(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate1811(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate1812(.a(N1815), .O(gate547inter7));
  inv1  gate1813(.a(N1707), .O(gate547inter8));
  nand2 gate1814(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate1815(.a(s_133), .b(gate547inter3), .O(gate547inter10));
  nor2  gate1816(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate1817(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate1818(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );

  xor2  gate2071(.a(N290), .b(N1798), .O(gate550inter0));
  nand2 gate2072(.a(gate550inter0), .b(s_170), .O(gate550inter1));
  and2  gate2073(.a(N290), .b(N1798), .O(gate550inter2));
  inv1  gate2074(.a(s_170), .O(gate550inter3));
  inv1  gate2075(.a(s_171), .O(gate550inter4));
  nand2 gate2076(.a(gate550inter4), .b(gate550inter3), .O(gate550inter5));
  nor2  gate2077(.a(gate550inter5), .b(gate550inter2), .O(gate550inter6));
  inv1  gate2078(.a(N1798), .O(gate550inter7));
  inv1  gate2079(.a(N290), .O(gate550inter8));
  nand2 gate2080(.a(gate550inter8), .b(gate550inter7), .O(gate550inter9));
  nand2 gate2081(.a(s_171), .b(gate550inter3), .O(gate550inter10));
  nor2  gate2082(.a(gate550inter10), .b(gate550inter9), .O(gate550inter11));
  nor2  gate2083(.a(gate550inter11), .b(gate550inter6), .O(gate550inter12));
  nand2 gate2084(.a(gate550inter12), .b(gate550inter1), .O(N1858));
inv1 gate551( .a(N1812), .O(N1864) );

  xor2  gate1623(.a(N1728), .b(N1812), .O(gate552inter0));
  nand2 gate1624(.a(gate552inter0), .b(s_106), .O(gate552inter1));
  and2  gate1625(.a(N1728), .b(N1812), .O(gate552inter2));
  inv1  gate1626(.a(s_106), .O(gate552inter3));
  inv1  gate1627(.a(s_107), .O(gate552inter4));
  nand2 gate1628(.a(gate552inter4), .b(gate552inter3), .O(gate552inter5));
  nor2  gate1629(.a(gate552inter5), .b(gate552inter2), .O(gate552inter6));
  inv1  gate1630(.a(N1812), .O(gate552inter7));
  inv1  gate1631(.a(N1728), .O(gate552inter8));
  nand2 gate1632(.a(gate552inter8), .b(gate552inter7), .O(gate552inter9));
  nand2 gate1633(.a(s_107), .b(gate552inter3), .O(gate552inter10));
  nor2  gate1634(.a(gate552inter10), .b(gate552inter9), .O(gate552inter11));
  nor2  gate1635(.a(gate552inter11), .b(gate552inter6), .O(gate552inter12));
  nand2 gate1636(.a(gate552inter12), .b(gate552inter1), .O(N1865));
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate1875(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate1876(.a(gate574inter0), .b(s_142), .O(gate574inter1));
  and2  gate1877(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate1878(.a(s_142), .O(gate574inter3));
  inv1  gate1879(.a(s_143), .O(gate574inter4));
  nand2 gate1880(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate1881(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate1882(.a(N1872), .O(gate574inter7));
  inv1  gate1883(.a(N919), .O(gate574inter8));
  nand2 gate1884(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate1885(.a(s_143), .b(gate574inter3), .O(gate574inter10));
  nor2  gate1886(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate1887(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate1888(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );

  xor2  gate1007(.a(N1911), .b(N1882), .O(gate583inter0));
  nand2 gate1008(.a(gate583inter0), .b(s_18), .O(gate583inter1));
  and2  gate1009(.a(N1911), .b(N1882), .O(gate583inter2));
  inv1  gate1010(.a(s_18), .O(gate583inter3));
  inv1  gate1011(.a(s_19), .O(gate583inter4));
  nand2 gate1012(.a(gate583inter4), .b(gate583inter3), .O(gate583inter5));
  nor2  gate1013(.a(gate583inter5), .b(gate583inter2), .O(gate583inter6));
  inv1  gate1014(.a(N1882), .O(gate583inter7));
  inv1  gate1015(.a(N1911), .O(gate583inter8));
  nand2 gate1016(.a(gate583inter8), .b(gate583inter7), .O(gate583inter9));
  nand2 gate1017(.a(s_19), .b(gate583inter3), .O(gate583inter10));
  nor2  gate1018(.a(gate583inter10), .b(gate583inter9), .O(gate583inter11));
  nor2  gate1019(.a(gate583inter11), .b(gate583inter6), .O(gate583inter12));
  nand2 gate1020(.a(gate583inter12), .b(gate583inter1), .O(N1936));
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );

  xor2  gate1119(.a(N1922), .b(N676), .O(gate587inter0));
  nand2 gate1120(.a(gate587inter0), .b(s_34), .O(gate587inter1));
  and2  gate1121(.a(N1922), .b(N676), .O(gate587inter2));
  inv1  gate1122(.a(s_34), .O(gate587inter3));
  inv1  gate1123(.a(s_35), .O(gate587inter4));
  nand2 gate1124(.a(gate587inter4), .b(gate587inter3), .O(gate587inter5));
  nor2  gate1125(.a(gate587inter5), .b(gate587inter2), .O(gate587inter6));
  inv1  gate1126(.a(N676), .O(gate587inter7));
  inv1  gate1127(.a(N1922), .O(gate587inter8));
  nand2 gate1128(.a(gate587inter8), .b(gate587inter7), .O(gate587inter9));
  nand2 gate1129(.a(s_35), .b(gate587inter3), .O(gate587inter10));
  nor2  gate1130(.a(gate587inter10), .b(gate587inter9), .O(gate587inter11));
  nor2  gate1131(.a(gate587inter11), .b(gate587inter6), .O(gate587inter12));
  nand2 gate1132(.a(gate587inter12), .b(gate587inter1), .O(N1942));
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );

  xor2  gate1581(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate1582(.a(gate601inter0), .b(s_100), .O(gate601inter1));
  and2  gate1583(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate1584(.a(s_100), .O(gate601inter3));
  inv1  gate1585(.a(s_101), .O(gate601inter4));
  nand2 gate1586(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate1587(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate1588(.a(N1921), .O(gate601inter7));
  inv1  gate1589(.a(N1942), .O(gate601inter8));
  nand2 gate1590(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate1591(.a(s_101), .b(gate601inter3), .O(gate601inter10));
  nor2  gate1592(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate1593(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate1594(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate1455(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate1456(.a(gate612inter0), .b(s_82), .O(gate612inter1));
  and2  gate1457(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate1458(.a(s_82), .O(gate612inter3));
  inv1  gate1459(.a(s_83), .O(gate612inter4));
  nand2 gate1460(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate1461(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate1462(.a(N673), .O(gate612inter7));
  inv1  gate1463(.a(N1976), .O(gate612inter8));
  nand2 gate1464(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate1465(.a(s_83), .b(gate612inter3), .O(gate612inter10));
  nor2  gate1466(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate1467(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate1468(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );

  xor2  gate1161(.a(N2013), .b(N1875), .O(gate631inter0));
  nand2 gate1162(.a(gate631inter0), .b(s_40), .O(gate631inter1));
  and2  gate1163(.a(N2013), .b(N1875), .O(gate631inter2));
  inv1  gate1164(.a(s_40), .O(gate631inter3));
  inv1  gate1165(.a(s_41), .O(gate631inter4));
  nand2 gate1166(.a(gate631inter4), .b(gate631inter3), .O(gate631inter5));
  nor2  gate1167(.a(gate631inter5), .b(gate631inter2), .O(gate631inter6));
  inv1  gate1168(.a(N1875), .O(gate631inter7));
  inv1  gate1169(.a(N2013), .O(gate631inter8));
  nand2 gate1170(.a(gate631inter8), .b(gate631inter7), .O(gate631inter9));
  nand2 gate1171(.a(s_41), .b(gate631inter3), .O(gate631inter10));
  nor2  gate1172(.a(gate631inter10), .b(gate631inter9), .O(gate631inter11));
  nor2  gate1173(.a(gate631inter11), .b(gate631inter6), .O(gate631inter12));
  nand2 gate1174(.a(gate631inter12), .b(gate631inter1), .O(N2036));
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );

  xor2  gate1217(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate1218(.a(gate634inter0), .b(s_48), .O(gate634inter1));
  and2  gate1219(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate1220(.a(s_48), .O(gate634inter3));
  inv1  gate1221(.a(s_49), .O(gate634inter4));
  nand2 gate1222(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate1223(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate1224(.a(N1534), .O(gate634inter7));
  inv1  gate1225(.a(N2021), .O(gate634inter8));
  nand2 gate1226(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate1227(.a(s_49), .b(gate634inter3), .O(gate634inter10));
  nor2  gate1228(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate1229(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate1230(.a(gate634inter12), .b(gate634inter1), .O(N2039));

  xor2  gate1931(.a(N2003), .b(N2023), .O(gate635inter0));
  nand2 gate1932(.a(gate635inter0), .b(s_150), .O(gate635inter1));
  and2  gate1933(.a(N2003), .b(N2023), .O(gate635inter2));
  inv1  gate1934(.a(s_150), .O(gate635inter3));
  inv1  gate1935(.a(s_151), .O(gate635inter4));
  nand2 gate1936(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate1937(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate1938(.a(N2023), .O(gate635inter7));
  inv1  gate1939(.a(N2003), .O(gate635inter8));
  nand2 gate1940(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate1941(.a(s_151), .b(gate635inter3), .O(gate635inter10));
  nor2  gate1942(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate1943(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate1944(.a(gate635inter12), .b(gate635inter1), .O(N2040));
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );

  xor2  gate1833(.a(N2022), .b(N2039), .O(gate642inter0));
  nand2 gate1834(.a(gate642inter0), .b(s_136), .O(gate642inter1));
  and2  gate1835(.a(N2022), .b(N2039), .O(gate642inter2));
  inv1  gate1836(.a(s_136), .O(gate642inter3));
  inv1  gate1837(.a(s_137), .O(gate642inter4));
  nand2 gate1838(.a(gate642inter4), .b(gate642inter3), .O(gate642inter5));
  nor2  gate1839(.a(gate642inter5), .b(gate642inter2), .O(gate642inter6));
  inv1  gate1840(.a(N2039), .O(gate642inter7));
  inv1  gate1841(.a(N2022), .O(gate642inter8));
  nand2 gate1842(.a(gate642inter8), .b(gate642inter7), .O(gate642inter9));
  nand2 gate1843(.a(s_137), .b(gate642inter3), .O(gate642inter10));
  nor2  gate1844(.a(gate642inter10), .b(gate642inter9), .O(gate642inter11));
  nor2  gate1845(.a(gate642inter11), .b(gate642inter6), .O(gate642inter12));
  nand2 gate1846(.a(gate642inter12), .b(gate642inter1), .O(N2061));

  xor2  gate1371(.a(N290), .b(N2040), .O(gate643inter0));
  nand2 gate1372(.a(gate643inter0), .b(s_70), .O(gate643inter1));
  and2  gate1373(.a(N290), .b(N2040), .O(gate643inter2));
  inv1  gate1374(.a(s_70), .O(gate643inter3));
  inv1  gate1375(.a(s_71), .O(gate643inter4));
  nand2 gate1376(.a(gate643inter4), .b(gate643inter3), .O(gate643inter5));
  nor2  gate1377(.a(gate643inter5), .b(gate643inter2), .O(gate643inter6));
  inv1  gate1378(.a(N2040), .O(gate643inter7));
  inv1  gate1379(.a(N290), .O(gate643inter8));
  nand2 gate1380(.a(gate643inter8), .b(gate643inter7), .O(gate643inter9));
  nand2 gate1381(.a(s_71), .b(gate643inter3), .O(gate643inter10));
  nor2  gate1382(.a(gate643inter10), .b(gate643inter9), .O(gate643inter11));
  nor2  gate1383(.a(gate643inter11), .b(gate643inter6), .O(gate643inter12));
  nand2 gate1384(.a(gate643inter12), .b(gate643inter1), .O(N2062));
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );

  xor2  gate1903(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate1904(.a(gate678inter0), .b(s_146), .O(gate678inter1));
  and2  gate1905(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate1906(.a(s_146), .O(gate678inter3));
  inv1  gate1907(.a(s_147), .O(gate678inter4));
  nand2 gate1908(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate1909(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate1910(.a(N1252), .O(gate678inter7));
  inv1  gate1911(.a(N2225), .O(gate678inter8));
  nand2 gate1912(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate1913(.a(s_147), .b(gate678inter3), .O(gate678inter10));
  nor2  gate1914(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate1915(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate1916(.a(gate678inter12), .b(gate678inter1), .O(N2233));
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );

  xor2  gate1693(.a(N2229), .b(N658), .O(gate680inter0));
  nand2 gate1694(.a(gate680inter0), .b(s_116), .O(gate680inter1));
  and2  gate1695(.a(N2229), .b(N658), .O(gate680inter2));
  inv1  gate1696(.a(s_116), .O(gate680inter3));
  inv1  gate1697(.a(s_117), .O(gate680inter4));
  nand2 gate1698(.a(gate680inter4), .b(gate680inter3), .O(gate680inter5));
  nor2  gate1699(.a(gate680inter5), .b(gate680inter2), .O(gate680inter6));
  inv1  gate1700(.a(N658), .O(gate680inter7));
  inv1  gate1701(.a(N2229), .O(gate680inter8));
  nand2 gate1702(.a(gate680inter8), .b(gate680inter7), .O(gate680inter9));
  nand2 gate1703(.a(s_117), .b(gate680inter3), .O(gate680inter10));
  nor2  gate1704(.a(gate680inter10), .b(gate680inter9), .O(gate680inter11));
  nor2  gate1705(.a(gate680inter11), .b(gate680inter6), .O(gate680inter12));
  nand2 gate1706(.a(gate680inter12), .b(gate680inter1), .O(N2235));
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );

  xor2  gate979(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate980(.a(gate684inter0), .b(s_14), .O(gate684inter1));
  and2  gate981(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate982(.a(s_14), .O(gate684inter3));
  inv1  gate983(.a(s_15), .O(gate684inter4));
  nand2 gate984(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate985(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate986(.a(N2224), .O(gate684inter7));
  inv1  gate987(.a(N2233), .O(gate684inter8));
  nand2 gate988(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate989(.a(s_15), .b(gate684inter3), .O(gate684inter10));
  nor2  gate990(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate991(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate992(.a(gate684inter12), .b(gate684inter1), .O(N2241));

  xor2  gate1665(.a(N2234), .b(N2226), .O(gate685inter0));
  nand2 gate1666(.a(gate685inter0), .b(s_112), .O(gate685inter1));
  and2  gate1667(.a(N2234), .b(N2226), .O(gate685inter2));
  inv1  gate1668(.a(s_112), .O(gate685inter3));
  inv1  gate1669(.a(s_113), .O(gate685inter4));
  nand2 gate1670(.a(gate685inter4), .b(gate685inter3), .O(gate685inter5));
  nor2  gate1671(.a(gate685inter5), .b(gate685inter2), .O(gate685inter6));
  inv1  gate1672(.a(N2226), .O(gate685inter7));
  inv1  gate1673(.a(N2234), .O(gate685inter8));
  nand2 gate1674(.a(gate685inter8), .b(gate685inter7), .O(gate685inter9));
  nand2 gate1675(.a(s_113), .b(gate685inter3), .O(gate685inter10));
  nor2  gate1676(.a(gate685inter10), .b(gate685inter9), .O(gate685inter11));
  nor2  gate1677(.a(gate685inter11), .b(gate685inter6), .O(gate685inter12));
  nand2 gate1678(.a(gate685inter12), .b(gate685inter1), .O(N2244));
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );

  xor2  gate909(.a(N534), .b(N2558), .O(gate750inter0));
  nand2 gate910(.a(gate750inter0), .b(s_4), .O(gate750inter1));
  and2  gate911(.a(N534), .b(N2558), .O(gate750inter2));
  inv1  gate912(.a(s_4), .O(gate750inter3));
  inv1  gate913(.a(s_5), .O(gate750inter4));
  nand2 gate914(.a(gate750inter4), .b(gate750inter3), .O(gate750inter5));
  nor2  gate915(.a(gate750inter5), .b(gate750inter2), .O(gate750inter6));
  inv1  gate916(.a(N2558), .O(gate750inter7));
  inv1  gate917(.a(N534), .O(gate750inter8));
  nand2 gate918(.a(gate750inter8), .b(gate750inter7), .O(gate750inter9));
  nand2 gate919(.a(s_5), .b(gate750inter3), .O(gate750inter10));
  nor2  gate920(.a(gate750inter10), .b(gate750inter9), .O(gate750inter11));
  nor2  gate921(.a(gate750inter11), .b(gate750inter6), .O(gate750inter12));
  nand2 gate922(.a(gate750inter12), .b(gate750inter1), .O(N2669));
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate1203(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate1204(.a(gate754inter0), .b(s_46), .O(gate754inter1));
  and2  gate1205(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate1206(.a(s_46), .O(gate754inter3));
  inv1  gate1207(.a(s_47), .O(gate754inter4));
  nand2 gate1208(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1209(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1210(.a(N2564), .O(gate754inter7));
  inv1  gate1211(.a(N536), .O(gate754inter8));
  nand2 gate1212(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1213(.a(s_47), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1214(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1215(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1216(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );

  xor2  gate1189(.a(N543), .b(N2570), .O(gate758inter0));
  nand2 gate1190(.a(gate758inter0), .b(s_44), .O(gate758inter1));
  and2  gate1191(.a(N543), .b(N2570), .O(gate758inter2));
  inv1  gate1192(.a(s_44), .O(gate758inter3));
  inv1  gate1193(.a(s_45), .O(gate758inter4));
  nand2 gate1194(.a(gate758inter4), .b(gate758inter3), .O(gate758inter5));
  nor2  gate1195(.a(gate758inter5), .b(gate758inter2), .O(gate758inter6));
  inv1  gate1196(.a(N2570), .O(gate758inter7));
  inv1  gate1197(.a(N543), .O(gate758inter8));
  nand2 gate1198(.a(gate758inter8), .b(gate758inter7), .O(gate758inter9));
  nand2 gate1199(.a(s_45), .b(gate758inter3), .O(gate758inter10));
  nor2  gate1200(.a(gate758inter10), .b(gate758inter9), .O(gate758inter11));
  nor2  gate1201(.a(gate758inter11), .b(gate758inter6), .O(gate758inter12));
  nand2 gate1202(.a(gate758inter12), .b(gate758inter1), .O(N2682));
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );

  xor2  gate2029(.a(N2670), .b(N343), .O(gate765inter0));
  nand2 gate2030(.a(gate765inter0), .b(s_164), .O(gate765inter1));
  and2  gate2031(.a(N2670), .b(N343), .O(gate765inter2));
  inv1  gate2032(.a(s_164), .O(gate765inter3));
  inv1  gate2033(.a(s_165), .O(gate765inter4));
  nand2 gate2034(.a(gate765inter4), .b(gate765inter3), .O(gate765inter5));
  nor2  gate2035(.a(gate765inter5), .b(gate765inter2), .O(gate765inter6));
  inv1  gate2036(.a(N343), .O(gate765inter7));
  inv1  gate2037(.a(N2670), .O(gate765inter8));
  nand2 gate2038(.a(gate765inter8), .b(gate765inter7), .O(gate765inter9));
  nand2 gate2039(.a(s_165), .b(gate765inter3), .O(gate765inter10));
  nor2  gate2040(.a(gate765inter10), .b(gate765inter9), .O(gate765inter11));
  nor2  gate2041(.a(gate765inter11), .b(gate765inter6), .O(gate765inter12));
  nand2 gate2042(.a(gate765inter12), .b(gate765inter1), .O(N2720));
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );

  xor2  gate881(.a(N2674), .b(N349), .O(gate767inter0));
  nand2 gate882(.a(gate767inter0), .b(s_0), .O(gate767inter1));
  and2  gate883(.a(N2674), .b(N349), .O(gate767inter2));
  inv1  gate884(.a(s_0), .O(gate767inter3));
  inv1  gate885(.a(s_1), .O(gate767inter4));
  nand2 gate886(.a(gate767inter4), .b(gate767inter3), .O(gate767inter5));
  nor2  gate887(.a(gate767inter5), .b(gate767inter2), .O(gate767inter6));
  inv1  gate888(.a(N349), .O(gate767inter7));
  inv1  gate889(.a(N2674), .O(gate767inter8));
  nand2 gate890(.a(gate767inter8), .b(gate767inter7), .O(gate767inter9));
  nand2 gate891(.a(s_1), .b(gate767inter3), .O(gate767inter10));
  nor2  gate892(.a(gate767inter10), .b(gate767inter9), .O(gate767inter11));
  nor2  gate893(.a(gate767inter11), .b(gate767inter6), .O(gate767inter12));
  nand2 gate894(.a(gate767inter12), .b(gate767inter1), .O(N2722));
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );

  xor2  gate1651(.a(N539), .b(N2642), .O(gate771inter0));
  nand2 gate1652(.a(gate771inter0), .b(s_110), .O(gate771inter1));
  and2  gate1653(.a(N539), .b(N2642), .O(gate771inter2));
  inv1  gate1654(.a(s_110), .O(gate771inter3));
  inv1  gate1655(.a(s_111), .O(gate771inter4));
  nand2 gate1656(.a(gate771inter4), .b(gate771inter3), .O(gate771inter5));
  nor2  gate1657(.a(gate771inter5), .b(gate771inter2), .O(gate771inter6));
  inv1  gate1658(.a(N2642), .O(gate771inter7));
  inv1  gate1659(.a(N539), .O(gate771inter8));
  nand2 gate1660(.a(gate771inter8), .b(gate771inter7), .O(gate771inter9));
  nand2 gate1661(.a(s_111), .b(gate771inter3), .O(gate771inter10));
  nor2  gate1662(.a(gate771inter10), .b(gate771inter9), .O(gate771inter11));
  nor2  gate1663(.a(gate771inter11), .b(gate771inter6), .O(gate771inter12));
  nand2 gate1664(.a(gate771inter12), .b(gate771inter1), .O(N2726));
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );

  xor2  gate1945(.a(N542), .b(N2651), .O(gate777inter0));
  nand2 gate1946(.a(gate777inter0), .b(s_152), .O(gate777inter1));
  and2  gate1947(.a(N542), .b(N2651), .O(gate777inter2));
  inv1  gate1948(.a(s_152), .O(gate777inter3));
  inv1  gate1949(.a(s_153), .O(gate777inter4));
  nand2 gate1950(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate1951(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate1952(.a(N2651), .O(gate777inter7));
  inv1  gate1953(.a(N542), .O(gate777inter8));
  nand2 gate1954(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate1955(.a(s_153), .b(gate777inter3), .O(gate777inter10));
  nor2  gate1956(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate1957(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate1958(.a(gate777inter12), .b(gate777inter1), .O(N2732));
inv1 gate778( .a(N2651), .O(N2733) );

  xor2  gate1721(.a(N2683), .b(N370), .O(gate779inter0));
  nand2 gate1722(.a(gate779inter0), .b(s_120), .O(gate779inter1));
  and2  gate1723(.a(N2683), .b(N370), .O(gate779inter2));
  inv1  gate1724(.a(s_120), .O(gate779inter3));
  inv1  gate1725(.a(s_121), .O(gate779inter4));
  nand2 gate1726(.a(gate779inter4), .b(gate779inter3), .O(gate779inter5));
  nor2  gate1727(.a(gate779inter5), .b(gate779inter2), .O(gate779inter6));
  inv1  gate1728(.a(N370), .O(gate779inter7));
  inv1  gate1729(.a(N2683), .O(gate779inter8));
  nand2 gate1730(.a(gate779inter8), .b(gate779inter7), .O(gate779inter9));
  nand2 gate1731(.a(s_121), .b(gate779inter3), .O(gate779inter10));
  nor2  gate1732(.a(gate779inter10), .b(gate779inter9), .O(gate779inter11));
  nor2  gate1733(.a(gate779inter11), .b(gate779inter6), .O(gate779inter12));
  nand2 gate1734(.a(gate779inter12), .b(gate779inter1), .O(N2734));
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );

  xor2  gate1273(.a(N546), .b(N2661), .O(gate784inter0));
  nand2 gate1274(.a(gate784inter0), .b(s_56), .O(gate784inter1));
  and2  gate1275(.a(N546), .b(N2661), .O(gate784inter2));
  inv1  gate1276(.a(s_56), .O(gate784inter3));
  inv1  gate1277(.a(s_57), .O(gate784inter4));
  nand2 gate1278(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate1279(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate1280(.a(N2661), .O(gate784inter7));
  inv1  gate1281(.a(N546), .O(gate784inter8));
  nand2 gate1282(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate1283(.a(s_57), .b(gate784inter3), .O(gate784inter10));
  nor2  gate1284(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate1285(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate1286(.a(gate784inter12), .b(gate784inter1), .O(N2739));
inv1 gate785( .a(N2661), .O(N2740) );

  xor2  gate1497(.a(N547), .b(N2664), .O(gate786inter0));
  nand2 gate1498(.a(gate786inter0), .b(s_88), .O(gate786inter1));
  and2  gate1499(.a(N547), .b(N2664), .O(gate786inter2));
  inv1  gate1500(.a(s_88), .O(gate786inter3));
  inv1  gate1501(.a(s_89), .O(gate786inter4));
  nand2 gate1502(.a(gate786inter4), .b(gate786inter3), .O(gate786inter5));
  nor2  gate1503(.a(gate786inter5), .b(gate786inter2), .O(gate786inter6));
  inv1  gate1504(.a(N2664), .O(gate786inter7));
  inv1  gate1505(.a(N547), .O(gate786inter8));
  nand2 gate1506(.a(gate786inter8), .b(gate786inter7), .O(gate786inter9));
  nand2 gate1507(.a(s_89), .b(gate786inter3), .O(gate786inter10));
  nor2  gate1508(.a(gate786inter10), .b(gate786inter9), .O(gate786inter11));
  nor2  gate1509(.a(gate786inter11), .b(gate786inter6), .O(gate786inter12));
  nand2 gate1510(.a(gate786inter12), .b(gate786inter1), .O(N2741));
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate1427(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate1428(.a(gate788inter0), .b(s_78), .O(gate788inter1));
  and2  gate1429(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate1430(.a(s_78), .O(gate788inter3));
  inv1  gate1431(.a(s_79), .O(gate788inter4));
  nand2 gate1432(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate1433(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate1434(.a(N385), .O(gate788inter7));
  inv1  gate1435(.a(N2689), .O(gate788inter8));
  nand2 gate1436(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate1437(.a(s_79), .b(gate788inter3), .O(gate788inter10));
  nor2  gate1438(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate1439(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate1440(.a(gate788inter12), .b(gate788inter1), .O(N2743));
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );

  xor2  gate965(.a(N2723), .b(N2675), .O(gate797inter0));
  nand2 gate966(.a(gate797inter0), .b(s_12), .O(gate797inter1));
  and2  gate967(.a(N2723), .b(N2675), .O(gate797inter2));
  inv1  gate968(.a(s_12), .O(gate797inter3));
  inv1  gate969(.a(s_13), .O(gate797inter4));
  nand2 gate970(.a(gate797inter4), .b(gate797inter3), .O(gate797inter5));
  nor2  gate971(.a(gate797inter5), .b(gate797inter2), .O(gate797inter6));
  inv1  gate972(.a(N2675), .O(gate797inter7));
  inv1  gate973(.a(N2723), .O(gate797inter8));
  nand2 gate974(.a(gate797inter8), .b(gate797inter7), .O(gate797inter9));
  nand2 gate975(.a(s_13), .b(gate797inter3), .O(gate797inter10));
  nor2  gate976(.a(gate797inter10), .b(gate797inter9), .O(gate797inter11));
  nor2  gate977(.a(gate797inter11), .b(gate797inter6), .O(gate797inter12));
  nand2 gate978(.a(gate797inter12), .b(gate797inter1), .O(N2756));

  xor2  gate1987(.a(N2725), .b(N355), .O(gate798inter0));
  nand2 gate1988(.a(gate798inter0), .b(s_158), .O(gate798inter1));
  and2  gate1989(.a(N2725), .b(N355), .O(gate798inter2));
  inv1  gate1990(.a(s_158), .O(gate798inter3));
  inv1  gate1991(.a(s_159), .O(gate798inter4));
  nand2 gate1992(.a(gate798inter4), .b(gate798inter3), .O(gate798inter5));
  nor2  gate1993(.a(gate798inter5), .b(gate798inter2), .O(gate798inter6));
  inv1  gate1994(.a(N355), .O(gate798inter7));
  inv1  gate1995(.a(N2725), .O(gate798inter8));
  nand2 gate1996(.a(gate798inter8), .b(gate798inter7), .O(gate798inter9));
  nand2 gate1997(.a(s_159), .b(gate798inter3), .O(gate798inter10));
  nor2  gate1998(.a(gate798inter10), .b(gate798inter9), .O(gate798inter11));
  nor2  gate1999(.a(gate798inter11), .b(gate798inter6), .O(gate798inter12));
  nand2 gate2000(.a(gate798inter12), .b(gate798inter1), .O(N2757));

  xor2  gate1357(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate1358(.a(gate799inter0), .b(s_68), .O(gate799inter1));
  and2  gate1359(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate1360(.a(s_68), .O(gate799inter3));
  inv1  gate1361(.a(s_69), .O(gate799inter4));
  nand2 gate1362(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate1363(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate1364(.a(N358), .O(gate799inter7));
  inv1  gate1365(.a(N2727), .O(gate799inter8));
  nand2 gate1366(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate1367(.a(s_69), .b(gate799inter3), .O(gate799inter10));
  nor2  gate1368(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate1369(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate1370(.a(gate799inter12), .b(gate799inter1), .O(N2758));

  xor2  gate1749(.a(N2729), .b(N361), .O(gate800inter0));
  nand2 gate1750(.a(gate800inter0), .b(s_124), .O(gate800inter1));
  and2  gate1751(.a(N2729), .b(N361), .O(gate800inter2));
  inv1  gate1752(.a(s_124), .O(gate800inter3));
  inv1  gate1753(.a(s_125), .O(gate800inter4));
  nand2 gate1754(.a(gate800inter4), .b(gate800inter3), .O(gate800inter5));
  nor2  gate1755(.a(gate800inter5), .b(gate800inter2), .O(gate800inter6));
  inv1  gate1756(.a(N361), .O(gate800inter7));
  inv1  gate1757(.a(N2729), .O(gate800inter8));
  nand2 gate1758(.a(gate800inter8), .b(gate800inter7), .O(gate800inter9));
  nand2 gate1759(.a(s_125), .b(gate800inter3), .O(gate800inter10));
  nor2  gate1760(.a(gate800inter10), .b(gate800inter9), .O(gate800inter11));
  nor2  gate1761(.a(gate800inter11), .b(gate800inter6), .O(gate800inter12));
  nand2 gate1762(.a(gate800inter12), .b(gate800inter1), .O(N2759));
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );

  xor2  gate1539(.a(N2736), .b(N373), .O(gate804inter0));
  nand2 gate1540(.a(gate804inter0), .b(s_94), .O(gate804inter1));
  and2  gate1541(.a(N2736), .b(N373), .O(gate804inter2));
  inv1  gate1542(.a(s_94), .O(gate804inter3));
  inv1  gate1543(.a(s_95), .O(gate804inter4));
  nand2 gate1544(.a(gate804inter4), .b(gate804inter3), .O(gate804inter5));
  nor2  gate1545(.a(gate804inter5), .b(gate804inter2), .O(gate804inter6));
  inv1  gate1546(.a(N373), .O(gate804inter7));
  inv1  gate1547(.a(N2736), .O(gate804inter8));
  nand2 gate1548(.a(gate804inter8), .b(gate804inter7), .O(gate804inter9));
  nand2 gate1549(.a(s_95), .b(gate804inter3), .O(gate804inter10));
  nor2  gate1550(.a(gate804inter10), .b(gate804inter9), .O(gate804inter11));
  nor2  gate1551(.a(gate804inter11), .b(gate804inter6), .O(gate804inter12));
  nand2 gate1552(.a(gate804inter12), .b(gate804inter1), .O(N2763));
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );

  xor2  gate1861(.a(N2742), .b(N382), .O(gate807inter0));
  nand2 gate1862(.a(gate807inter0), .b(s_140), .O(gate807inter1));
  and2  gate1863(.a(N2742), .b(N382), .O(gate807inter2));
  inv1  gate1864(.a(s_140), .O(gate807inter3));
  inv1  gate1865(.a(s_141), .O(gate807inter4));
  nand2 gate1866(.a(gate807inter4), .b(gate807inter3), .O(gate807inter5));
  nor2  gate1867(.a(gate807inter5), .b(gate807inter2), .O(gate807inter6));
  inv1  gate1868(.a(N382), .O(gate807inter7));
  inv1  gate1869(.a(N2742), .O(gate807inter8));
  nand2 gate1870(.a(gate807inter8), .b(gate807inter7), .O(gate807inter9));
  nand2 gate1871(.a(s_141), .b(gate807inter3), .O(gate807inter10));
  nor2  gate1872(.a(gate807inter10), .b(gate807inter9), .O(gate807inter11));
  nor2  gate1873(.a(gate807inter11), .b(gate807inter6), .O(gate807inter12));
  nand2 gate1874(.a(gate807inter12), .b(gate807inter1), .O(N2766));
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );

  xor2  gate1091(.a(N2759), .b(N2728), .O(gate814inter0));
  nand2 gate1092(.a(gate814inter0), .b(s_30), .O(gate814inter1));
  and2  gate1093(.a(N2759), .b(N2728), .O(gate814inter2));
  inv1  gate1094(.a(s_30), .O(gate814inter3));
  inv1  gate1095(.a(s_31), .O(gate814inter4));
  nand2 gate1096(.a(gate814inter4), .b(gate814inter3), .O(gate814inter5));
  nor2  gate1097(.a(gate814inter5), .b(gate814inter2), .O(gate814inter6));
  inv1  gate1098(.a(N2728), .O(gate814inter7));
  inv1  gate1099(.a(N2759), .O(gate814inter8));
  nand2 gate1100(.a(gate814inter8), .b(gate814inter7), .O(gate814inter9));
  nand2 gate1101(.a(s_31), .b(gate814inter3), .O(gate814inter10));
  nor2  gate1102(.a(gate814inter10), .b(gate814inter9), .O(gate814inter11));
  nor2  gate1103(.a(gate814inter11), .b(gate814inter6), .O(gate814inter12));
  nand2 gate1104(.a(gate814inter12), .b(gate814inter1), .O(N2781));

  xor2  gate895(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate896(.a(gate815inter0), .b(s_2), .O(gate815inter1));
  and2  gate897(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate898(.a(s_2), .O(gate815inter3));
  inv1  gate899(.a(s_3), .O(gate815inter4));
  nand2 gate900(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate901(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate902(.a(N2730), .O(gate815inter7));
  inv1  gate903(.a(N2760), .O(gate815inter8));
  nand2 gate904(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate905(.a(s_3), .b(gate815inter3), .O(gate815inter10));
  nor2  gate906(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate907(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate908(.a(gate815inter12), .b(gate815inter1), .O(N2782));
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );

  xor2  gate1763(.a(N2764), .b(N2737), .O(gate818inter0));
  nand2 gate1764(.a(gate818inter0), .b(s_126), .O(gate818inter1));
  and2  gate1765(.a(N2764), .b(N2737), .O(gate818inter2));
  inv1  gate1766(.a(s_126), .O(gate818inter3));
  inv1  gate1767(.a(s_127), .O(gate818inter4));
  nand2 gate1768(.a(gate818inter4), .b(gate818inter3), .O(gate818inter5));
  nor2  gate1769(.a(gate818inter5), .b(gate818inter2), .O(gate818inter6));
  inv1  gate1770(.a(N2737), .O(gate818inter7));
  inv1  gate1771(.a(N2764), .O(gate818inter8));
  nand2 gate1772(.a(gate818inter8), .b(gate818inter7), .O(gate818inter9));
  nand2 gate1773(.a(s_127), .b(gate818inter3), .O(gate818inter10));
  nor2  gate1774(.a(gate818inter10), .b(gate818inter9), .O(gate818inter11));
  nor2  gate1775(.a(gate818inter11), .b(gate818inter6), .O(gate818inter12));
  nand2 gate1776(.a(gate818inter12), .b(gate818inter1), .O(N2785));
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );

  xor2  gate1245(.a(N2808), .b(N1965), .O(gate834inter0));
  nand2 gate1246(.a(gate834inter0), .b(s_52), .O(gate834inter1));
  and2  gate1247(.a(N2808), .b(N1965), .O(gate834inter2));
  inv1  gate1248(.a(s_52), .O(gate834inter3));
  inv1  gate1249(.a(s_53), .O(gate834inter4));
  nand2 gate1250(.a(gate834inter4), .b(gate834inter3), .O(gate834inter5));
  nor2  gate1251(.a(gate834inter5), .b(gate834inter2), .O(gate834inter6));
  inv1  gate1252(.a(N1965), .O(gate834inter7));
  inv1  gate1253(.a(N2808), .O(gate834inter8));
  nand2 gate1254(.a(gate834inter8), .b(gate834inter7), .O(gate834inter9));
  nand2 gate1255(.a(s_53), .b(gate834inter3), .O(gate834inter10));
  nor2  gate1256(.a(gate834inter10), .b(gate834inter9), .O(gate834inter11));
  nor2  gate1257(.a(gate834inter11), .b(gate834inter6), .O(gate834inter12));
  nand2 gate1258(.a(gate834inter12), .b(gate834inter1), .O(N2827));
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );

  xor2  gate1707(.a(N1857), .b(N2821), .O(gate842inter0));
  nand2 gate1708(.a(gate842inter0), .b(s_118), .O(gate842inter1));
  and2  gate1709(.a(N1857), .b(N2821), .O(gate842inter2));
  inv1  gate1710(.a(s_118), .O(gate842inter3));
  inv1  gate1711(.a(s_119), .O(gate842inter4));
  nand2 gate1712(.a(gate842inter4), .b(gate842inter3), .O(gate842inter5));
  nor2  gate1713(.a(gate842inter5), .b(gate842inter2), .O(gate842inter6));
  inv1  gate1714(.a(N2821), .O(gate842inter7));
  inv1  gate1715(.a(N1857), .O(gate842inter8));
  nand2 gate1716(.a(gate842inter8), .b(gate842inter7), .O(gate842inter9));
  nand2 gate1717(.a(s_119), .b(gate842inter3), .O(gate842inter10));
  nor2  gate1718(.a(gate842inter10), .b(gate842inter9), .O(gate842inter11));
  nor2  gate1719(.a(gate842inter11), .b(gate842inter6), .O(gate842inter12));
  nand2 gate1720(.a(gate842inter12), .b(gate842inter1), .O(N2853));
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );

  xor2  gate1917(.a(N2861), .b(N1902), .O(gate855inter0));
  nand2 gate1918(.a(gate855inter0), .b(s_148), .O(gate855inter1));
  and2  gate1919(.a(N2861), .b(N1902), .O(gate855inter2));
  inv1  gate1920(.a(s_148), .O(gate855inter3));
  inv1  gate1921(.a(s_149), .O(gate855inter4));
  nand2 gate1922(.a(gate855inter4), .b(gate855inter3), .O(gate855inter5));
  nor2  gate1923(.a(gate855inter5), .b(gate855inter2), .O(gate855inter6));
  inv1  gate1924(.a(N1902), .O(gate855inter7));
  inv1  gate1925(.a(N2861), .O(gate855inter8));
  nand2 gate1926(.a(gate855inter8), .b(gate855inter7), .O(gate855inter9));
  nand2 gate1927(.a(s_149), .b(gate855inter3), .O(gate855inter10));
  nor2  gate1928(.a(gate855inter10), .b(gate855inter9), .O(gate855inter11));
  nor2  gate1929(.a(gate855inter11), .b(gate855inter6), .O(gate855inter12));
  nand2 gate1930(.a(gate855inter12), .b(gate855inter1), .O(N2870));
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );

  xor2  gate2043(.a(N2853), .b(N2869), .O(gate864inter0));
  nand2 gate2044(.a(gate864inter0), .b(s_166), .O(gate864inter1));
  and2  gate2045(.a(N2853), .b(N2869), .O(gate864inter2));
  inv1  gate2046(.a(s_166), .O(gate864inter3));
  inv1  gate2047(.a(s_167), .O(gate864inter4));
  nand2 gate2048(.a(gate864inter4), .b(gate864inter3), .O(gate864inter5));
  nor2  gate2049(.a(gate864inter5), .b(gate864inter2), .O(gate864inter6));
  inv1  gate2050(.a(N2869), .O(gate864inter7));
  inv1  gate2051(.a(N2853), .O(gate864inter8));
  nand2 gate2052(.a(gate864inter8), .b(gate864inter7), .O(gate864inter9));
  nand2 gate2053(.a(s_167), .b(gate864inter3), .O(gate864inter10));
  nor2  gate2054(.a(gate864inter10), .b(gate864inter9), .O(gate864inter11));
  nor2  gate2055(.a(gate864inter11), .b(gate864inter6), .O(gate864inter12));
  nand2 gate2056(.a(gate864inter12), .b(gate864inter1), .O(N2879));
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );

  xor2  gate937(.a(N2872), .b(N682), .O(gate866inter0));
  nand2 gate938(.a(gate866inter0), .b(s_8), .O(gate866inter1));
  and2  gate939(.a(N2872), .b(N682), .O(gate866inter2));
  inv1  gate940(.a(s_8), .O(gate866inter3));
  inv1  gate941(.a(s_9), .O(gate866inter4));
  nand2 gate942(.a(gate866inter4), .b(gate866inter3), .O(gate866inter5));
  nor2  gate943(.a(gate866inter5), .b(gate866inter2), .O(gate866inter6));
  inv1  gate944(.a(N682), .O(gate866inter7));
  inv1  gate945(.a(N2872), .O(gate866inter8));
  nand2 gate946(.a(gate866inter8), .b(gate866inter7), .O(gate866inter9));
  nand2 gate947(.a(s_9), .b(gate866inter3), .O(gate866inter10));
  nor2  gate948(.a(gate866inter10), .b(gate866inter9), .O(gate866inter11));
  nor2  gate949(.a(gate866inter11), .b(gate866inter6), .O(gate866inter12));
  nand2 gate950(.a(gate866inter12), .b(gate866inter1), .O(N2881));

  xor2  gate1315(.a(N2874), .b(N685), .O(gate867inter0));
  nand2 gate1316(.a(gate867inter0), .b(s_62), .O(gate867inter1));
  and2  gate1317(.a(N2874), .b(N685), .O(gate867inter2));
  inv1  gate1318(.a(s_62), .O(gate867inter3));
  inv1  gate1319(.a(s_63), .O(gate867inter4));
  nand2 gate1320(.a(gate867inter4), .b(gate867inter3), .O(gate867inter5));
  nor2  gate1321(.a(gate867inter5), .b(gate867inter2), .O(gate867inter6));
  inv1  gate1322(.a(N685), .O(gate867inter7));
  inv1  gate1323(.a(N2874), .O(gate867inter8));
  nand2 gate1324(.a(gate867inter8), .b(gate867inter7), .O(gate867inter9));
  nand2 gate1325(.a(s_63), .b(gate867inter3), .O(gate867inter10));
  nor2  gate1326(.a(gate867inter10), .b(gate867inter9), .O(gate867inter11));
  nor2  gate1327(.a(gate867inter11), .b(gate867inter6), .O(gate867inter12));
  nand2 gate1328(.a(gate867inter12), .b(gate867inter1), .O(N2882));
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate1679(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate1680(.a(gate874inter0), .b(s_114), .O(gate874inter1));
  and2  gate1681(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate1682(.a(s_114), .O(gate874inter3));
  inv1  gate1683(.a(s_115), .O(gate874inter4));
  nand2 gate1684(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate1685(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate1686(.a(N2871), .O(gate874inter7));
  inv1  gate1687(.a(N2881), .O(gate874inter8));
  nand2 gate1688(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate1689(.a(s_115), .b(gate874inter3), .O(gate874inter10));
  nor2  gate1690(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate1691(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate1692(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );

  xor2  gate1889(.a(N2897), .b(N2895), .O(gate879inter0));
  nand2 gate1890(.a(gate879inter0), .b(s_144), .O(gate879inter1));
  and2  gate1891(.a(N2897), .b(N2895), .O(gate879inter2));
  inv1  gate1892(.a(s_144), .O(gate879inter3));
  inv1  gate1893(.a(s_145), .O(gate879inter4));
  nand2 gate1894(.a(gate879inter4), .b(gate879inter3), .O(gate879inter5));
  nor2  gate1895(.a(gate879inter5), .b(gate879inter2), .O(gate879inter6));
  inv1  gate1896(.a(N2895), .O(gate879inter7));
  inv1  gate1897(.a(N2897), .O(gate879inter8));
  nand2 gate1898(.a(gate879inter8), .b(gate879inter7), .O(gate879inter9));
  nand2 gate1899(.a(s_145), .b(gate879inter3), .O(gate879inter10));
  nor2  gate1900(.a(gate879inter10), .b(gate879inter9), .O(gate879inter11));
  nor2  gate1901(.a(gate879inter11), .b(gate879inter6), .O(gate879inter12));
  nand2 gate1902(.a(gate879inter12), .b(gate879inter1), .O(N2898));
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule