module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1835(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1836(.a(gate11inter0), .b(s_184), .O(gate11inter1));
  and2  gate1837(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1838(.a(s_184), .O(gate11inter3));
  inv1  gate1839(.a(s_185), .O(gate11inter4));
  nand2 gate1840(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1841(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1842(.a(G5), .O(gate11inter7));
  inv1  gate1843(.a(G6), .O(gate11inter8));
  nand2 gate1844(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1845(.a(s_185), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1846(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1847(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1848(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate659(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate660(.a(gate13inter0), .b(s_16), .O(gate13inter1));
  and2  gate661(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate662(.a(s_16), .O(gate13inter3));
  inv1  gate663(.a(s_17), .O(gate13inter4));
  nand2 gate664(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate665(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate666(.a(G9), .O(gate13inter7));
  inv1  gate667(.a(G10), .O(gate13inter8));
  nand2 gate668(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate669(.a(s_17), .b(gate13inter3), .O(gate13inter10));
  nor2  gate670(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate671(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate672(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1639(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1640(.a(gate16inter0), .b(s_156), .O(gate16inter1));
  and2  gate1641(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1642(.a(s_156), .O(gate16inter3));
  inv1  gate1643(.a(s_157), .O(gate16inter4));
  nand2 gate1644(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1645(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1646(.a(G15), .O(gate16inter7));
  inv1  gate1647(.a(G16), .O(gate16inter8));
  nand2 gate1648(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1649(.a(s_157), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1650(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1651(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1652(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1415(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1416(.a(gate23inter0), .b(s_124), .O(gate23inter1));
  and2  gate1417(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1418(.a(s_124), .O(gate23inter3));
  inv1  gate1419(.a(s_125), .O(gate23inter4));
  nand2 gate1420(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1421(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1422(.a(G29), .O(gate23inter7));
  inv1  gate1423(.a(G30), .O(gate23inter8));
  nand2 gate1424(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1425(.a(s_125), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1426(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1427(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1428(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate2073(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2074(.a(gate30inter0), .b(s_218), .O(gate30inter1));
  and2  gate2075(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2076(.a(s_218), .O(gate30inter3));
  inv1  gate2077(.a(s_219), .O(gate30inter4));
  nand2 gate2078(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2079(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2080(.a(G11), .O(gate30inter7));
  inv1  gate2081(.a(G15), .O(gate30inter8));
  nand2 gate2082(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2083(.a(s_219), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2084(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2085(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2086(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate911(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate912(.a(gate35inter0), .b(s_52), .O(gate35inter1));
  and2  gate913(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate914(.a(s_52), .O(gate35inter3));
  inv1  gate915(.a(s_53), .O(gate35inter4));
  nand2 gate916(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate917(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate918(.a(G18), .O(gate35inter7));
  inv1  gate919(.a(G22), .O(gate35inter8));
  nand2 gate920(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate921(.a(s_53), .b(gate35inter3), .O(gate35inter10));
  nor2  gate922(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate923(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate924(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1401(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1402(.a(gate36inter0), .b(s_122), .O(gate36inter1));
  and2  gate1403(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1404(.a(s_122), .O(gate36inter3));
  inv1  gate1405(.a(s_123), .O(gate36inter4));
  nand2 gate1406(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1407(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1408(.a(G26), .O(gate36inter7));
  inv1  gate1409(.a(G30), .O(gate36inter8));
  nand2 gate1410(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1411(.a(s_123), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1412(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1413(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1414(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2157(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2158(.a(gate46inter0), .b(s_230), .O(gate46inter1));
  and2  gate2159(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2160(.a(s_230), .O(gate46inter3));
  inv1  gate2161(.a(s_231), .O(gate46inter4));
  nand2 gate2162(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2163(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2164(.a(G6), .O(gate46inter7));
  inv1  gate2165(.a(G272), .O(gate46inter8));
  nand2 gate2166(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2167(.a(s_231), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2168(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2169(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2170(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1261(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1262(.a(gate47inter0), .b(s_102), .O(gate47inter1));
  and2  gate1263(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1264(.a(s_102), .O(gate47inter3));
  inv1  gate1265(.a(s_103), .O(gate47inter4));
  nand2 gate1266(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1267(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1268(.a(G7), .O(gate47inter7));
  inv1  gate1269(.a(G275), .O(gate47inter8));
  nand2 gate1270(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1271(.a(s_103), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1272(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1273(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1274(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate771(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate772(.a(gate49inter0), .b(s_32), .O(gate49inter1));
  and2  gate773(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate774(.a(s_32), .O(gate49inter3));
  inv1  gate775(.a(s_33), .O(gate49inter4));
  nand2 gate776(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate777(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate778(.a(G9), .O(gate49inter7));
  inv1  gate779(.a(G278), .O(gate49inter8));
  nand2 gate780(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate781(.a(s_33), .b(gate49inter3), .O(gate49inter10));
  nor2  gate782(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate783(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate784(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2227(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2228(.a(gate51inter0), .b(s_240), .O(gate51inter1));
  and2  gate2229(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2230(.a(s_240), .O(gate51inter3));
  inv1  gate2231(.a(s_241), .O(gate51inter4));
  nand2 gate2232(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2233(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2234(.a(G11), .O(gate51inter7));
  inv1  gate2235(.a(G281), .O(gate51inter8));
  nand2 gate2236(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2237(.a(s_241), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2238(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2239(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2240(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1443(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1444(.a(gate52inter0), .b(s_128), .O(gate52inter1));
  and2  gate1445(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1446(.a(s_128), .O(gate52inter3));
  inv1  gate1447(.a(s_129), .O(gate52inter4));
  nand2 gate1448(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1449(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1450(.a(G12), .O(gate52inter7));
  inv1  gate1451(.a(G281), .O(gate52inter8));
  nand2 gate1452(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1453(.a(s_129), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1454(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1455(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1456(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate729(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate730(.a(gate57inter0), .b(s_26), .O(gate57inter1));
  and2  gate731(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate732(.a(s_26), .O(gate57inter3));
  inv1  gate733(.a(s_27), .O(gate57inter4));
  nand2 gate734(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate735(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate736(.a(G17), .O(gate57inter7));
  inv1  gate737(.a(G290), .O(gate57inter8));
  nand2 gate738(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate739(.a(s_27), .b(gate57inter3), .O(gate57inter10));
  nor2  gate740(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate741(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate742(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1345(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1346(.a(gate58inter0), .b(s_114), .O(gate58inter1));
  and2  gate1347(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1348(.a(s_114), .O(gate58inter3));
  inv1  gate1349(.a(s_115), .O(gate58inter4));
  nand2 gate1350(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1351(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1352(.a(G18), .O(gate58inter7));
  inv1  gate1353(.a(G290), .O(gate58inter8));
  nand2 gate1354(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1355(.a(s_115), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1356(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1357(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1358(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate827(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate828(.a(gate59inter0), .b(s_40), .O(gate59inter1));
  and2  gate829(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate830(.a(s_40), .O(gate59inter3));
  inv1  gate831(.a(s_41), .O(gate59inter4));
  nand2 gate832(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate833(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate834(.a(G19), .O(gate59inter7));
  inv1  gate835(.a(G293), .O(gate59inter8));
  nand2 gate836(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate837(.a(s_41), .b(gate59inter3), .O(gate59inter10));
  nor2  gate838(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate839(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate840(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate785(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate786(.a(gate64inter0), .b(s_34), .O(gate64inter1));
  and2  gate787(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate788(.a(s_34), .O(gate64inter3));
  inv1  gate789(.a(s_35), .O(gate64inter4));
  nand2 gate790(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate791(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate792(.a(G24), .O(gate64inter7));
  inv1  gate793(.a(G299), .O(gate64inter8));
  nand2 gate794(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate795(.a(s_35), .b(gate64inter3), .O(gate64inter10));
  nor2  gate796(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate797(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate798(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1779(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1780(.a(gate68inter0), .b(s_176), .O(gate68inter1));
  and2  gate1781(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1782(.a(s_176), .O(gate68inter3));
  inv1  gate1783(.a(s_177), .O(gate68inter4));
  nand2 gate1784(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1785(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1786(.a(G28), .O(gate68inter7));
  inv1  gate1787(.a(G305), .O(gate68inter8));
  nand2 gate1788(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1789(.a(s_177), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1790(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1791(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1792(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1457(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1458(.a(gate71inter0), .b(s_130), .O(gate71inter1));
  and2  gate1459(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1460(.a(s_130), .O(gate71inter3));
  inv1  gate1461(.a(s_131), .O(gate71inter4));
  nand2 gate1462(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1463(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1464(.a(G31), .O(gate71inter7));
  inv1  gate1465(.a(G311), .O(gate71inter8));
  nand2 gate1466(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1467(.a(s_131), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1468(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1469(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1470(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate813(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate814(.a(gate74inter0), .b(s_38), .O(gate74inter1));
  and2  gate815(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate816(.a(s_38), .O(gate74inter3));
  inv1  gate817(.a(s_39), .O(gate74inter4));
  nand2 gate818(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate819(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate820(.a(G5), .O(gate74inter7));
  inv1  gate821(.a(G314), .O(gate74inter8));
  nand2 gate822(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate823(.a(s_39), .b(gate74inter3), .O(gate74inter10));
  nor2  gate824(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate825(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate826(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1653(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1654(.a(gate76inter0), .b(s_158), .O(gate76inter1));
  and2  gate1655(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1656(.a(s_158), .O(gate76inter3));
  inv1  gate1657(.a(s_159), .O(gate76inter4));
  nand2 gate1658(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1659(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1660(.a(G13), .O(gate76inter7));
  inv1  gate1661(.a(G317), .O(gate76inter8));
  nand2 gate1662(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1663(.a(s_159), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1664(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1665(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1666(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1135(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1136(.a(gate80inter0), .b(s_84), .O(gate80inter1));
  and2  gate1137(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1138(.a(s_84), .O(gate80inter3));
  inv1  gate1139(.a(s_85), .O(gate80inter4));
  nand2 gate1140(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1141(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1142(.a(G14), .O(gate80inter7));
  inv1  gate1143(.a(G323), .O(gate80inter8));
  nand2 gate1144(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1145(.a(s_85), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1146(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1147(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1148(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate995(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate996(.a(gate85inter0), .b(s_64), .O(gate85inter1));
  and2  gate997(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate998(.a(s_64), .O(gate85inter3));
  inv1  gate999(.a(s_65), .O(gate85inter4));
  nand2 gate1000(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1001(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1002(.a(G4), .O(gate85inter7));
  inv1  gate1003(.a(G332), .O(gate85inter8));
  nand2 gate1004(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1005(.a(s_65), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1006(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1007(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1008(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1737(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1738(.a(gate88inter0), .b(s_170), .O(gate88inter1));
  and2  gate1739(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1740(.a(s_170), .O(gate88inter3));
  inv1  gate1741(.a(s_171), .O(gate88inter4));
  nand2 gate1742(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1743(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1744(.a(G16), .O(gate88inter7));
  inv1  gate1745(.a(G335), .O(gate88inter8));
  nand2 gate1746(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1747(.a(s_171), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1748(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1749(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1750(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1667(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1668(.a(gate92inter0), .b(s_160), .O(gate92inter1));
  and2  gate1669(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1670(.a(s_160), .O(gate92inter3));
  inv1  gate1671(.a(s_161), .O(gate92inter4));
  nand2 gate1672(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1673(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1674(.a(G29), .O(gate92inter7));
  inv1  gate1675(.a(G341), .O(gate92inter8));
  nand2 gate1676(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1677(.a(s_161), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1678(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1679(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1680(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1121(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1122(.a(gate95inter0), .b(s_82), .O(gate95inter1));
  and2  gate1123(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1124(.a(s_82), .O(gate95inter3));
  inv1  gate1125(.a(s_83), .O(gate95inter4));
  nand2 gate1126(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1127(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1128(.a(G26), .O(gate95inter7));
  inv1  gate1129(.a(G347), .O(gate95inter8));
  nand2 gate1130(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1131(.a(s_83), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1132(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1133(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1134(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2045(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2046(.a(gate96inter0), .b(s_214), .O(gate96inter1));
  and2  gate2047(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2048(.a(s_214), .O(gate96inter3));
  inv1  gate2049(.a(s_215), .O(gate96inter4));
  nand2 gate2050(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2051(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2052(.a(G30), .O(gate96inter7));
  inv1  gate2053(.a(G347), .O(gate96inter8));
  nand2 gate2054(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2055(.a(s_215), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2056(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2057(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2058(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2185(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2186(.a(gate98inter0), .b(s_234), .O(gate98inter1));
  and2  gate2187(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2188(.a(s_234), .O(gate98inter3));
  inv1  gate2189(.a(s_235), .O(gate98inter4));
  nand2 gate2190(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2191(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2192(.a(G23), .O(gate98inter7));
  inv1  gate2193(.a(G350), .O(gate98inter8));
  nand2 gate2194(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2195(.a(s_235), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2196(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2197(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2198(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1863(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1864(.a(gate99inter0), .b(s_188), .O(gate99inter1));
  and2  gate1865(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1866(.a(s_188), .O(gate99inter3));
  inv1  gate1867(.a(s_189), .O(gate99inter4));
  nand2 gate1868(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1869(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1870(.a(G27), .O(gate99inter7));
  inv1  gate1871(.a(G353), .O(gate99inter8));
  nand2 gate1872(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1873(.a(s_189), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1874(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1875(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1876(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1485(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1486(.a(gate102inter0), .b(s_134), .O(gate102inter1));
  and2  gate1487(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1488(.a(s_134), .O(gate102inter3));
  inv1  gate1489(.a(s_135), .O(gate102inter4));
  nand2 gate1490(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1491(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1492(.a(G24), .O(gate102inter7));
  inv1  gate1493(.a(G356), .O(gate102inter8));
  nand2 gate1494(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1495(.a(s_135), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1496(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1497(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1498(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2115(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2116(.a(gate104inter0), .b(s_224), .O(gate104inter1));
  and2  gate2117(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2118(.a(s_224), .O(gate104inter3));
  inv1  gate2119(.a(s_225), .O(gate104inter4));
  nand2 gate2120(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2121(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2122(.a(G32), .O(gate104inter7));
  inv1  gate2123(.a(G359), .O(gate104inter8));
  nand2 gate2124(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2125(.a(s_225), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2126(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2127(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2128(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1499(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1500(.a(gate105inter0), .b(s_136), .O(gate105inter1));
  and2  gate1501(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1502(.a(s_136), .O(gate105inter3));
  inv1  gate1503(.a(s_137), .O(gate105inter4));
  nand2 gate1504(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1505(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1506(.a(G362), .O(gate105inter7));
  inv1  gate1507(.a(G363), .O(gate105inter8));
  nand2 gate1508(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1509(.a(s_137), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1510(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1511(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1512(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1009(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1010(.a(gate108inter0), .b(s_66), .O(gate108inter1));
  and2  gate1011(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1012(.a(s_66), .O(gate108inter3));
  inv1  gate1013(.a(s_67), .O(gate108inter4));
  nand2 gate1014(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1015(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1016(.a(G368), .O(gate108inter7));
  inv1  gate1017(.a(G369), .O(gate108inter8));
  nand2 gate1018(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1019(.a(s_67), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1020(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1021(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1022(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate883(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate884(.a(gate111inter0), .b(s_48), .O(gate111inter1));
  and2  gate885(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate886(.a(s_48), .O(gate111inter3));
  inv1  gate887(.a(s_49), .O(gate111inter4));
  nand2 gate888(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate889(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate890(.a(G374), .O(gate111inter7));
  inv1  gate891(.a(G375), .O(gate111inter8));
  nand2 gate892(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate893(.a(s_49), .b(gate111inter3), .O(gate111inter10));
  nor2  gate894(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate895(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate896(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2241(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2242(.a(gate112inter0), .b(s_242), .O(gate112inter1));
  and2  gate2243(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2244(.a(s_242), .O(gate112inter3));
  inv1  gate2245(.a(s_243), .O(gate112inter4));
  nand2 gate2246(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2247(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2248(.a(G376), .O(gate112inter7));
  inv1  gate2249(.a(G377), .O(gate112inter8));
  nand2 gate2250(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2251(.a(s_243), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2252(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2253(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2254(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1317(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1318(.a(gate113inter0), .b(s_110), .O(gate113inter1));
  and2  gate1319(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1320(.a(s_110), .O(gate113inter3));
  inv1  gate1321(.a(s_111), .O(gate113inter4));
  nand2 gate1322(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1323(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1324(.a(G378), .O(gate113inter7));
  inv1  gate1325(.a(G379), .O(gate113inter8));
  nand2 gate1326(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1327(.a(s_111), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1328(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1329(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1330(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate757(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate758(.a(gate114inter0), .b(s_30), .O(gate114inter1));
  and2  gate759(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate760(.a(s_30), .O(gate114inter3));
  inv1  gate761(.a(s_31), .O(gate114inter4));
  nand2 gate762(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate763(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate764(.a(G380), .O(gate114inter7));
  inv1  gate765(.a(G381), .O(gate114inter8));
  nand2 gate766(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate767(.a(s_31), .b(gate114inter3), .O(gate114inter10));
  nor2  gate768(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate769(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate770(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate925(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate926(.a(gate117inter0), .b(s_54), .O(gate117inter1));
  and2  gate927(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate928(.a(s_54), .O(gate117inter3));
  inv1  gate929(.a(s_55), .O(gate117inter4));
  nand2 gate930(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate931(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate932(.a(G386), .O(gate117inter7));
  inv1  gate933(.a(G387), .O(gate117inter8));
  nand2 gate934(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate935(.a(s_55), .b(gate117inter3), .O(gate117inter10));
  nor2  gate936(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate937(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate938(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1681(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1682(.a(gate120inter0), .b(s_162), .O(gate120inter1));
  and2  gate1683(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1684(.a(s_162), .O(gate120inter3));
  inv1  gate1685(.a(s_163), .O(gate120inter4));
  nand2 gate1686(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1687(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1688(.a(G392), .O(gate120inter7));
  inv1  gate1689(.a(G393), .O(gate120inter8));
  nand2 gate1690(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1691(.a(s_163), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1692(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1693(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1694(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate2269(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2270(.a(gate121inter0), .b(s_246), .O(gate121inter1));
  and2  gate2271(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2272(.a(s_246), .O(gate121inter3));
  inv1  gate2273(.a(s_247), .O(gate121inter4));
  nand2 gate2274(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2275(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2276(.a(G394), .O(gate121inter7));
  inv1  gate2277(.a(G395), .O(gate121inter8));
  nand2 gate2278(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2279(.a(s_247), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2280(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2281(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2282(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1709(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1710(.a(gate126inter0), .b(s_166), .O(gate126inter1));
  and2  gate1711(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1712(.a(s_166), .O(gate126inter3));
  inv1  gate1713(.a(s_167), .O(gate126inter4));
  nand2 gate1714(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1715(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1716(.a(G404), .O(gate126inter7));
  inv1  gate1717(.a(G405), .O(gate126inter8));
  nand2 gate1718(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1719(.a(s_167), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1720(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1721(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1722(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1303(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1304(.a(gate132inter0), .b(s_108), .O(gate132inter1));
  and2  gate1305(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1306(.a(s_108), .O(gate132inter3));
  inv1  gate1307(.a(s_109), .O(gate132inter4));
  nand2 gate1308(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1309(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1310(.a(G416), .O(gate132inter7));
  inv1  gate1311(.a(G417), .O(gate132inter8));
  nand2 gate1312(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1313(.a(s_109), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1314(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1315(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1316(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2087(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2088(.a(gate134inter0), .b(s_220), .O(gate134inter1));
  and2  gate2089(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2090(.a(s_220), .O(gate134inter3));
  inv1  gate2091(.a(s_221), .O(gate134inter4));
  nand2 gate2092(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2093(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2094(.a(G420), .O(gate134inter7));
  inv1  gate2095(.a(G421), .O(gate134inter8));
  nand2 gate2096(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2097(.a(s_221), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2098(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2099(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2100(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1975(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1976(.a(gate137inter0), .b(s_204), .O(gate137inter1));
  and2  gate1977(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1978(.a(s_204), .O(gate137inter3));
  inv1  gate1979(.a(s_205), .O(gate137inter4));
  nand2 gate1980(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1981(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1982(.a(G426), .O(gate137inter7));
  inv1  gate1983(.a(G429), .O(gate137inter8));
  nand2 gate1984(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1985(.a(s_205), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1986(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1987(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1988(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1555(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1556(.a(gate142inter0), .b(s_144), .O(gate142inter1));
  and2  gate1557(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1558(.a(s_144), .O(gate142inter3));
  inv1  gate1559(.a(s_145), .O(gate142inter4));
  nand2 gate1560(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1561(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1562(.a(G456), .O(gate142inter7));
  inv1  gate1563(.a(G459), .O(gate142inter8));
  nand2 gate1564(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1565(.a(s_145), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1566(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1567(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1568(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1429(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1430(.a(gate145inter0), .b(s_126), .O(gate145inter1));
  and2  gate1431(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1432(.a(s_126), .O(gate145inter3));
  inv1  gate1433(.a(s_127), .O(gate145inter4));
  nand2 gate1434(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1435(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1436(.a(G474), .O(gate145inter7));
  inv1  gate1437(.a(G477), .O(gate145inter8));
  nand2 gate1438(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1439(.a(s_127), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1440(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1441(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1442(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1177(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1178(.a(gate153inter0), .b(s_90), .O(gate153inter1));
  and2  gate1179(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1180(.a(s_90), .O(gate153inter3));
  inv1  gate1181(.a(s_91), .O(gate153inter4));
  nand2 gate1182(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1183(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1184(.a(G426), .O(gate153inter7));
  inv1  gate1185(.a(G522), .O(gate153inter8));
  nand2 gate1186(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1187(.a(s_91), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1188(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1189(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1190(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate967(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate968(.a(gate161inter0), .b(s_60), .O(gate161inter1));
  and2  gate969(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate970(.a(s_60), .O(gate161inter3));
  inv1  gate971(.a(s_61), .O(gate161inter4));
  nand2 gate972(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate973(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate974(.a(G450), .O(gate161inter7));
  inv1  gate975(.a(G534), .O(gate161inter8));
  nand2 gate976(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate977(.a(s_61), .b(gate161inter3), .O(gate161inter10));
  nor2  gate978(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate979(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate980(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate2101(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2102(.a(gate162inter0), .b(s_222), .O(gate162inter1));
  and2  gate2103(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2104(.a(s_222), .O(gate162inter3));
  inv1  gate2105(.a(s_223), .O(gate162inter4));
  nand2 gate2106(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2107(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2108(.a(G453), .O(gate162inter7));
  inv1  gate2109(.a(G534), .O(gate162inter8));
  nand2 gate2110(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2111(.a(s_223), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2112(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2113(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2114(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate1093(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1094(.a(gate163inter0), .b(s_78), .O(gate163inter1));
  and2  gate1095(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1096(.a(s_78), .O(gate163inter3));
  inv1  gate1097(.a(s_79), .O(gate163inter4));
  nand2 gate1098(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1099(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1100(.a(G456), .O(gate163inter7));
  inv1  gate1101(.a(G537), .O(gate163inter8));
  nand2 gate1102(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1103(.a(s_79), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1104(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1105(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1106(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2003(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2004(.a(gate167inter0), .b(s_208), .O(gate167inter1));
  and2  gate2005(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2006(.a(s_208), .O(gate167inter3));
  inv1  gate2007(.a(s_209), .O(gate167inter4));
  nand2 gate2008(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2009(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2010(.a(G468), .O(gate167inter7));
  inv1  gate2011(.a(G543), .O(gate167inter8));
  nand2 gate2012(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2013(.a(s_209), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2014(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2015(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2016(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1807(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1808(.a(gate169inter0), .b(s_180), .O(gate169inter1));
  and2  gate1809(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1810(.a(s_180), .O(gate169inter3));
  inv1  gate1811(.a(s_181), .O(gate169inter4));
  nand2 gate1812(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1813(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1814(.a(G474), .O(gate169inter7));
  inv1  gate1815(.a(G546), .O(gate169inter8));
  nand2 gate1816(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1817(.a(s_181), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1818(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1819(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1820(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1233(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1234(.a(gate172inter0), .b(s_98), .O(gate172inter1));
  and2  gate1235(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1236(.a(s_98), .O(gate172inter3));
  inv1  gate1237(.a(s_99), .O(gate172inter4));
  nand2 gate1238(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1239(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1240(.a(G483), .O(gate172inter7));
  inv1  gate1241(.a(G549), .O(gate172inter8));
  nand2 gate1242(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1243(.a(s_99), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1244(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1245(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1246(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2017(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2018(.a(gate176inter0), .b(s_210), .O(gate176inter1));
  and2  gate2019(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2020(.a(s_210), .O(gate176inter3));
  inv1  gate2021(.a(s_211), .O(gate176inter4));
  nand2 gate2022(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2023(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2024(.a(G495), .O(gate176inter7));
  inv1  gate2025(.a(G555), .O(gate176inter8));
  nand2 gate2026(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2027(.a(s_211), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2028(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2029(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2030(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1219(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1220(.a(gate183inter0), .b(s_96), .O(gate183inter1));
  and2  gate1221(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1222(.a(s_96), .O(gate183inter3));
  inv1  gate1223(.a(s_97), .O(gate183inter4));
  nand2 gate1224(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1225(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1226(.a(G516), .O(gate183inter7));
  inv1  gate1227(.a(G567), .O(gate183inter8));
  nand2 gate1228(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1229(.a(s_97), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1230(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1231(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1232(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1611(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1612(.a(gate193inter0), .b(s_152), .O(gate193inter1));
  and2  gate1613(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1614(.a(s_152), .O(gate193inter3));
  inv1  gate1615(.a(s_153), .O(gate193inter4));
  nand2 gate1616(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1617(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1618(.a(G586), .O(gate193inter7));
  inv1  gate1619(.a(G587), .O(gate193inter8));
  nand2 gate1620(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1621(.a(s_153), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1622(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1623(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1624(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1023(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1024(.a(gate195inter0), .b(s_68), .O(gate195inter1));
  and2  gate1025(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1026(.a(s_68), .O(gate195inter3));
  inv1  gate1027(.a(s_69), .O(gate195inter4));
  nand2 gate1028(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1029(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1030(.a(G590), .O(gate195inter7));
  inv1  gate1031(.a(G591), .O(gate195inter8));
  nand2 gate1032(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1033(.a(s_69), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1034(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1035(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1036(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate841(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate842(.a(gate196inter0), .b(s_42), .O(gate196inter1));
  and2  gate843(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate844(.a(s_42), .O(gate196inter3));
  inv1  gate845(.a(s_43), .O(gate196inter4));
  nand2 gate846(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate847(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate848(.a(G592), .O(gate196inter7));
  inv1  gate849(.a(G593), .O(gate196inter8));
  nand2 gate850(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate851(.a(s_43), .b(gate196inter3), .O(gate196inter10));
  nor2  gate852(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate853(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate854(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate673(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate674(.a(gate199inter0), .b(s_18), .O(gate199inter1));
  and2  gate675(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate676(.a(s_18), .O(gate199inter3));
  inv1  gate677(.a(s_19), .O(gate199inter4));
  nand2 gate678(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate679(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate680(.a(G598), .O(gate199inter7));
  inv1  gate681(.a(G599), .O(gate199inter8));
  nand2 gate682(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate683(.a(s_19), .b(gate199inter3), .O(gate199inter10));
  nor2  gate684(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate685(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate686(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1205(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1206(.a(gate205inter0), .b(s_94), .O(gate205inter1));
  and2  gate1207(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1208(.a(s_94), .O(gate205inter3));
  inv1  gate1209(.a(s_95), .O(gate205inter4));
  nand2 gate1210(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1211(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1212(.a(G622), .O(gate205inter7));
  inv1  gate1213(.a(G627), .O(gate205inter8));
  nand2 gate1214(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1215(.a(s_95), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1216(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1217(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1218(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate645(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate646(.a(gate207inter0), .b(s_14), .O(gate207inter1));
  and2  gate647(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate648(.a(s_14), .O(gate207inter3));
  inv1  gate649(.a(s_15), .O(gate207inter4));
  nand2 gate650(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate651(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate652(.a(G622), .O(gate207inter7));
  inv1  gate653(.a(G632), .O(gate207inter8));
  nand2 gate654(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate655(.a(s_15), .b(gate207inter3), .O(gate207inter10));
  nor2  gate656(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate657(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate658(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1751(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1752(.a(gate208inter0), .b(s_172), .O(gate208inter1));
  and2  gate1753(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1754(.a(s_172), .O(gate208inter3));
  inv1  gate1755(.a(s_173), .O(gate208inter4));
  nand2 gate1756(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1757(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1758(.a(G627), .O(gate208inter7));
  inv1  gate1759(.a(G637), .O(gate208inter8));
  nand2 gate1760(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1761(.a(s_173), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1762(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1763(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1764(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1359(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1360(.a(gate211inter0), .b(s_116), .O(gate211inter1));
  and2  gate1361(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1362(.a(s_116), .O(gate211inter3));
  inv1  gate1363(.a(s_117), .O(gate211inter4));
  nand2 gate1364(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1365(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1366(.a(G612), .O(gate211inter7));
  inv1  gate1367(.a(G669), .O(gate211inter8));
  nand2 gate1368(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1369(.a(s_117), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1370(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1371(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1372(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1163(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1164(.a(gate216inter0), .b(s_88), .O(gate216inter1));
  and2  gate1165(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1166(.a(s_88), .O(gate216inter3));
  inv1  gate1167(.a(s_89), .O(gate216inter4));
  nand2 gate1168(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1169(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1170(.a(G617), .O(gate216inter7));
  inv1  gate1171(.a(G675), .O(gate216inter8));
  nand2 gate1172(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1173(.a(s_89), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1174(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1175(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1176(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2199(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2200(.a(gate217inter0), .b(s_236), .O(gate217inter1));
  and2  gate2201(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2202(.a(s_236), .O(gate217inter3));
  inv1  gate2203(.a(s_237), .O(gate217inter4));
  nand2 gate2204(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2205(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2206(.a(G622), .O(gate217inter7));
  inv1  gate2207(.a(G678), .O(gate217inter8));
  nand2 gate2208(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2209(.a(s_237), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2210(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2211(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2212(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1331(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1332(.a(gate218inter0), .b(s_112), .O(gate218inter1));
  and2  gate1333(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1334(.a(s_112), .O(gate218inter3));
  inv1  gate1335(.a(s_113), .O(gate218inter4));
  nand2 gate1336(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1337(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1338(.a(G627), .O(gate218inter7));
  inv1  gate1339(.a(G678), .O(gate218inter8));
  nand2 gate1340(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1341(.a(s_113), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1342(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1343(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1344(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate575(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate576(.a(gate219inter0), .b(s_4), .O(gate219inter1));
  and2  gate577(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate578(.a(s_4), .O(gate219inter3));
  inv1  gate579(.a(s_5), .O(gate219inter4));
  nand2 gate580(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate581(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate582(.a(G632), .O(gate219inter7));
  inv1  gate583(.a(G681), .O(gate219inter8));
  nand2 gate584(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate585(.a(s_5), .b(gate219inter3), .O(gate219inter10));
  nor2  gate586(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate587(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate588(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1191(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1192(.a(gate222inter0), .b(s_92), .O(gate222inter1));
  and2  gate1193(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1194(.a(s_92), .O(gate222inter3));
  inv1  gate1195(.a(s_93), .O(gate222inter4));
  nand2 gate1196(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1197(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1198(.a(G632), .O(gate222inter7));
  inv1  gate1199(.a(G684), .O(gate222inter8));
  nand2 gate1200(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1201(.a(s_93), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1202(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1203(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1204(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate701(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate702(.a(gate240inter0), .b(s_22), .O(gate240inter1));
  and2  gate703(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate704(.a(s_22), .O(gate240inter3));
  inv1  gate705(.a(s_23), .O(gate240inter4));
  nand2 gate706(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate707(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate708(.a(G263), .O(gate240inter7));
  inv1  gate709(.a(G715), .O(gate240inter8));
  nand2 gate710(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate711(.a(s_23), .b(gate240inter3), .O(gate240inter10));
  nor2  gate712(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate713(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate714(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2255(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2256(.a(gate242inter0), .b(s_244), .O(gate242inter1));
  and2  gate2257(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2258(.a(s_244), .O(gate242inter3));
  inv1  gate2259(.a(s_245), .O(gate242inter4));
  nand2 gate2260(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2261(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2262(.a(G718), .O(gate242inter7));
  inv1  gate2263(.a(G730), .O(gate242inter8));
  nand2 gate2264(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2265(.a(s_245), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2266(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2267(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2268(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2213(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2214(.a(gate249inter0), .b(s_238), .O(gate249inter1));
  and2  gate2215(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2216(.a(s_238), .O(gate249inter3));
  inv1  gate2217(.a(s_239), .O(gate249inter4));
  nand2 gate2218(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2219(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2220(.a(G254), .O(gate249inter7));
  inv1  gate2221(.a(G742), .O(gate249inter8));
  nand2 gate2222(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2223(.a(s_239), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2224(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2225(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2226(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate981(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate982(.a(gate251inter0), .b(s_62), .O(gate251inter1));
  and2  gate983(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate984(.a(s_62), .O(gate251inter3));
  inv1  gate985(.a(s_63), .O(gate251inter4));
  nand2 gate986(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate987(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate988(.a(G257), .O(gate251inter7));
  inv1  gate989(.a(G745), .O(gate251inter8));
  nand2 gate990(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate991(.a(s_63), .b(gate251inter3), .O(gate251inter10));
  nor2  gate992(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate993(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate994(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1723(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1724(.a(gate255inter0), .b(s_168), .O(gate255inter1));
  and2  gate1725(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1726(.a(s_168), .O(gate255inter3));
  inv1  gate1727(.a(s_169), .O(gate255inter4));
  nand2 gate1728(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1729(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1730(.a(G263), .O(gate255inter7));
  inv1  gate1731(.a(G751), .O(gate255inter8));
  nand2 gate1732(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1733(.a(s_169), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1734(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1735(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1736(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate897(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate898(.a(gate256inter0), .b(s_50), .O(gate256inter1));
  and2  gate899(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate900(.a(s_50), .O(gate256inter3));
  inv1  gate901(.a(s_51), .O(gate256inter4));
  nand2 gate902(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate903(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate904(.a(G715), .O(gate256inter7));
  inv1  gate905(.a(G751), .O(gate256inter8));
  nand2 gate906(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate907(.a(s_51), .b(gate256inter3), .O(gate256inter10));
  nor2  gate908(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate909(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate910(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2143(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2144(.a(gate258inter0), .b(s_228), .O(gate258inter1));
  and2  gate2145(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2146(.a(s_228), .O(gate258inter3));
  inv1  gate2147(.a(s_229), .O(gate258inter4));
  nand2 gate2148(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2149(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2150(.a(G756), .O(gate258inter7));
  inv1  gate2151(.a(G757), .O(gate258inter8));
  nand2 gate2152(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2153(.a(s_229), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2154(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2155(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2156(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1625(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1626(.a(gate259inter0), .b(s_154), .O(gate259inter1));
  and2  gate1627(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1628(.a(s_154), .O(gate259inter3));
  inv1  gate1629(.a(s_155), .O(gate259inter4));
  nand2 gate1630(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1631(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1632(.a(G758), .O(gate259inter7));
  inv1  gate1633(.a(G759), .O(gate259inter8));
  nand2 gate1634(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1635(.a(s_155), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1636(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1637(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1638(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1051(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1052(.a(gate260inter0), .b(s_72), .O(gate260inter1));
  and2  gate1053(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1054(.a(s_72), .O(gate260inter3));
  inv1  gate1055(.a(s_73), .O(gate260inter4));
  nand2 gate1056(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1057(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1058(.a(G760), .O(gate260inter7));
  inv1  gate1059(.a(G761), .O(gate260inter8));
  nand2 gate1060(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1061(.a(s_73), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1062(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1063(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1064(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate603(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate604(.a(gate266inter0), .b(s_8), .O(gate266inter1));
  and2  gate605(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate606(.a(s_8), .O(gate266inter3));
  inv1  gate607(.a(s_9), .O(gate266inter4));
  nand2 gate608(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate609(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate610(.a(G645), .O(gate266inter7));
  inv1  gate611(.a(G773), .O(gate266inter8));
  nand2 gate612(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate613(.a(s_9), .b(gate266inter3), .O(gate266inter10));
  nor2  gate614(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate615(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate616(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1905(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1906(.a(gate273inter0), .b(s_194), .O(gate273inter1));
  and2  gate1907(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1908(.a(s_194), .O(gate273inter3));
  inv1  gate1909(.a(s_195), .O(gate273inter4));
  nand2 gate1910(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1911(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1912(.a(G642), .O(gate273inter7));
  inv1  gate1913(.a(G794), .O(gate273inter8));
  nand2 gate1914(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1915(.a(s_195), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1916(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1917(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1918(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate547(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate548(.a(gate274inter0), .b(s_0), .O(gate274inter1));
  and2  gate549(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate550(.a(s_0), .O(gate274inter3));
  inv1  gate551(.a(s_1), .O(gate274inter4));
  nand2 gate552(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate553(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate554(.a(G770), .O(gate274inter7));
  inv1  gate555(.a(G794), .O(gate274inter8));
  nand2 gate556(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate557(.a(s_1), .b(gate274inter3), .O(gate274inter10));
  nor2  gate558(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate559(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate560(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1947(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1948(.a(gate276inter0), .b(s_200), .O(gate276inter1));
  and2  gate1949(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1950(.a(s_200), .O(gate276inter3));
  inv1  gate1951(.a(s_201), .O(gate276inter4));
  nand2 gate1952(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1953(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1954(.a(G773), .O(gate276inter7));
  inv1  gate1955(.a(G797), .O(gate276inter8));
  nand2 gate1956(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1957(.a(s_201), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1958(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1959(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1960(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1107(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1108(.a(gate283inter0), .b(s_80), .O(gate283inter1));
  and2  gate1109(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1110(.a(s_80), .O(gate283inter3));
  inv1  gate1111(.a(s_81), .O(gate283inter4));
  nand2 gate1112(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1113(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1114(.a(G657), .O(gate283inter7));
  inv1  gate1115(.a(G809), .O(gate283inter8));
  nand2 gate1116(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1117(.a(s_81), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1118(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1119(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1120(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1821(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1822(.a(gate287inter0), .b(s_182), .O(gate287inter1));
  and2  gate1823(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1824(.a(s_182), .O(gate287inter3));
  inv1  gate1825(.a(s_183), .O(gate287inter4));
  nand2 gate1826(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1827(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1828(.a(G663), .O(gate287inter7));
  inv1  gate1829(.a(G815), .O(gate287inter8));
  nand2 gate1830(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1831(.a(s_183), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1832(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1833(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1834(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1541(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1542(.a(gate387inter0), .b(s_142), .O(gate387inter1));
  and2  gate1543(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1544(.a(s_142), .O(gate387inter3));
  inv1  gate1545(.a(s_143), .O(gate387inter4));
  nand2 gate1546(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1547(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1548(.a(G1), .O(gate387inter7));
  inv1  gate1549(.a(G1036), .O(gate387inter8));
  nand2 gate1550(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1551(.a(s_143), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1552(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1553(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1554(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1933(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1934(.a(gate388inter0), .b(s_198), .O(gate388inter1));
  and2  gate1935(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1936(.a(s_198), .O(gate388inter3));
  inv1  gate1937(.a(s_199), .O(gate388inter4));
  nand2 gate1938(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1939(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1940(.a(G2), .O(gate388inter7));
  inv1  gate1941(.a(G1039), .O(gate388inter8));
  nand2 gate1942(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1943(.a(s_199), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1944(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1945(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1946(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1989(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1990(.a(gate395inter0), .b(s_206), .O(gate395inter1));
  and2  gate1991(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1992(.a(s_206), .O(gate395inter3));
  inv1  gate1993(.a(s_207), .O(gate395inter4));
  nand2 gate1994(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1995(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1996(.a(G9), .O(gate395inter7));
  inv1  gate1997(.a(G1060), .O(gate395inter8));
  nand2 gate1998(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1999(.a(s_207), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2000(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2001(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2002(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1149(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1150(.a(gate400inter0), .b(s_86), .O(gate400inter1));
  and2  gate1151(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1152(.a(s_86), .O(gate400inter3));
  inv1  gate1153(.a(s_87), .O(gate400inter4));
  nand2 gate1154(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1155(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1156(.a(G14), .O(gate400inter7));
  inv1  gate1157(.a(G1075), .O(gate400inter8));
  nand2 gate1158(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1159(.a(s_87), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1160(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1161(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1162(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate939(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate940(.a(gate402inter0), .b(s_56), .O(gate402inter1));
  and2  gate941(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate942(.a(s_56), .O(gate402inter3));
  inv1  gate943(.a(s_57), .O(gate402inter4));
  nand2 gate944(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate945(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate946(.a(G16), .O(gate402inter7));
  inv1  gate947(.a(G1081), .O(gate402inter8));
  nand2 gate948(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate949(.a(s_57), .b(gate402inter3), .O(gate402inter10));
  nor2  gate950(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate951(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate952(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1793(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1794(.a(gate403inter0), .b(s_178), .O(gate403inter1));
  and2  gate1795(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1796(.a(s_178), .O(gate403inter3));
  inv1  gate1797(.a(s_179), .O(gate403inter4));
  nand2 gate1798(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1799(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1800(.a(G17), .O(gate403inter7));
  inv1  gate1801(.a(G1084), .O(gate403inter8));
  nand2 gate1802(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1803(.a(s_179), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1804(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1805(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1806(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate561(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate562(.a(gate404inter0), .b(s_2), .O(gate404inter1));
  and2  gate563(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate564(.a(s_2), .O(gate404inter3));
  inv1  gate565(.a(s_3), .O(gate404inter4));
  nand2 gate566(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate567(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate568(.a(G18), .O(gate404inter7));
  inv1  gate569(.a(G1087), .O(gate404inter8));
  nand2 gate570(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate571(.a(s_3), .b(gate404inter3), .O(gate404inter10));
  nor2  gate572(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate573(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate574(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2283(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2284(.a(gate406inter0), .b(s_248), .O(gate406inter1));
  and2  gate2285(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2286(.a(s_248), .O(gate406inter3));
  inv1  gate2287(.a(s_249), .O(gate406inter4));
  nand2 gate2288(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2289(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2290(.a(G20), .O(gate406inter7));
  inv1  gate2291(.a(G1093), .O(gate406inter8));
  nand2 gate2292(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2293(.a(s_249), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2294(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2295(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2296(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1569(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1570(.a(gate409inter0), .b(s_146), .O(gate409inter1));
  and2  gate1571(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1572(.a(s_146), .O(gate409inter3));
  inv1  gate1573(.a(s_147), .O(gate409inter4));
  nand2 gate1574(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1575(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1576(.a(G23), .O(gate409inter7));
  inv1  gate1577(.a(G1102), .O(gate409inter8));
  nand2 gate1578(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1579(.a(s_147), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1580(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1581(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1582(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2171(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2172(.a(gate411inter0), .b(s_232), .O(gate411inter1));
  and2  gate2173(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2174(.a(s_232), .O(gate411inter3));
  inv1  gate2175(.a(s_233), .O(gate411inter4));
  nand2 gate2176(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2177(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2178(.a(G25), .O(gate411inter7));
  inv1  gate2179(.a(G1108), .O(gate411inter8));
  nand2 gate2180(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2181(.a(s_233), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2182(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2183(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2184(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1513(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1514(.a(gate412inter0), .b(s_138), .O(gate412inter1));
  and2  gate1515(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1516(.a(s_138), .O(gate412inter3));
  inv1  gate1517(.a(s_139), .O(gate412inter4));
  nand2 gate1518(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1519(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1520(.a(G26), .O(gate412inter7));
  inv1  gate1521(.a(G1111), .O(gate412inter8));
  nand2 gate1522(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1523(.a(s_139), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1524(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1525(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1526(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1289(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1290(.a(gate415inter0), .b(s_106), .O(gate415inter1));
  and2  gate1291(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1292(.a(s_106), .O(gate415inter3));
  inv1  gate1293(.a(s_107), .O(gate415inter4));
  nand2 gate1294(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1295(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1296(.a(G29), .O(gate415inter7));
  inv1  gate1297(.a(G1120), .O(gate415inter8));
  nand2 gate1298(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1299(.a(s_107), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1300(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1301(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1302(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1583(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1584(.a(gate417inter0), .b(s_148), .O(gate417inter1));
  and2  gate1585(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1586(.a(s_148), .O(gate417inter3));
  inv1  gate1587(.a(s_149), .O(gate417inter4));
  nand2 gate1588(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1589(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1590(.a(G31), .O(gate417inter7));
  inv1  gate1591(.a(G1126), .O(gate417inter8));
  nand2 gate1592(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1593(.a(s_149), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1594(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1595(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1596(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1387(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1388(.a(gate418inter0), .b(s_120), .O(gate418inter1));
  and2  gate1389(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1390(.a(s_120), .O(gate418inter3));
  inv1  gate1391(.a(s_121), .O(gate418inter4));
  nand2 gate1392(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1393(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1394(.a(G32), .O(gate418inter7));
  inv1  gate1395(.a(G1129), .O(gate418inter8));
  nand2 gate1396(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1397(.a(s_121), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1398(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1399(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1400(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1373(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1374(.a(gate420inter0), .b(s_118), .O(gate420inter1));
  and2  gate1375(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1376(.a(s_118), .O(gate420inter3));
  inv1  gate1377(.a(s_119), .O(gate420inter4));
  nand2 gate1378(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1379(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1380(.a(G1036), .O(gate420inter7));
  inv1  gate1381(.a(G1132), .O(gate420inter8));
  nand2 gate1382(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1383(.a(s_119), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1384(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1385(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1386(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1765(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1766(.a(gate422inter0), .b(s_174), .O(gate422inter1));
  and2  gate1767(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1768(.a(s_174), .O(gate422inter3));
  inv1  gate1769(.a(s_175), .O(gate422inter4));
  nand2 gate1770(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1771(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1772(.a(G1039), .O(gate422inter7));
  inv1  gate1773(.a(G1135), .O(gate422inter8));
  nand2 gate1774(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1775(.a(s_175), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1776(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1777(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1778(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1877(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1878(.a(gate429inter0), .b(s_190), .O(gate429inter1));
  and2  gate1879(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1880(.a(s_190), .O(gate429inter3));
  inv1  gate1881(.a(s_191), .O(gate429inter4));
  nand2 gate1882(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1883(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1884(.a(G6), .O(gate429inter7));
  inv1  gate1885(.a(G1147), .O(gate429inter8));
  nand2 gate1886(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1887(.a(s_191), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1888(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1889(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1890(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1079(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1080(.a(gate431inter0), .b(s_76), .O(gate431inter1));
  and2  gate1081(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1082(.a(s_76), .O(gate431inter3));
  inv1  gate1083(.a(s_77), .O(gate431inter4));
  nand2 gate1084(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1085(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1086(.a(G7), .O(gate431inter7));
  inv1  gate1087(.a(G1150), .O(gate431inter8));
  nand2 gate1088(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1089(.a(s_77), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1090(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1091(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1092(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1247(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1248(.a(gate432inter0), .b(s_100), .O(gate432inter1));
  and2  gate1249(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1250(.a(s_100), .O(gate432inter3));
  inv1  gate1251(.a(s_101), .O(gate432inter4));
  nand2 gate1252(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1253(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1254(.a(G1054), .O(gate432inter7));
  inv1  gate1255(.a(G1150), .O(gate432inter8));
  nand2 gate1256(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1257(.a(s_101), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1258(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1259(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1260(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2129(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2130(.a(gate433inter0), .b(s_226), .O(gate433inter1));
  and2  gate2131(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2132(.a(s_226), .O(gate433inter3));
  inv1  gate2133(.a(s_227), .O(gate433inter4));
  nand2 gate2134(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2135(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2136(.a(G8), .O(gate433inter7));
  inv1  gate2137(.a(G1153), .O(gate433inter8));
  nand2 gate2138(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2139(.a(s_227), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2140(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2141(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2142(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1275(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1276(.a(gate437inter0), .b(s_104), .O(gate437inter1));
  and2  gate1277(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1278(.a(s_104), .O(gate437inter3));
  inv1  gate1279(.a(s_105), .O(gate437inter4));
  nand2 gate1280(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1281(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1282(.a(G10), .O(gate437inter7));
  inv1  gate1283(.a(G1159), .O(gate437inter8));
  nand2 gate1284(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1285(.a(s_105), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1286(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1287(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1288(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate855(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate856(.a(gate438inter0), .b(s_44), .O(gate438inter1));
  and2  gate857(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate858(.a(s_44), .O(gate438inter3));
  inv1  gate859(.a(s_45), .O(gate438inter4));
  nand2 gate860(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate861(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate862(.a(G1063), .O(gate438inter7));
  inv1  gate863(.a(G1159), .O(gate438inter8));
  nand2 gate864(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate865(.a(s_45), .b(gate438inter3), .O(gate438inter10));
  nor2  gate866(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate867(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate868(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2297(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2298(.a(gate440inter0), .b(s_250), .O(gate440inter1));
  and2  gate2299(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2300(.a(s_250), .O(gate440inter3));
  inv1  gate2301(.a(s_251), .O(gate440inter4));
  nand2 gate2302(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2303(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2304(.a(G1066), .O(gate440inter7));
  inv1  gate2305(.a(G1162), .O(gate440inter8));
  nand2 gate2306(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2307(.a(s_251), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2308(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2309(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2310(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate743(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate744(.a(gate444inter0), .b(s_28), .O(gate444inter1));
  and2  gate745(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate746(.a(s_28), .O(gate444inter3));
  inv1  gate747(.a(s_29), .O(gate444inter4));
  nand2 gate748(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate749(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate750(.a(G1072), .O(gate444inter7));
  inv1  gate751(.a(G1168), .O(gate444inter8));
  nand2 gate752(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate753(.a(s_29), .b(gate444inter3), .O(gate444inter10));
  nor2  gate754(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate755(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate756(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate953(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate954(.a(gate445inter0), .b(s_58), .O(gate445inter1));
  and2  gate955(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate956(.a(s_58), .O(gate445inter3));
  inv1  gate957(.a(s_59), .O(gate445inter4));
  nand2 gate958(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate959(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate960(.a(G14), .O(gate445inter7));
  inv1  gate961(.a(G1171), .O(gate445inter8));
  nand2 gate962(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate963(.a(s_59), .b(gate445inter3), .O(gate445inter10));
  nor2  gate964(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate965(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate966(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1695(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1696(.a(gate446inter0), .b(s_164), .O(gate446inter1));
  and2  gate1697(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1698(.a(s_164), .O(gate446inter3));
  inv1  gate1699(.a(s_165), .O(gate446inter4));
  nand2 gate1700(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1701(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1702(.a(G1075), .O(gate446inter7));
  inv1  gate1703(.a(G1171), .O(gate446inter8));
  nand2 gate1704(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1705(.a(s_165), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1706(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1707(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1708(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1527(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1528(.a(gate448inter0), .b(s_140), .O(gate448inter1));
  and2  gate1529(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1530(.a(s_140), .O(gate448inter3));
  inv1  gate1531(.a(s_141), .O(gate448inter4));
  nand2 gate1532(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1533(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1534(.a(G1078), .O(gate448inter7));
  inv1  gate1535(.a(G1174), .O(gate448inter8));
  nand2 gate1536(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1537(.a(s_141), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1538(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1539(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1540(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2031(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2032(.a(gate449inter0), .b(s_212), .O(gate449inter1));
  and2  gate2033(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2034(.a(s_212), .O(gate449inter3));
  inv1  gate2035(.a(s_213), .O(gate449inter4));
  nand2 gate2036(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2037(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2038(.a(G16), .O(gate449inter7));
  inv1  gate2039(.a(G1177), .O(gate449inter8));
  nand2 gate2040(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2041(.a(s_213), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2042(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2043(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2044(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate869(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate870(.a(gate453inter0), .b(s_46), .O(gate453inter1));
  and2  gate871(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate872(.a(s_46), .O(gate453inter3));
  inv1  gate873(.a(s_47), .O(gate453inter4));
  nand2 gate874(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate875(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate876(.a(G18), .O(gate453inter7));
  inv1  gate877(.a(G1183), .O(gate453inter8));
  nand2 gate878(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate879(.a(s_47), .b(gate453inter3), .O(gate453inter10));
  nor2  gate880(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate881(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate882(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1919(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1920(.a(gate462inter0), .b(s_196), .O(gate462inter1));
  and2  gate1921(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1922(.a(s_196), .O(gate462inter3));
  inv1  gate1923(.a(s_197), .O(gate462inter4));
  nand2 gate1924(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1925(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1926(.a(G1099), .O(gate462inter7));
  inv1  gate1927(.a(G1195), .O(gate462inter8));
  nand2 gate1928(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1929(.a(s_197), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1930(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1931(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1932(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1597(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1598(.a(gate467inter0), .b(s_150), .O(gate467inter1));
  and2  gate1599(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1600(.a(s_150), .O(gate467inter3));
  inv1  gate1601(.a(s_151), .O(gate467inter4));
  nand2 gate1602(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1603(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1604(.a(G25), .O(gate467inter7));
  inv1  gate1605(.a(G1204), .O(gate467inter8));
  nand2 gate1606(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1607(.a(s_151), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1608(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1609(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1610(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1961(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1962(.a(gate468inter0), .b(s_202), .O(gate468inter1));
  and2  gate1963(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1964(.a(s_202), .O(gate468inter3));
  inv1  gate1965(.a(s_203), .O(gate468inter4));
  nand2 gate1966(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1967(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1968(.a(G1108), .O(gate468inter7));
  inv1  gate1969(.a(G1204), .O(gate468inter8));
  nand2 gate1970(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1971(.a(s_203), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1972(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1973(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1974(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1065(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1066(.a(gate473inter0), .b(s_74), .O(gate473inter1));
  and2  gate1067(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1068(.a(s_74), .O(gate473inter3));
  inv1  gate1069(.a(s_75), .O(gate473inter4));
  nand2 gate1070(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1071(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1072(.a(G28), .O(gate473inter7));
  inv1  gate1073(.a(G1213), .O(gate473inter8));
  nand2 gate1074(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1075(.a(s_75), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1076(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1077(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1078(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2059(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2060(.a(gate474inter0), .b(s_216), .O(gate474inter1));
  and2  gate2061(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2062(.a(s_216), .O(gate474inter3));
  inv1  gate2063(.a(s_217), .O(gate474inter4));
  nand2 gate2064(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2065(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2066(.a(G1117), .O(gate474inter7));
  inv1  gate2067(.a(G1213), .O(gate474inter8));
  nand2 gate2068(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2069(.a(s_217), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2070(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2071(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2072(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1471(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1472(.a(gate477inter0), .b(s_132), .O(gate477inter1));
  and2  gate1473(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1474(.a(s_132), .O(gate477inter3));
  inv1  gate1475(.a(s_133), .O(gate477inter4));
  nand2 gate1476(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1477(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1478(.a(G30), .O(gate477inter7));
  inv1  gate1479(.a(G1219), .O(gate477inter8));
  nand2 gate1480(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1481(.a(s_133), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1482(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1483(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1484(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1037(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1038(.a(gate482inter0), .b(s_70), .O(gate482inter1));
  and2  gate1039(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1040(.a(s_70), .O(gate482inter3));
  inv1  gate1041(.a(s_71), .O(gate482inter4));
  nand2 gate1042(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1043(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1044(.a(G1129), .O(gate482inter7));
  inv1  gate1045(.a(G1225), .O(gate482inter8));
  nand2 gate1046(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1047(.a(s_71), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1048(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1049(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1050(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate589(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate590(.a(gate484inter0), .b(s_6), .O(gate484inter1));
  and2  gate591(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate592(.a(s_6), .O(gate484inter3));
  inv1  gate593(.a(s_7), .O(gate484inter4));
  nand2 gate594(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate595(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate596(.a(G1230), .O(gate484inter7));
  inv1  gate597(.a(G1231), .O(gate484inter8));
  nand2 gate598(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate599(.a(s_7), .b(gate484inter3), .O(gate484inter10));
  nor2  gate600(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate601(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate602(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate715(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate716(.a(gate488inter0), .b(s_24), .O(gate488inter1));
  and2  gate717(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate718(.a(s_24), .O(gate488inter3));
  inv1  gate719(.a(s_25), .O(gate488inter4));
  nand2 gate720(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate721(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate722(.a(G1238), .O(gate488inter7));
  inv1  gate723(.a(G1239), .O(gate488inter8));
  nand2 gate724(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate725(.a(s_25), .b(gate488inter3), .O(gate488inter10));
  nor2  gate726(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate727(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate728(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1891(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1892(.a(gate490inter0), .b(s_192), .O(gate490inter1));
  and2  gate1893(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1894(.a(s_192), .O(gate490inter3));
  inv1  gate1895(.a(s_193), .O(gate490inter4));
  nand2 gate1896(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1897(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1898(.a(G1242), .O(gate490inter7));
  inv1  gate1899(.a(G1243), .O(gate490inter8));
  nand2 gate1900(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1901(.a(s_193), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1902(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1903(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1904(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate687(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate688(.a(gate505inter0), .b(s_20), .O(gate505inter1));
  and2  gate689(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate690(.a(s_20), .O(gate505inter3));
  inv1  gate691(.a(s_21), .O(gate505inter4));
  nand2 gate692(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate693(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate694(.a(G1272), .O(gate505inter7));
  inv1  gate695(.a(G1273), .O(gate505inter8));
  nand2 gate696(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate697(.a(s_21), .b(gate505inter3), .O(gate505inter10));
  nor2  gate698(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate699(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate700(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1849(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1850(.a(gate507inter0), .b(s_186), .O(gate507inter1));
  and2  gate1851(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1852(.a(s_186), .O(gate507inter3));
  inv1  gate1853(.a(s_187), .O(gate507inter4));
  nand2 gate1854(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1855(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1856(.a(G1276), .O(gate507inter7));
  inv1  gate1857(.a(G1277), .O(gate507inter8));
  nand2 gate1858(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1859(.a(s_187), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1860(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1861(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1862(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate617(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate618(.a(gate508inter0), .b(s_10), .O(gate508inter1));
  and2  gate619(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate620(.a(s_10), .O(gate508inter3));
  inv1  gate621(.a(s_11), .O(gate508inter4));
  nand2 gate622(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate623(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate624(.a(G1278), .O(gate508inter7));
  inv1  gate625(.a(G1279), .O(gate508inter8));
  nand2 gate626(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate627(.a(s_11), .b(gate508inter3), .O(gate508inter10));
  nor2  gate628(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate629(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate630(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate799(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate800(.a(gate511inter0), .b(s_36), .O(gate511inter1));
  and2  gate801(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate802(.a(s_36), .O(gate511inter3));
  inv1  gate803(.a(s_37), .O(gate511inter4));
  nand2 gate804(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate805(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate806(.a(G1284), .O(gate511inter7));
  inv1  gate807(.a(G1285), .O(gate511inter8));
  nand2 gate808(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate809(.a(s_37), .b(gate511inter3), .O(gate511inter10));
  nor2  gate810(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate811(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate812(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate631(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate632(.a(gate512inter0), .b(s_12), .O(gate512inter1));
  and2  gate633(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate634(.a(s_12), .O(gate512inter3));
  inv1  gate635(.a(s_13), .O(gate512inter4));
  nand2 gate636(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate637(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate638(.a(G1286), .O(gate512inter7));
  inv1  gate639(.a(G1287), .O(gate512inter8));
  nand2 gate640(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate641(.a(s_13), .b(gate512inter3), .O(gate512inter10));
  nor2  gate642(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate643(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate644(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule