module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate217(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate218(.a(gate4inter0), .b(s_2), .O(gate4inter1));
  and2  gate219(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate220(.a(s_2), .O(gate4inter3));
  inv1  gate221(.a(s_3), .O(gate4inter4));
  nand2 gate222(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate223(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate224(.a(N25), .O(gate4inter7));
  inv1  gate225(.a(N29), .O(gate4inter8));
  nand2 gate226(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate227(.a(s_3), .b(gate4inter3), .O(gate4inter10));
  nor2  gate228(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate229(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate230(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate203(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate204(.a(gate8inter0), .b(s_0), .O(gate8inter1));
  and2  gate205(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate206(.a(s_0), .O(gate8inter3));
  inv1  gate207(.a(s_1), .O(gate8inter4));
  nand2 gate208(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate209(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate210(.a(N57), .O(gate8inter7));
  inv1  gate211(.a(N61), .O(gate8inter8));
  nand2 gate212(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate213(.a(s_1), .b(gate8inter3), .O(gate8inter10));
  nor2  gate214(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate215(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate216(.a(gate8inter12), .b(gate8inter1), .O(N257));

  xor2  gate315(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate316(.a(gate9inter0), .b(s_16), .O(gate9inter1));
  and2  gate317(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate318(.a(s_16), .O(gate9inter3));
  inv1  gate319(.a(s_17), .O(gate9inter4));
  nand2 gate320(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate321(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate322(.a(N65), .O(gate9inter7));
  inv1  gate323(.a(N69), .O(gate9inter8));
  nand2 gate324(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate325(.a(s_17), .b(gate9inter3), .O(gate9inter10));
  nor2  gate326(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate327(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate328(.a(gate9inter12), .b(gate9inter1), .O(N258));
xor2 gate10( .a(N73), .b(N77), .O(N259) );

  xor2  gate343(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate344(.a(gate11inter0), .b(s_20), .O(gate11inter1));
  and2  gate345(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate346(.a(s_20), .O(gate11inter3));
  inv1  gate347(.a(s_21), .O(gate11inter4));
  nand2 gate348(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate349(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate350(.a(N81), .O(gate11inter7));
  inv1  gate351(.a(N85), .O(gate11inter8));
  nand2 gate352(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate353(.a(s_21), .b(gate11inter3), .O(gate11inter10));
  nor2  gate354(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate355(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate356(.a(gate11inter12), .b(gate11inter1), .O(N260));
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );

  xor2  gate329(.a(N21), .b(N5), .O(gate27inter0));
  nand2 gate330(.a(gate27inter0), .b(s_18), .O(gate27inter1));
  and2  gate331(.a(N21), .b(N5), .O(gate27inter2));
  inv1  gate332(.a(s_18), .O(gate27inter3));
  inv1  gate333(.a(s_19), .O(gate27inter4));
  nand2 gate334(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate335(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate336(.a(N5), .O(gate27inter7));
  inv1  gate337(.a(N21), .O(gate27inter8));
  nand2 gate338(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate339(.a(s_19), .b(gate27inter3), .O(gate27inter10));
  nor2  gate340(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate341(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate342(.a(gate27inter12), .b(gate27inter1), .O(N276));
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate245(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate246(.a(gate30inter0), .b(s_6), .O(gate30inter1));
  and2  gate247(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate248(.a(s_6), .O(gate30inter3));
  inv1  gate249(.a(s_7), .O(gate30inter4));
  nand2 gate250(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate251(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate252(.a(N41), .O(gate30inter7));
  inv1  gate253(.a(N57), .O(gate30inter8));
  nand2 gate254(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate255(.a(s_7), .b(gate30inter3), .O(gate30inter10));
  nor2  gate256(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate257(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate258(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );

  xor2  gate385(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate386(.a(gate34inter0), .b(s_26), .O(gate34inter1));
  and2  gate387(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate388(.a(s_26), .O(gate34inter3));
  inv1  gate389(.a(s_27), .O(gate34inter4));
  nand2 gate390(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate391(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate392(.a(N97), .O(gate34inter7));
  inv1  gate393(.a(N113), .O(gate34inter8));
  nand2 gate394(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate395(.a(s_27), .b(gate34inter3), .O(gate34inter10));
  nor2  gate396(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate397(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate398(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate399(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate400(.a(gate50inter0), .b(s_28), .O(gate50inter1));
  and2  gate401(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate402(.a(s_28), .O(gate50inter3));
  inv1  gate403(.a(s_29), .O(gate50inter4));
  nand2 gate404(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate405(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate406(.a(N276), .O(gate50inter7));
  inv1  gate407(.a(N277), .O(gate50inter8));
  nand2 gate408(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate409(.a(s_29), .b(gate50inter3), .O(gate50inter10));
  nor2  gate410(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate411(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate412(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );

  xor2  gate273(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate274(.a(gate58inter0), .b(s_10), .O(gate58inter1));
  and2  gate275(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate276(.a(s_10), .O(gate58inter3));
  inv1  gate277(.a(s_11), .O(gate58inter4));
  nand2 gate278(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate279(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate280(.a(N296), .O(gate58inter7));
  inv1  gate281(.a(N299), .O(gate58inter8));
  nand2 gate282(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate283(.a(s_11), .b(gate58inter3), .O(gate58inter10));
  nor2  gate284(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate285(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate286(.a(gate58inter12), .b(gate58inter1), .O(N339));
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );

  xor2  gate259(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate260(.a(gate64inter0), .b(s_8), .O(gate64inter1));
  and2  gate261(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate262(.a(s_8), .O(gate64inter3));
  inv1  gate263(.a(s_9), .O(gate64inter4));
  nand2 gate264(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate265(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate266(.a(N305), .O(gate64inter7));
  inv1  gate267(.a(N311), .O(gate64inter8));
  nand2 gate268(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate269(.a(s_9), .b(gate64inter3), .O(gate64inter10));
  nor2  gate270(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate271(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate272(.a(gate64inter12), .b(gate64inter1), .O(N345));
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate231(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate232(.a(gate70inter0), .b(s_4), .O(gate70inter1));
  and2  gate233(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate234(.a(s_4), .O(gate70inter3));
  inv1  gate235(.a(s_5), .O(gate70inter4));
  nand2 gate236(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate237(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate238(.a(N271), .O(gate70inter7));
  inv1  gate239(.a(N339), .O(gate70inter8));
  nand2 gate240(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate241(.a(s_5), .b(gate70inter3), .O(gate70inter10));
  nor2  gate242(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate243(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate244(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );

  xor2  gate287(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate288(.a(gate74inter0), .b(s_12), .O(gate74inter1));
  and2  gate289(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate290(.a(s_12), .O(gate74inter3));
  inv1  gate291(.a(s_13), .O(gate74inter4));
  nand2 gate292(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate293(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate294(.a(N315), .O(gate74inter7));
  inv1  gate295(.a(N347), .O(gate74inter8));
  nand2 gate296(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate297(.a(s_13), .b(gate74inter3), .O(gate74inter10));
  nor2  gate298(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate299(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate300(.a(gate74inter12), .b(gate74inter1), .O(N367));
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );

  xor2  gate301(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate302(.a(gate173inter0), .b(s_14), .O(gate173inter1));
  and2  gate303(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate304(.a(s_14), .O(gate173inter3));
  inv1  gate305(.a(s_15), .O(gate173inter4));
  nand2 gate306(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate307(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate308(.a(N9), .O(gate173inter7));
  inv1  gate309(.a(N694), .O(gate173inter8));
  nand2 gate310(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate311(.a(s_15), .b(gate173inter3), .O(gate173inter10));
  nor2  gate312(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate313(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate314(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );

  xor2  gate413(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate414(.a(gate188inter0), .b(s_30), .O(gate188inter1));
  and2  gate415(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate416(.a(s_30), .O(gate188inter3));
  inv1  gate417(.a(s_31), .O(gate188inter4));
  nand2 gate418(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate419(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate420(.a(N69), .O(gate188inter7));
  inv1  gate421(.a(N709), .O(gate188inter8));
  nand2 gate422(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate423(.a(s_31), .b(gate188inter3), .O(gate188inter10));
  nor2  gate424(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate425(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate426(.a(gate188inter12), .b(gate188inter1), .O(N741));
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );

  xor2  gate357(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate358(.a(gate197inter0), .b(s_22), .O(gate197inter1));
  and2  gate359(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate360(.a(s_22), .O(gate197inter3));
  inv1  gate361(.a(s_23), .O(gate197inter4));
  nand2 gate362(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate363(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate364(.a(N105), .O(gate197inter7));
  inv1  gate365(.a(N718), .O(gate197inter8));
  nand2 gate366(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate367(.a(s_23), .b(gate197inter3), .O(gate197inter10));
  nor2  gate368(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate369(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate370(.a(gate197inter12), .b(gate197inter1), .O(N750));
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate371(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate372(.a(gate201inter0), .b(s_24), .O(gate201inter1));
  and2  gate373(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate374(.a(s_24), .O(gate201inter3));
  inv1  gate375(.a(s_25), .O(gate201inter4));
  nand2 gate376(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate377(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate378(.a(N121), .O(gate201inter7));
  inv1  gate379(.a(N722), .O(gate201inter8));
  nand2 gate380(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate381(.a(s_25), .b(gate201inter3), .O(gate201inter10));
  nor2  gate382(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate383(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate384(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule