module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate357(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate358(.a(gate22inter0), .b(s_28), .O(gate22inter1));
  and2  gate359(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate360(.a(s_28), .O(gate22inter3));
  inv1  gate361(.a(s_29), .O(gate22inter4));
  nand2 gate362(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate363(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate364(.a(N122), .O(gate22inter7));
  inv1  gate365(.a(N17), .O(gate22inter8));
  nand2 gate366(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate367(.a(s_29), .b(gate22inter3), .O(gate22inter10));
  nor2  gate368(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate369(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate370(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate259(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate260(.a(gate36inter0), .b(s_14), .O(gate36inter1));
  and2  gate261(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate262(.a(s_14), .O(gate36inter3));
  inv1  gate263(.a(s_15), .O(gate36inter4));
  nand2 gate264(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate265(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate266(.a(N60), .O(gate36inter7));
  inv1  gate267(.a(N135), .O(gate36inter8));
  nand2 gate268(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate269(.a(s_15), .b(gate36inter3), .O(gate36inter10));
  nor2  gate270(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate271(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate272(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate287(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate288(.a(gate38inter0), .b(s_18), .O(gate38inter1));
  and2  gate289(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate290(.a(s_18), .O(gate38inter3));
  inv1  gate291(.a(s_19), .O(gate38inter4));
  nand2 gate292(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate293(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate294(.a(N73), .O(gate38inter7));
  inv1  gate295(.a(N139), .O(gate38inter8));
  nand2 gate296(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate297(.a(s_19), .b(gate38inter3), .O(gate38inter10));
  nor2  gate298(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate299(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate300(.a(gate38inter12), .b(gate38inter1), .O(N191));

  xor2  gate315(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate316(.a(gate39inter0), .b(s_22), .O(gate39inter1));
  and2  gate317(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate318(.a(s_22), .O(gate39inter3));
  inv1  gate319(.a(s_23), .O(gate39inter4));
  nand2 gate320(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate321(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate322(.a(N79), .O(gate39inter7));
  inv1  gate323(.a(N139), .O(gate39inter8));
  nand2 gate324(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate325(.a(s_23), .b(gate39inter3), .O(gate39inter10));
  nor2  gate326(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate327(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate328(.a(gate39inter12), .b(gate39inter1), .O(N192));
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate413(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate414(.a(gate50inter0), .b(s_36), .O(gate50inter1));
  and2  gate415(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate416(.a(s_36), .O(gate50inter3));
  inv1  gate417(.a(s_37), .O(gate50inter4));
  nand2 gate418(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate419(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate420(.a(N203), .O(gate50inter7));
  inv1  gate421(.a(N154), .O(gate50inter8));
  nand2 gate422(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate423(.a(s_37), .b(gate50inter3), .O(gate50inter10));
  nor2  gate424(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate425(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate426(.a(gate50inter12), .b(gate50inter1), .O(N224));

  xor2  gate273(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate274(.a(gate51inter0), .b(s_16), .O(gate51inter1));
  and2  gate275(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate276(.a(s_16), .O(gate51inter3));
  inv1  gate277(.a(s_17), .O(gate51inter4));
  nand2 gate278(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate279(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate280(.a(N203), .O(gate51inter7));
  inv1  gate281(.a(N159), .O(gate51inter8));
  nand2 gate282(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate283(.a(s_17), .b(gate51inter3), .O(gate51inter10));
  nor2  gate284(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate285(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate286(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );

  xor2  gate161(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate162(.a(gate55inter0), .b(s_0), .O(gate55inter1));
  and2  gate163(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate164(.a(s_0), .O(gate55inter3));
  inv1  gate165(.a(s_1), .O(gate55inter4));
  nand2 gate166(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate167(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate168(.a(N203), .O(gate55inter7));
  inv1  gate169(.a(N171), .O(gate55inter8));
  nand2 gate170(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate171(.a(s_1), .b(gate55inter3), .O(gate55inter10));
  nor2  gate172(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate173(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate174(.a(gate55inter12), .b(gate55inter1), .O(N239));
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );

  xor2  gate399(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate400(.a(gate58inter0), .b(s_34), .O(gate58inter1));
  and2  gate401(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate402(.a(s_34), .O(gate58inter3));
  inv1  gate403(.a(s_35), .O(gate58inter4));
  nand2 gate404(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate405(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate406(.a(N213), .O(gate58inter7));
  inv1  gate407(.a(N11), .O(gate58inter8));
  nand2 gate408(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate409(.a(s_35), .b(gate58inter3), .O(gate58inter10));
  nor2  gate410(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate411(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate412(.a(gate58inter12), .b(gate58inter1), .O(N246));
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );

  xor2  gate189(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate190(.a(gate66inter0), .b(s_4), .O(gate66inter1));
  and2  gate191(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate192(.a(s_4), .O(gate66inter3));
  inv1  gate193(.a(s_5), .O(gate66inter4));
  nand2 gate194(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate195(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate196(.a(N213), .O(gate66inter7));
  inv1  gate197(.a(N89), .O(gate66inter8));
  nand2 gate198(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate199(.a(s_5), .b(gate66inter3), .O(gate66inter10));
  nor2  gate200(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate201(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate202(.a(gate66inter12), .b(gate66inter1), .O(N258));
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate203(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate204(.a(gate68inter0), .b(s_6), .O(gate68inter1));
  and2  gate205(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate206(.a(s_6), .O(gate68inter3));
  inv1  gate207(.a(s_7), .O(gate68inter4));
  nand2 gate208(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate209(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate210(.a(N224), .O(gate68inter7));
  inv1  gate211(.a(N157), .O(gate68inter8));
  nand2 gate212(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate213(.a(s_7), .b(gate68inter3), .O(gate68inter10));
  nor2  gate214(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate215(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate216(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate385(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate386(.a(gate72inter0), .b(s_32), .O(gate72inter1));
  and2  gate387(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate388(.a(s_32), .O(gate72inter3));
  inv1  gate389(.a(s_33), .O(gate72inter4));
  nand2 gate390(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate391(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate392(.a(N233), .O(gate72inter7));
  inv1  gate393(.a(N187), .O(gate72inter8));
  nand2 gate394(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate395(.a(s_33), .b(gate72inter3), .O(gate72inter10));
  nor2  gate396(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate397(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate398(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );

  xor2  gate329(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate330(.a(gate76inter0), .b(s_24), .O(gate76inter1));
  and2  gate331(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate332(.a(s_24), .O(gate76inter3));
  inv1  gate333(.a(s_25), .O(gate76inter4));
  nand2 gate334(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate335(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate336(.a(N247), .O(gate76inter7));
  inv1  gate337(.a(N195), .O(gate76inter8));
  nand2 gate338(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate339(.a(s_25), .b(gate76inter3), .O(gate76inter10));
  nor2  gate340(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate341(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate342(.a(gate76inter12), .b(gate76inter1), .O(N282));
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate231(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate232(.a(gate80inter0), .b(s_10), .O(gate80inter1));
  and2  gate233(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate234(.a(s_10), .O(gate80inter3));
  inv1  gate235(.a(s_11), .O(gate80inter4));
  nand2 gate236(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate237(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate238(.a(N233), .O(gate80inter7));
  inv1  gate239(.a(N188), .O(gate80inter8));
  nand2 gate240(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate241(.a(s_11), .b(gate80inter3), .O(gate80inter10));
  nor2  gate242(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate243(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate244(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate441(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate442(.a(gate83inter0), .b(s_40), .O(gate83inter1));
  and2  gate443(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate444(.a(s_40), .O(gate83inter3));
  inv1  gate445(.a(s_41), .O(gate83inter4));
  nand2 gate446(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate447(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate448(.a(N243), .O(gate83inter7));
  inv1  gate449(.a(N194), .O(gate83inter8));
  nand2 gate450(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate451(.a(s_41), .b(gate83inter3), .O(gate83inter10));
  nor2  gate452(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate453(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate454(.a(gate83inter12), .b(gate83inter1), .O(N293));

  xor2  gate175(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate176(.a(gate84inter0), .b(s_2), .O(gate84inter1));
  and2  gate177(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate178(.a(s_2), .O(gate84inter3));
  inv1  gate179(.a(s_3), .O(gate84inter4));
  nand2 gate180(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate181(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate182(.a(N247), .O(gate84inter7));
  inv1  gate183(.a(N196), .O(gate84inter8));
  nand2 gate184(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate185(.a(s_3), .b(gate84inter3), .O(gate84inter10));
  nor2  gate186(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate187(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate188(.a(gate84inter12), .b(gate84inter1), .O(N294));

  xor2  gate245(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate246(.a(gate85inter0), .b(s_12), .O(gate85inter1));
  and2  gate247(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate248(.a(s_12), .O(gate85inter3));
  inv1  gate249(.a(s_13), .O(gate85inter4));
  nand2 gate250(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate251(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate252(.a(N251), .O(gate85inter7));
  inv1  gate253(.a(N198), .O(gate85inter8));
  nand2 gate254(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate255(.a(s_13), .b(gate85inter3), .O(gate85inter10));
  nor2  gate256(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate257(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate258(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate427(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate428(.a(gate99inter0), .b(s_38), .O(gate99inter1));
  and2  gate429(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate430(.a(s_38), .O(gate99inter3));
  inv1  gate431(.a(s_39), .O(gate99inter4));
  nand2 gate432(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate433(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate434(.a(N309), .O(gate99inter7));
  inv1  gate435(.a(N260), .O(gate99inter8));
  nand2 gate436(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate437(.a(s_39), .b(gate99inter3), .O(gate99inter10));
  nor2  gate438(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate439(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate440(.a(gate99inter12), .b(gate99inter1), .O(N330));
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );

  xor2  gate371(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate372(.a(gate125inter0), .b(s_30), .O(gate125inter1));
  and2  gate373(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate374(.a(s_30), .O(gate125inter3));
  inv1  gate375(.a(s_31), .O(gate125inter4));
  nand2 gate376(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate377(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate378(.a(N343), .O(gate125inter7));
  inv1  gate379(.a(N308), .O(gate125inter8));
  nand2 gate380(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate381(.a(s_31), .b(gate125inter3), .O(gate125inter10));
  nor2  gate382(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate383(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate384(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate301(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate302(.a(gate129inter0), .b(s_20), .O(gate129inter1));
  and2  gate303(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate304(.a(s_20), .O(gate129inter3));
  inv1  gate305(.a(s_21), .O(gate129inter4));
  nand2 gate306(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate307(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate308(.a(N14), .O(gate129inter7));
  inv1  gate309(.a(N360), .O(gate129inter8));
  nand2 gate310(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate311(.a(s_21), .b(gate129inter3), .O(gate129inter10));
  nor2  gate312(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate313(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate314(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );

  xor2  gate217(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate218(.a(gate133inter0), .b(s_8), .O(gate133inter1));
  and2  gate219(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate220(.a(s_8), .O(gate133inter3));
  inv1  gate221(.a(s_9), .O(gate133inter4));
  nand2 gate222(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate223(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate224(.a(N360), .O(gate133inter7));
  inv1  gate225(.a(N66), .O(gate133inter8));
  nand2 gate226(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate227(.a(s_9), .b(gate133inter3), .O(gate133inter10));
  nor2  gate228(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate229(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate230(.a(gate133inter12), .b(gate133inter1), .O(N375));

  xor2  gate343(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate344(.a(gate134inter0), .b(s_26), .O(gate134inter1));
  and2  gate345(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate346(.a(s_26), .O(gate134inter3));
  inv1  gate347(.a(s_27), .O(gate134inter4));
  nand2 gate348(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate349(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate350(.a(N360), .O(gate134inter7));
  inv1  gate351(.a(N79), .O(gate134inter8));
  nand2 gate352(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate353(.a(s_27), .b(gate134inter3), .O(gate134inter10));
  nor2  gate354(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate355(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate356(.a(gate134inter12), .b(gate134inter1), .O(N376));
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule