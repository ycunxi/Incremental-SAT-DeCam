module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12, gate851inter0, gate851inter1, gate851inter2, gate851inter3, gate851inter4, gate851inter5, gate851inter6, gate851inter7, gate851inter8, gate851inter9, gate851inter10, gate851inter11, gate851inter12, gate556inter0, gate556inter1, gate556inter2, gate556inter3, gate556inter4, gate556inter5, gate556inter6, gate556inter7, gate556inter8, gate556inter9, gate556inter10, gate556inter11, gate556inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate539inter0, gate539inter1, gate539inter2, gate539inter3, gate539inter4, gate539inter5, gate539inter6, gate539inter7, gate539inter8, gate539inter9, gate539inter10, gate539inter11, gate539inter12, gate380inter0, gate380inter1, gate380inter2, gate380inter3, gate380inter4, gate380inter5, gate380inter6, gate380inter7, gate380inter8, gate380inter9, gate380inter10, gate380inter11, gate380inter12, gate570inter0, gate570inter1, gate570inter2, gate570inter3, gate570inter4, gate570inter5, gate570inter6, gate570inter7, gate570inter8, gate570inter9, gate570inter10, gate570inter11, gate570inter12, gate561inter0, gate561inter1, gate561inter2, gate561inter3, gate561inter4, gate561inter5, gate561inter6, gate561inter7, gate561inter8, gate561inter9, gate561inter10, gate561inter11, gate561inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate608inter0, gate608inter1, gate608inter2, gate608inter3, gate608inter4, gate608inter5, gate608inter6, gate608inter7, gate608inter8, gate608inter9, gate608inter10, gate608inter11, gate608inter12, gate650inter0, gate650inter1, gate650inter2, gate650inter3, gate650inter4, gate650inter5, gate650inter6, gate650inter7, gate650inter8, gate650inter9, gate650inter10, gate650inter11, gate650inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate540inter0, gate540inter1, gate540inter2, gate540inter3, gate540inter4, gate540inter5, gate540inter6, gate540inter7, gate540inter8, gate540inter9, gate540inter10, gate540inter11, gate540inter12, gate765inter0, gate765inter1, gate765inter2, gate765inter3, gate765inter4, gate765inter5, gate765inter6, gate765inter7, gate765inter8, gate765inter9, gate765inter10, gate765inter11, gate765inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate758inter0, gate758inter1, gate758inter2, gate758inter3, gate758inter4, gate758inter5, gate758inter6, gate758inter7, gate758inter8, gate758inter9, gate758inter10, gate758inter11, gate758inter12, gate616inter0, gate616inter1, gate616inter2, gate616inter3, gate616inter4, gate616inter5, gate616inter6, gate616inter7, gate616inter8, gate616inter9, gate616inter10, gate616inter11, gate616inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate800inter0, gate800inter1, gate800inter2, gate800inter3, gate800inter4, gate800inter5, gate800inter6, gate800inter7, gate800inter8, gate800inter9, gate800inter10, gate800inter11, gate800inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate843inter0, gate843inter1, gate843inter2, gate843inter3, gate843inter4, gate843inter5, gate843inter6, gate843inter7, gate843inter8, gate843inter9, gate843inter10, gate843inter11, gate843inter12, gate357inter0, gate357inter1, gate357inter2, gate357inter3, gate357inter4, gate357inter5, gate357inter6, gate357inter7, gate357inter8, gate357inter9, gate357inter10, gate357inter11, gate357inter12, gate818inter0, gate818inter1, gate818inter2, gate818inter3, gate818inter4, gate818inter5, gate818inter6, gate818inter7, gate818inter8, gate818inter9, gate818inter10, gate818inter11, gate818inter12, gate819inter0, gate819inter1, gate819inter2, gate819inter3, gate819inter4, gate819inter5, gate819inter6, gate819inter7, gate819inter8, gate819inter9, gate819inter10, gate819inter11, gate819inter12, gate324inter0, gate324inter1, gate324inter2, gate324inter3, gate324inter4, gate324inter5, gate324inter6, gate324inter7, gate324inter8, gate324inter9, gate324inter10, gate324inter11, gate324inter12, gate868inter0, gate868inter1, gate868inter2, gate868inter3, gate868inter4, gate868inter5, gate868inter6, gate868inter7, gate868inter8, gate868inter9, gate868inter10, gate868inter11, gate868inter12, gate814inter0, gate814inter1, gate814inter2, gate814inter3, gate814inter4, gate814inter5, gate814inter6, gate814inter7, gate814inter8, gate814inter9, gate814inter10, gate814inter11, gate814inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate524inter0, gate524inter1, gate524inter2, gate524inter3, gate524inter4, gate524inter5, gate524inter6, gate524inter7, gate524inter8, gate524inter9, gate524inter10, gate524inter11, gate524inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate626inter0, gate626inter1, gate626inter2, gate626inter3, gate626inter4, gate626inter5, gate626inter6, gate626inter7, gate626inter8, gate626inter9, gate626inter10, gate626inter11, gate626inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate797inter0, gate797inter1, gate797inter2, gate797inter3, gate797inter4, gate797inter5, gate797inter6, gate797inter7, gate797inter8, gate797inter9, gate797inter10, gate797inter11, gate797inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate351inter0, gate351inter1, gate351inter2, gate351inter3, gate351inter4, gate351inter5, gate351inter6, gate351inter7, gate351inter8, gate351inter9, gate351inter10, gate351inter11, gate351inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate541inter0, gate541inter1, gate541inter2, gate541inter3, gate541inter4, gate541inter5, gate541inter6, gate541inter7, gate541inter8, gate541inter9, gate541inter10, gate541inter11, gate541inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate817inter0, gate817inter1, gate817inter2, gate817inter3, gate817inter4, gate817inter5, gate817inter6, gate817inter7, gate817inter8, gate817inter9, gate817inter10, gate817inter11, gate817inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate804inter0, gate804inter1, gate804inter2, gate804inter3, gate804inter4, gate804inter5, gate804inter6, gate804inter7, gate804inter8, gate804inter9, gate804inter10, gate804inter11, gate804inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate587inter0, gate587inter1, gate587inter2, gate587inter3, gate587inter4, gate587inter5, gate587inter6, gate587inter7, gate587inter8, gate587inter9, gate587inter10, gate587inter11, gate587inter12, gate516inter0, gate516inter1, gate516inter2, gate516inter3, gate516inter4, gate516inter5, gate516inter6, gate516inter7, gate516inter8, gate516inter9, gate516inter10, gate516inter11, gate516inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate682inter0, gate682inter1, gate682inter2, gate682inter3, gate682inter4, gate682inter5, gate682inter6, gate682inter7, gate682inter8, gate682inter9, gate682inter10, gate682inter11, gate682inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate808inter0, gate808inter1, gate808inter2, gate808inter3, gate808inter4, gate808inter5, gate808inter6, gate808inter7, gate808inter8, gate808inter9, gate808inter10, gate808inter11, gate808inter12, gate586inter0, gate586inter1, gate586inter2, gate586inter3, gate586inter4, gate586inter5, gate586inter6, gate586inter7, gate586inter8, gate586inter9, gate586inter10, gate586inter11, gate586inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate355inter0, gate355inter1, gate355inter2, gate355inter3, gate355inter4, gate355inter5, gate355inter6, gate355inter7, gate355inter8, gate355inter9, gate355inter10, gate355inter11, gate355inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate677inter0, gate677inter1, gate677inter2, gate677inter3, gate677inter4, gate677inter5, gate677inter6, gate677inter7, gate677inter8, gate677inter9, gate677inter10, gate677inter11, gate677inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate378inter0, gate378inter1, gate378inter2, gate378inter3, gate378inter4, gate378inter5, gate378inter6, gate378inter7, gate378inter8, gate378inter9, gate378inter10, gate378inter11, gate378inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate519inter0, gate519inter1, gate519inter2, gate519inter3, gate519inter4, gate519inter5, gate519inter6, gate519inter7, gate519inter8, gate519inter9, gate519inter10, gate519inter11, gate519inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate528inter0, gate528inter1, gate528inter2, gate528inter3, gate528inter4, gate528inter5, gate528inter6, gate528inter7, gate528inter8, gate528inter9, gate528inter10, gate528inter11, gate528inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate864inter0, gate864inter1, gate864inter2, gate864inter3, gate864inter4, gate864inter5, gate864inter6, gate864inter7, gate864inter8, gate864inter9, gate864inter10, gate864inter11, gate864inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate526inter0, gate526inter1, gate526inter2, gate526inter3, gate526inter4, gate526inter5, gate526inter6, gate526inter7, gate526inter8, gate526inter9, gate526inter10, gate526inter11, gate526inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate816inter0, gate816inter1, gate816inter2, gate816inter3, gate816inter4, gate816inter5, gate816inter6, gate816inter7, gate816inter8, gate816inter9, gate816inter10, gate816inter11, gate816inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate794inter0, gate794inter1, gate794inter2, gate794inter3, gate794inter4, gate794inter5, gate794inter6, gate794inter7, gate794inter8, gate794inter9, gate794inter10, gate794inter11, gate794inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate879inter0, gate879inter1, gate879inter2, gate879inter3, gate879inter4, gate879inter5, gate879inter6, gate879inter7, gate879inter8, gate879inter9, gate879inter10, gate879inter11, gate879inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate769inter0, gate769inter1, gate769inter2, gate769inter3, gate769inter4, gate769inter5, gate769inter6, gate769inter7, gate769inter8, gate769inter9, gate769inter10, gate769inter11, gate769inter12, gate366inter0, gate366inter1, gate366inter2, gate366inter3, gate366inter4, gate366inter5, gate366inter6, gate366inter7, gate366inter8, gate366inter9, gate366inter10, gate366inter11, gate366inter12, gate576inter0, gate576inter1, gate576inter2, gate576inter3, gate576inter4, gate576inter5, gate576inter6, gate576inter7, gate576inter8, gate576inter9, gate576inter10, gate576inter11, gate576inter12, gate306inter0, gate306inter1, gate306inter2, gate306inter3, gate306inter4, gate306inter5, gate306inter6, gate306inter7, gate306inter8, gate306inter9, gate306inter10, gate306inter11, gate306inter12, gate683inter0, gate683inter1, gate683inter2, gate683inter3, gate683inter4, gate683inter5, gate683inter6, gate683inter7, gate683inter8, gate683inter9, gate683inter10, gate683inter11, gate683inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate340inter0, gate340inter1, gate340inter2, gate340inter3, gate340inter4, gate340inter5, gate340inter6, gate340inter7, gate340inter8, gate340inter9, gate340inter10, gate340inter11, gate340inter12, gate341inter0, gate341inter1, gate341inter2, gate341inter3, gate341inter4, gate341inter5, gate341inter6, gate341inter7, gate341inter8, gate341inter9, gate341inter10, gate341inter11, gate341inter12, gate807inter0, gate807inter1, gate807inter2, gate807inter3, gate807inter4, gate807inter5, gate807inter6, gate807inter7, gate807inter8, gate807inter9, gate807inter10, gate807inter11, gate807inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate530inter0, gate530inter1, gate530inter2, gate530inter3, gate530inter4, gate530inter5, gate530inter6, gate530inter7, gate530inter8, gate530inter9, gate530inter10, gate530inter11, gate530inter12, gate320inter0, gate320inter1, gate320inter2, gate320inter3, gate320inter4, gate320inter5, gate320inter6, gate320inter7, gate320inter8, gate320inter9, gate320inter10, gate320inter11, gate320inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate600inter0, gate600inter1, gate600inter2, gate600inter3, gate600inter4, gate600inter5, gate600inter6, gate600inter7, gate600inter8, gate600inter9, gate600inter10, gate600inter11, gate600inter12, gate370inter0, gate370inter1, gate370inter2, gate370inter3, gate370inter4, gate370inter5, gate370inter6, gate370inter7, gate370inter8, gate370inter9, gate370inter10, gate370inter11, gate370inter12, gate605inter0, gate605inter1, gate605inter2, gate605inter3, gate605inter4, gate605inter5, gate605inter6, gate605inter7, gate605inter8, gate605inter9, gate605inter10, gate605inter11, gate605inter12, gate801inter0, gate801inter1, gate801inter2, gate801inter3, gate801inter4, gate801inter5, gate801inter6, gate801inter7, gate801inter8, gate801inter9, gate801inter10, gate801inter11, gate801inter12, gate305inter0, gate305inter1, gate305inter2, gate305inter3, gate305inter4, gate305inter5, gate305inter6, gate305inter7, gate305inter8, gate305inter9, gate305inter10, gate305inter11, gate305inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12, gate867inter0, gate867inter1, gate867inter2, gate867inter3, gate867inter4, gate867inter5, gate867inter6, gate867inter7, gate867inter8, gate867inter9, gate867inter10, gate867inter11, gate867inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );

  xor2  gate2001(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate2002(.a(gate77inter0), .b(s_160), .O(gate77inter1));
  and2  gate2003(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate2004(.a(s_160), .O(gate77inter3));
  inv1  gate2005(.a(s_161), .O(gate77inter4));
  nand2 gate2006(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2007(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2008(.a(N306), .O(gate77inter7));
  inv1  gate2009(.a(N331), .O(gate77inter8));
  nand2 gate2010(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2011(.a(s_161), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2012(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2013(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2014(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );

  xor2  gate1609(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate1610(.a(gate79inter0), .b(s_104), .O(gate79inter1));
  and2  gate1611(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate1612(.a(s_104), .O(gate79inter3));
  inv1  gate1613(.a(s_105), .O(gate79inter4));
  nand2 gate1614(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1615(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1616(.a(N306), .O(gate79inter7));
  inv1  gate1617(.a(N331), .O(gate79inter8));
  nand2 gate1618(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1619(.a(s_105), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1620(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1621(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1622(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate2071(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate2072(.a(gate96inter0), .b(s_170), .O(gate96inter1));
  and2  gate2073(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate2074(.a(s_170), .O(gate96inter3));
  inv1  gate2075(.a(s_171), .O(gate96inter4));
  nand2 gate2076(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2077(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2078(.a(N326), .O(gate96inter7));
  inv1  gate2079(.a(N277), .O(gate96inter8));
  nand2 gate2080(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2081(.a(s_171), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2082(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2083(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2084(.a(gate96inter12), .b(gate96inter1), .O(N601));
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );

  xor2  gate1147(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate1148(.a(gate99inter0), .b(s_38), .O(gate99inter1));
  and2  gate1149(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate1150(.a(s_38), .O(gate99inter3));
  inv1  gate1151(.a(s_39), .O(gate99inter4));
  nand2 gate1152(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1153(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1154(.a(N260), .O(gate99inter7));
  inv1  gate1155(.a(N300), .O(gate99inter8));
  nand2 gate1156(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1157(.a(s_39), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1158(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1159(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1160(.a(gate99inter12), .b(gate99inter1), .O(N608));
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );

  xor2  gate2281(.a(N612), .b(N53), .O(gate160inter0));
  nand2 gate2282(.a(gate160inter0), .b(s_200), .O(gate160inter1));
  and2  gate2283(.a(N612), .b(N53), .O(gate160inter2));
  inv1  gate2284(.a(s_200), .O(gate160inter3));
  inv1  gate2285(.a(s_201), .O(gate160inter4));
  nand2 gate2286(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2287(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2288(.a(N53), .O(gate160inter7));
  inv1  gate2289(.a(N612), .O(gate160inter8));
  nand2 gate2290(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2291(.a(s_201), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2292(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2293(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2294(.a(gate160inter12), .b(gate160inter1), .O(N899));

  xor2  gate2827(.a(N608), .b(N60), .O(gate161inter0));
  nand2 gate2828(.a(gate161inter0), .b(s_278), .O(gate161inter1));
  and2  gate2829(.a(N608), .b(N60), .O(gate161inter2));
  inv1  gate2830(.a(s_278), .O(gate161inter3));
  inv1  gate2831(.a(s_279), .O(gate161inter4));
  nand2 gate2832(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2833(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2834(.a(N60), .O(gate161inter7));
  inv1  gate2835(.a(N608), .O(gate161inter8));
  nand2 gate2836(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2837(.a(s_279), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2838(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2839(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2840(.a(gate161inter12), .b(gate161inter1), .O(N903));
nand2 gate162( .a(N49), .b(N612), .O(N907) );

  xor2  gate1035(.a(N608), .b(N56), .O(gate163inter0));
  nand2 gate1036(.a(gate163inter0), .b(s_22), .O(gate163inter1));
  and2  gate1037(.a(N608), .b(N56), .O(gate163inter2));
  inv1  gate1038(.a(s_22), .O(gate163inter3));
  inv1  gate1039(.a(s_23), .O(gate163inter4));
  nand2 gate1040(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1041(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1042(.a(N56), .O(gate163inter7));
  inv1  gate1043(.a(N608), .O(gate163inter8));
  nand2 gate1044(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1045(.a(s_23), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1046(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1047(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1048(.a(gate163inter12), .b(gate163inter1), .O(N910));
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );

  xor2  gate1651(.a(N888), .b(N619), .O(gate233inter0));
  nand2 gate1652(.a(gate233inter0), .b(s_110), .O(gate233inter1));
  and2  gate1653(.a(N888), .b(N619), .O(gate233inter2));
  inv1  gate1654(.a(s_110), .O(gate233inter3));
  inv1  gate1655(.a(s_111), .O(gate233inter4));
  nand2 gate1656(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1657(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1658(.a(N619), .O(gate233inter7));
  inv1  gate1659(.a(N888), .O(gate233inter8));
  nand2 gate1660(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1661(.a(s_111), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1662(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1663(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1664(.a(gate233inter12), .b(gate233inter1), .O(N1054));

  xor2  gate2099(.a(N889), .b(N616), .O(gate234inter0));
  nand2 gate2100(.a(gate234inter0), .b(s_174), .O(gate234inter1));
  and2  gate2101(.a(N889), .b(N616), .O(gate234inter2));
  inv1  gate2102(.a(s_174), .O(gate234inter3));
  inv1  gate2103(.a(s_175), .O(gate234inter4));
  nand2 gate2104(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2105(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2106(.a(N616), .O(gate234inter7));
  inv1  gate2107(.a(N889), .O(gate234inter8));
  nand2 gate2108(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2109(.a(s_175), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2110(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2111(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2112(.a(gate234inter12), .b(gate234inter1), .O(N1055));
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );

  xor2  gate1091(.a(N895), .b(N655), .O(gate237inter0));
  nand2 gate1092(.a(gate237inter0), .b(s_30), .O(gate237inter1));
  and2  gate1093(.a(N895), .b(N655), .O(gate237inter2));
  inv1  gate1094(.a(s_30), .O(gate237inter3));
  inv1  gate1095(.a(s_31), .O(gate237inter4));
  nand2 gate1096(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1097(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1098(.a(N655), .O(gate237inter7));
  inv1  gate1099(.a(N895), .O(gate237inter8));
  nand2 gate1100(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1101(.a(s_31), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1102(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1103(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1104(.a(gate237inter12), .b(gate237inter1), .O(N1067));

  xor2  gate2659(.a(N896), .b(N652), .O(gate238inter0));
  nand2 gate2660(.a(gate238inter0), .b(s_254), .O(gate238inter1));
  and2  gate2661(.a(N896), .b(N652), .O(gate238inter2));
  inv1  gate2662(.a(s_254), .O(gate238inter3));
  inv1  gate2663(.a(s_255), .O(gate238inter4));
  nand2 gate2664(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2665(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2666(.a(N652), .O(gate238inter7));
  inv1  gate2667(.a(N896), .O(gate238inter8));
  nand2 gate2668(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2669(.a(s_255), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2670(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2671(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2672(.a(gate238inter12), .b(gate238inter1), .O(N1068));
nand2 gate239( .a(N721), .b(N988), .O(N1119) );

  xor2  gate2897(.a(N989), .b(N718), .O(gate240inter0));
  nand2 gate2898(.a(gate240inter0), .b(s_288), .O(gate240inter1));
  and2  gate2899(.a(N989), .b(N718), .O(gate240inter2));
  inv1  gate2900(.a(s_288), .O(gate240inter3));
  inv1  gate2901(.a(s_289), .O(gate240inter4));
  nand2 gate2902(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2903(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2904(.a(N718), .O(gate240inter7));
  inv1  gate2905(.a(N989), .O(gate240inter8));
  nand2 gate2906(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2907(.a(s_289), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2908(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2909(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2910(.a(gate240inter12), .b(gate240inter1), .O(N1120));

  xor2  gate2645(.a(N991), .b(N727), .O(gate241inter0));
  nand2 gate2646(.a(gate241inter0), .b(s_252), .O(gate241inter1));
  and2  gate2647(.a(N991), .b(N727), .O(gate241inter2));
  inv1  gate2648(.a(s_252), .O(gate241inter3));
  inv1  gate2649(.a(s_253), .O(gate241inter4));
  nand2 gate2650(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2651(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2652(.a(N727), .O(gate241inter7));
  inv1  gate2653(.a(N991), .O(gate241inter8));
  nand2 gate2654(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2655(.a(s_253), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2656(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2657(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2658(.a(gate241inter12), .b(gate241inter1), .O(N1121));
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );

  xor2  gate1763(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate1764(.a(gate244inter0), .b(s_126), .O(gate244inter1));
  and2  gate1765(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate1766(.a(s_126), .O(gate244inter3));
  inv1  gate1767(.a(s_127), .O(gate244inter4));
  nand2 gate1768(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1769(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1770(.a(N736), .O(gate244inter7));
  inv1  gate1771(.a(N1003), .O(gate244inter8));
  nand2 gate1772(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1773(.a(s_127), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1774(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1775(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1776(.a(gate244inter12), .b(gate244inter1), .O(N1129));

  xor2  gate2463(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate2464(.a(gate245inter0), .b(s_226), .O(gate245inter1));
  and2  gate2465(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate2466(.a(s_226), .O(gate245inter3));
  inv1  gate2467(.a(s_227), .O(gate245inter4));
  nand2 gate2468(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2469(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2470(.a(N745), .O(gate245inter7));
  inv1  gate2471(.a(N1005), .O(gate245inter8));
  nand2 gate2472(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2473(.a(s_227), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2474(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2475(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2476(.a(gate245inter12), .b(gate245inter1), .O(N1130));
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );

  xor2  gate2253(.a(N1068), .b(N1067), .O(gate263inter0));
  nand2 gate2254(.a(gate263inter0), .b(s_196), .O(gate263inter1));
  and2  gate2255(.a(N1068), .b(N1067), .O(gate263inter2));
  inv1  gate2256(.a(s_196), .O(gate263inter3));
  inv1  gate2257(.a(s_197), .O(gate263inter4));
  nand2 gate2258(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2259(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2260(.a(N1067), .O(gate263inter7));
  inv1  gate2261(.a(N1068), .O(gate263inter8));
  nand2 gate2262(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2263(.a(s_197), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2264(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2265(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2266(.a(gate263inter12), .b(gate263inter1), .O(N1162));
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate2169(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate2170(.a(gate268inter0), .b(s_184), .O(gate268inter1));
  and2  gate2171(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate2172(.a(s_184), .O(gate268inter3));
  inv1  gate2173(.a(s_185), .O(gate268inter4));
  nand2 gate2174(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2175(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2176(.a(N921), .O(gate268inter7));
  inv1  gate2177(.a(N923), .O(gate268inter8));
  nand2 gate2178(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2179(.a(s_185), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2180(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2181(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2182(.a(gate268inter12), .b(gate268inter1), .O(N1171));

  xor2  gate2029(.a(N923), .b(N922), .O(gate269inter0));
  nand2 gate2030(.a(gate269inter0), .b(s_164), .O(gate269inter1));
  and2  gate2031(.a(N923), .b(N922), .O(gate269inter2));
  inv1  gate2032(.a(s_164), .O(gate269inter3));
  inv1  gate2033(.a(s_165), .O(gate269inter4));
  nand2 gate2034(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2035(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2036(.a(N922), .O(gate269inter7));
  inv1  gate2037(.a(N923), .O(gate269inter8));
  nand2 gate2038(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2039(.a(s_165), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2040(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2041(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2042(.a(gate269inter12), .b(gate269inter1), .O(N1188));
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate1175(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate1176(.a(gate273inter0), .b(s_42), .O(gate273inter1));
  and2  gate1177(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate1178(.a(s_42), .O(gate273inter3));
  inv1  gate1179(.a(s_43), .O(gate273inter4));
  nand2 gate1180(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1181(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1182(.a(N1013), .O(gate273inter7));
  inv1  gate1183(.a(N942), .O(gate273inter8));
  nand2 gate1184(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1185(.a(s_43), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1186(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1187(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1188(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate1497(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate1498(.a(gate275inter0), .b(s_88), .O(gate275inter1));
  and2  gate1499(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate1500(.a(s_88), .O(gate275inter3));
  inv1  gate1501(.a(s_89), .O(gate275inter4));
  nand2 gate1502(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1503(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1504(.a(N1016), .O(gate275inter7));
  inv1  gate1505(.a(N946), .O(gate275inter8));
  nand2 gate1506(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1507(.a(s_89), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1508(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1509(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1510(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate2505(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate2506(.a(gate277inter0), .b(s_232), .O(gate277inter1));
  and2  gate2507(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate2508(.a(s_232), .O(gate277inter3));
  inv1  gate2509(.a(s_233), .O(gate277inter4));
  nand2 gate2510(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2511(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2512(.a(N1019), .O(gate277inter7));
  inv1  gate2513(.a(N950), .O(gate277inter8));
  nand2 gate2514(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2515(.a(s_233), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2516(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2517(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2518(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );

  xor2  gate2155(.a(N968), .b(N1034), .O(gate286inter0));
  nand2 gate2156(.a(gate286inter0), .b(s_182), .O(gate286inter1));
  and2  gate2157(.a(N968), .b(N1034), .O(gate286inter2));
  inv1  gate2158(.a(s_182), .O(gate286inter3));
  inv1  gate2159(.a(s_183), .O(gate286inter4));
  nand2 gate2160(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2161(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2162(.a(N1034), .O(gate286inter7));
  inv1  gate2163(.a(N968), .O(gate286inter8));
  nand2 gate2164(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2165(.a(s_183), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2166(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2167(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2168(.a(gate286inter12), .b(gate286inter1), .O(N1221));
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );

  xor2  gate1903(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate1904(.a(gate297inter0), .b(s_146), .O(gate297inter1));
  and2  gate1905(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate1906(.a(s_146), .O(gate297inter3));
  inv1  gate1907(.a(s_147), .O(gate297inter4));
  nand2 gate1908(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate1909(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate1910(.a(N1119), .O(gate297inter7));
  inv1  gate1911(.a(N1120), .O(gate297inter8));
  nand2 gate1912(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate1913(.a(s_147), .b(gate297inter3), .O(gate297inter10));
  nor2  gate1914(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate1915(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate1916(.a(gate297inter12), .b(gate297inter1), .O(N1232));
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );

  xor2  gate2883(.a(N997), .b(N1046), .O(gate300inter0));
  nand2 gate2884(.a(gate300inter0), .b(s_286), .O(gate300inter1));
  and2  gate2885(.a(N997), .b(N1046), .O(gate300inter2));
  inv1  gate2886(.a(s_286), .O(gate300inter3));
  inv1  gate2887(.a(s_287), .O(gate300inter4));
  nand2 gate2888(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate2889(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate2890(.a(N1046), .O(gate300inter7));
  inv1  gate2891(.a(N997), .O(gate300inter8));
  nand2 gate2892(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate2893(.a(s_287), .b(gate300inter3), .O(gate300inter10));
  nor2  gate2894(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate2895(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate2896(.a(gate300inter12), .b(gate300inter1), .O(N1239));
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );

  xor2  gate2813(.a(N1131), .b(N1130), .O(gate305inter0));
  nand2 gate2814(.a(gate305inter0), .b(s_276), .O(gate305inter1));
  and2  gate2815(.a(N1131), .b(N1130), .O(gate305inter2));
  inv1  gate2816(.a(s_276), .O(gate305inter3));
  inv1  gate2817(.a(s_277), .O(gate305inter4));
  nand2 gate2818(.a(gate305inter4), .b(gate305inter3), .O(gate305inter5));
  nor2  gate2819(.a(gate305inter5), .b(gate305inter2), .O(gate305inter6));
  inv1  gate2820(.a(N1130), .O(gate305inter7));
  inv1  gate2821(.a(N1131), .O(gate305inter8));
  nand2 gate2822(.a(gate305inter8), .b(gate305inter7), .O(gate305inter9));
  nand2 gate2823(.a(s_277), .b(gate305inter3), .O(gate305inter10));
  nor2  gate2824(.a(gate305inter10), .b(gate305inter9), .O(gate305inter11));
  nor2  gate2825(.a(gate305inter11), .b(gate305inter6), .O(gate305inter12));
  nand2 gate2826(.a(gate305inter12), .b(gate305inter1), .O(N1246));

  xor2  gate2561(.a(N1133), .b(N1132), .O(gate306inter0));
  nand2 gate2562(.a(gate306inter0), .b(s_240), .O(gate306inter1));
  and2  gate2563(.a(N1133), .b(N1132), .O(gate306inter2));
  inv1  gate2564(.a(s_240), .O(gate306inter3));
  inv1  gate2565(.a(s_241), .O(gate306inter4));
  nand2 gate2566(.a(gate306inter4), .b(gate306inter3), .O(gate306inter5));
  nor2  gate2567(.a(gate306inter5), .b(gate306inter2), .O(gate306inter6));
  inv1  gate2568(.a(N1132), .O(gate306inter7));
  inv1  gate2569(.a(N1133), .O(gate306inter8));
  nand2 gate2570(.a(gate306inter8), .b(gate306inter7), .O(gate306inter9));
  nand2 gate2571(.a(s_241), .b(gate306inter3), .O(gate306inter10));
  nor2  gate2572(.a(gate306inter10), .b(gate306inter9), .O(gate306inter11));
  nor2  gate2573(.a(gate306inter11), .b(gate306inter6), .O(gate306inter12));
  nand2 gate2574(.a(gate306inter12), .b(gate306inter1), .O(N1249));
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );

  xor2  gate2057(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate2058(.a(gate316inter0), .b(s_168), .O(gate316inter1));
  and2  gate2059(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate2060(.a(s_168), .O(gate316inter3));
  inv1  gate2061(.a(s_169), .O(gate316inter4));
  nand2 gate2062(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate2063(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate2064(.a(N697), .O(gate316inter7));
  inv1  gate2065(.a(N1211), .O(gate316inter8));
  nand2 gate2066(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate2067(.a(s_169), .b(gate316inter3), .O(gate316inter10));
  nor2  gate2068(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate2069(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate2070(.a(gate316inter12), .b(gate316inter1), .O(N1312));

  xor2  gate2729(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate2730(.a(gate317inter0), .b(s_264), .O(gate317inter1));
  and2  gate2731(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate2732(.a(s_264), .O(gate317inter3));
  inv1  gate2733(.a(s_265), .O(gate317inter4));
  nand2 gate2734(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate2735(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate2736(.a(N700), .O(gate317inter7));
  inv1  gate2737(.a(N1213), .O(gate317inter8));
  nand2 gate2738(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate2739(.a(s_265), .b(gate317inter3), .O(gate317inter10));
  nor2  gate2740(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate2741(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate2742(.a(gate317inter12), .b(gate317inter1), .O(N1313));
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );

  xor2  gate2715(.a(N1223), .b(N709), .O(gate320inter0));
  nand2 gate2716(.a(gate320inter0), .b(s_262), .O(gate320inter1));
  and2  gate2717(.a(N1223), .b(N709), .O(gate320inter2));
  inv1  gate2718(.a(s_262), .O(gate320inter3));
  inv1  gate2719(.a(s_263), .O(gate320inter4));
  nand2 gate2720(.a(gate320inter4), .b(gate320inter3), .O(gate320inter5));
  nor2  gate2721(.a(gate320inter5), .b(gate320inter2), .O(gate320inter6));
  inv1  gate2722(.a(N709), .O(gate320inter7));
  inv1  gate2723(.a(N1223), .O(gate320inter8));
  nand2 gate2724(.a(gate320inter8), .b(gate320inter7), .O(gate320inter9));
  nand2 gate2725(.a(s_263), .b(gate320inter3), .O(gate320inter10));
  nor2  gate2726(.a(gate320inter10), .b(gate320inter9), .O(gate320inter11));
  nor2  gate2727(.a(gate320inter11), .b(gate320inter6), .O(gate320inter12));
  nand2 gate2728(.a(gate320inter12), .b(gate320inter1), .O(N1316));
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );

  xor2  gate2351(.a(N1228), .b(N715), .O(gate322inter0));
  nand2 gate2352(.a(gate322inter0), .b(s_210), .O(gate322inter1));
  and2  gate2353(.a(N1228), .b(N715), .O(gate322inter2));
  inv1  gate2354(.a(s_210), .O(gate322inter3));
  inv1  gate2355(.a(s_211), .O(gate322inter4));
  nand2 gate2356(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate2357(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate2358(.a(N715), .O(gate322inter7));
  inv1  gate2359(.a(N1228), .O(gate322inter8));
  nand2 gate2360(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate2361(.a(s_211), .b(gate322inter3), .O(gate322inter10));
  nor2  gate2362(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate2363(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate2364(.a(gate322inter12), .b(gate322inter1), .O(N1318));
inv1 gate323( .a(N1158), .O(N1319) );

  xor2  gate1371(.a(N1230), .b(N628), .O(gate324inter0));
  nand2 gate1372(.a(gate324inter0), .b(s_70), .O(gate324inter1));
  and2  gate1373(.a(N1230), .b(N628), .O(gate324inter2));
  inv1  gate1374(.a(s_70), .O(gate324inter3));
  inv1  gate1375(.a(s_71), .O(gate324inter4));
  nand2 gate1376(.a(gate324inter4), .b(gate324inter3), .O(gate324inter5));
  nor2  gate1377(.a(gate324inter5), .b(gate324inter2), .O(gate324inter6));
  inv1  gate1378(.a(N628), .O(gate324inter7));
  inv1  gate1379(.a(N1230), .O(gate324inter8));
  nand2 gate1380(.a(gate324inter8), .b(gate324inter7), .O(gate324inter9));
  nand2 gate1381(.a(s_71), .b(gate324inter3), .O(gate324inter10));
  nor2  gate1382(.a(gate324inter10), .b(gate324inter9), .O(gate324inter11));
  nor2  gate1383(.a(gate324inter11), .b(gate324inter6), .O(gate324inter12));
  nand2 gate1384(.a(gate324inter12), .b(gate324inter1), .O(N1322));
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );

  xor2  gate2183(.a(N1206), .b(N1309), .O(gate335inter0));
  nand2 gate2184(.a(gate335inter0), .b(s_186), .O(gate335inter1));
  and2  gate2185(.a(N1206), .b(N1309), .O(gate335inter2));
  inv1  gate2186(.a(s_186), .O(gate335inter3));
  inv1  gate2187(.a(s_187), .O(gate335inter4));
  nand2 gate2188(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate2189(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate2190(.a(N1309), .O(gate335inter7));
  inv1  gate2191(.a(N1206), .O(gate335inter8));
  nand2 gate2192(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate2193(.a(s_187), .b(gate335inter3), .O(gate335inter10));
  nor2  gate2194(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate2195(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate2196(.a(gate335inter12), .b(gate335inter1), .O(N1352));
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );

  xor2  gate951(.a(N1210), .b(N1311), .O(gate337inter0));
  nand2 gate952(.a(gate337inter0), .b(s_10), .O(gate337inter1));
  and2  gate953(.a(N1210), .b(N1311), .O(gate337inter2));
  inv1  gate954(.a(s_10), .O(gate337inter3));
  inv1  gate955(.a(s_11), .O(gate337inter4));
  nand2 gate956(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate957(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate958(.a(N1311), .O(gate337inter7));
  inv1  gate959(.a(N1210), .O(gate337inter8));
  nand2 gate960(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate961(.a(s_11), .b(gate337inter3), .O(gate337inter10));
  nor2  gate962(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate963(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate964(.a(gate337inter12), .b(gate337inter1), .O(N1358));
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );

  xor2  gate2603(.a(N1216), .b(N1314), .O(gate340inter0));
  nand2 gate2604(.a(gate340inter0), .b(s_246), .O(gate340inter1));
  and2  gate2605(.a(N1216), .b(N1314), .O(gate340inter2));
  inv1  gate2606(.a(s_246), .O(gate340inter3));
  inv1  gate2607(.a(s_247), .O(gate340inter4));
  nand2 gate2608(.a(gate340inter4), .b(gate340inter3), .O(gate340inter5));
  nor2  gate2609(.a(gate340inter5), .b(gate340inter2), .O(gate340inter6));
  inv1  gate2610(.a(N1314), .O(gate340inter7));
  inv1  gate2611(.a(N1216), .O(gate340inter8));
  nand2 gate2612(.a(gate340inter8), .b(gate340inter7), .O(gate340inter9));
  nand2 gate2613(.a(s_247), .b(gate340inter3), .O(gate340inter10));
  nor2  gate2614(.a(gate340inter10), .b(gate340inter9), .O(gate340inter11));
  nor2  gate2615(.a(gate340inter11), .b(gate340inter6), .O(gate340inter12));
  nand2 gate2616(.a(gate340inter12), .b(gate340inter1), .O(N1367));

  xor2  gate2617(.a(N1221), .b(N1315), .O(gate341inter0));
  nand2 gate2618(.a(gate341inter0), .b(s_248), .O(gate341inter1));
  and2  gate2619(.a(N1221), .b(N1315), .O(gate341inter2));
  inv1  gate2620(.a(s_248), .O(gate341inter3));
  inv1  gate2621(.a(s_249), .O(gate341inter4));
  nand2 gate2622(.a(gate341inter4), .b(gate341inter3), .O(gate341inter5));
  nor2  gate2623(.a(gate341inter5), .b(gate341inter2), .O(gate341inter6));
  inv1  gate2624(.a(N1315), .O(gate341inter7));
  inv1  gate2625(.a(N1221), .O(gate341inter8));
  nand2 gate2626(.a(gate341inter8), .b(gate341inter7), .O(gate341inter9));
  nand2 gate2627(.a(s_249), .b(gate341inter3), .O(gate341inter10));
  nor2  gate2628(.a(gate341inter10), .b(gate341inter9), .O(gate341inter11));
  nor2  gate2629(.a(gate341inter11), .b(gate341inter6), .O(gate341inter12));
  nand2 gate2630(.a(gate341inter12), .b(gate341inter1), .O(N1370));
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate1189(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate1190(.a(gate347inter0), .b(s_44), .O(gate347inter1));
  and2  gate1191(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate1192(.a(s_44), .O(gate347inter3));
  inv1  gate1193(.a(s_45), .O(gate347inter4));
  nand2 gate1194(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate1195(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate1196(.a(N1232), .O(gate347inter7));
  inv1  gate1197(.a(N990), .O(gate347inter8));
  nand2 gate1198(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate1199(.a(s_45), .b(gate347inter3), .O(gate347inter10));
  nor2  gate1200(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate1201(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate1202(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );

  xor2  gate1581(.a(N1242), .b(N1328), .O(gate351inter0));
  nand2 gate1582(.a(gate351inter0), .b(s_100), .O(gate351inter1));
  and2  gate1583(.a(N1242), .b(N1328), .O(gate351inter2));
  inv1  gate1584(.a(s_100), .O(gate351inter3));
  inv1  gate1585(.a(s_101), .O(gate351inter4));
  nand2 gate1586(.a(gate351inter4), .b(gate351inter3), .O(gate351inter5));
  nor2  gate1587(.a(gate351inter5), .b(gate351inter2), .O(gate351inter6));
  inv1  gate1588(.a(N1328), .O(gate351inter7));
  inv1  gate1589(.a(N1242), .O(gate351inter8));
  nand2 gate1590(.a(gate351inter8), .b(gate351inter7), .O(gate351inter9));
  nand2 gate1591(.a(s_101), .b(gate351inter3), .O(gate351inter10));
  nor2  gate1592(.a(gate351inter10), .b(gate351inter9), .O(gate351inter11));
  nor2  gate1593(.a(gate351inter11), .b(gate351inter6), .O(gate351inter12));
  nand2 gate1594(.a(gate351inter12), .b(gate351inter1), .O(N1393));
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );

  xor2  gate1987(.a(N1007), .b(N1246), .O(gate355inter0));
  nand2 gate1988(.a(gate355inter0), .b(s_158), .O(gate355inter1));
  and2  gate1989(.a(N1007), .b(N1246), .O(gate355inter2));
  inv1  gate1990(.a(s_158), .O(gate355inter3));
  inv1  gate1991(.a(s_159), .O(gate355inter4));
  nand2 gate1992(.a(gate355inter4), .b(gate355inter3), .O(gate355inter5));
  nor2  gate1993(.a(gate355inter5), .b(gate355inter2), .O(gate355inter6));
  inv1  gate1994(.a(N1246), .O(gate355inter7));
  inv1  gate1995(.a(N1007), .O(gate355inter8));
  nand2 gate1996(.a(gate355inter8), .b(gate355inter7), .O(gate355inter9));
  nand2 gate1997(.a(s_159), .b(gate355inter3), .O(gate355inter10));
  nor2  gate1998(.a(gate355inter10), .b(gate355inter9), .O(gate355inter11));
  nor2  gate1999(.a(gate355inter11), .b(gate355inter6), .O(gate355inter12));
  nand2 gate2000(.a(gate355inter12), .b(gate355inter1), .O(N1399));
inv1 gate356( .a(N1319), .O(N1409) );

  xor2  gate1329(.a(N1346), .b(N649), .O(gate357inter0));
  nand2 gate1330(.a(gate357inter0), .b(s_64), .O(gate357inter1));
  and2  gate1331(.a(N1346), .b(N649), .O(gate357inter2));
  inv1  gate1332(.a(s_64), .O(gate357inter3));
  inv1  gate1333(.a(s_65), .O(gate357inter4));
  nand2 gate1334(.a(gate357inter4), .b(gate357inter3), .O(gate357inter5));
  nor2  gate1335(.a(gate357inter5), .b(gate357inter2), .O(gate357inter6));
  inv1  gate1336(.a(N649), .O(gate357inter7));
  inv1  gate1337(.a(N1346), .O(gate357inter8));
  nand2 gate1338(.a(gate357inter8), .b(gate357inter7), .O(gate357inter9));
  nand2 gate1339(.a(s_65), .b(gate357inter3), .O(gate357inter10));
  nor2  gate1340(.a(gate357inter10), .b(gate357inter9), .O(gate357inter11));
  nor2  gate1341(.a(gate357inter11), .b(gate357inter6), .O(gate357inter12));
  nand2 gate1342(.a(gate357inter12), .b(gate357inter1), .O(N1412));
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );

  xor2  gate2673(.a(N1388), .b(N637), .O(gate362inter0));
  nand2 gate2674(.a(gate362inter0), .b(s_256), .O(gate362inter1));
  and2  gate2675(.a(N1388), .b(N637), .O(gate362inter2));
  inv1  gate2676(.a(s_256), .O(gate362inter3));
  inv1  gate2677(.a(s_257), .O(gate362inter4));
  nand2 gate2678(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate2679(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate2680(.a(N637), .O(gate362inter7));
  inv1  gate2681(.a(N1388), .O(gate362inter8));
  nand2 gate2682(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate2683(.a(s_257), .b(gate362inter3), .O(gate362inter10));
  nor2  gate2684(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate2685(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate2686(.a(gate362inter12), .b(gate362inter1), .O(N1434));
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );

  xor2  gate1567(.a(N1398), .b(N646), .O(gate364inter0));
  nand2 gate1568(.a(gate364inter0), .b(s_98), .O(gate364inter1));
  and2  gate1569(.a(N1398), .b(N646), .O(gate364inter2));
  inv1  gate1570(.a(s_98), .O(gate364inter3));
  inv1  gate1571(.a(s_99), .O(gate364inter4));
  nand2 gate1572(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate1573(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate1574(.a(N646), .O(gate364inter7));
  inv1  gate1575(.a(N1398), .O(gate364inter8));
  nand2 gate1576(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate1577(.a(s_99), .b(gate364inter3), .O(gate364inter10));
  nor2  gate1578(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate1579(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate1580(.a(gate364inter12), .b(gate364inter1), .O(N1439));
inv1 gate365( .a(N1344), .O(N1440) );

  xor2  gate2533(.a(N1148), .b(N1355), .O(gate366inter0));
  nand2 gate2534(.a(gate366inter0), .b(s_236), .O(gate366inter1));
  and2  gate2535(.a(N1148), .b(N1355), .O(gate366inter2));
  inv1  gate2536(.a(s_236), .O(gate366inter3));
  inv1  gate2537(.a(s_237), .O(gate366inter4));
  nand2 gate2538(.a(gate366inter4), .b(gate366inter3), .O(gate366inter5));
  nor2  gate2539(.a(gate366inter5), .b(gate366inter2), .O(gate366inter6));
  inv1  gate2540(.a(N1355), .O(gate366inter7));
  inv1  gate2541(.a(N1148), .O(gate366inter8));
  nand2 gate2542(.a(gate366inter8), .b(gate366inter7), .O(gate366inter9));
  nand2 gate2543(.a(s_237), .b(gate366inter3), .O(gate366inter10));
  nor2  gate2544(.a(gate366inter10), .b(gate366inter9), .O(gate366inter11));
  nor2  gate2545(.a(gate366inter11), .b(gate366inter6), .O(gate366inter12));
  nand2 gate2546(.a(gate366inter12), .b(gate366inter1), .O(N1443));
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );

  xor2  gate2771(.a(N1151), .b(N1358), .O(gate370inter0));
  nand2 gate2772(.a(gate370inter0), .b(s_270), .O(gate370inter1));
  and2  gate2773(.a(N1151), .b(N1358), .O(gate370inter2));
  inv1  gate2774(.a(s_270), .O(gate370inter3));
  inv1  gate2775(.a(s_271), .O(gate370inter4));
  nand2 gate2776(.a(gate370inter4), .b(gate370inter3), .O(gate370inter5));
  nor2  gate2777(.a(gate370inter5), .b(gate370inter2), .O(gate370inter6));
  inv1  gate2778(.a(N1358), .O(gate370inter7));
  inv1  gate2779(.a(N1151), .O(gate370inter8));
  nand2 gate2780(.a(gate370inter8), .b(gate370inter7), .O(gate370inter9));
  nand2 gate2781(.a(s_271), .b(gate370inter3), .O(gate370inter10));
  nor2  gate2782(.a(gate370inter10), .b(gate370inter9), .O(gate370inter11));
  nor2  gate2783(.a(gate370inter11), .b(gate370inter6), .O(gate370inter12));
  nand2 gate2784(.a(gate370inter12), .b(gate370inter1), .O(N1447));
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate1553(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate1554(.a(gate376inter0), .b(s_96), .O(gate376inter1));
  and2  gate1555(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate1556(.a(s_96), .O(gate376inter3));
  inv1  gate1557(.a(s_97), .O(gate376inter4));
  nand2 gate1558(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate1559(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate1560(.a(N1364), .O(gate376inter7));
  inv1  gate1561(.a(N1154), .O(gate376inter8));
  nand2 gate1562(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate1563(.a(s_97), .b(gate376inter3), .O(gate376inter10));
  nor2  gate1564(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate1565(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate1566(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );

  xor2  gate2043(.a(N1156), .b(N1373), .O(gate378inter0));
  nand2 gate2044(.a(gate378inter0), .b(s_166), .O(gate378inter1));
  and2  gate2045(.a(N1156), .b(N1373), .O(gate378inter2));
  inv1  gate2046(.a(s_166), .O(gate378inter3));
  inv1  gate2047(.a(s_167), .O(gate378inter4));
  nand2 gate2048(.a(gate378inter4), .b(gate378inter3), .O(gate378inter5));
  nor2  gate2049(.a(gate378inter5), .b(gate378inter2), .O(gate378inter6));
  inv1  gate2050(.a(N1373), .O(gate378inter7));
  inv1  gate2051(.a(N1156), .O(gate378inter8));
  nand2 gate2052(.a(gate378inter8), .b(gate378inter7), .O(gate378inter9));
  nand2 gate2053(.a(s_167), .b(gate378inter3), .O(gate378inter10));
  nor2  gate2054(.a(gate378inter10), .b(gate378inter9), .O(gate378inter11));
  nor2  gate2055(.a(gate378inter11), .b(gate378inter6), .O(gate378inter12));
  nand2 gate2056(.a(gate378inter12), .b(gate378inter1), .O(N1457));
inv1 gate379( .a(N1373), .O(N1458) );

  xor2  gate993(.a(N1157), .b(N1379), .O(gate380inter0));
  nand2 gate994(.a(gate380inter0), .b(s_16), .O(gate380inter1));
  and2  gate995(.a(N1157), .b(N1379), .O(gate380inter2));
  inv1  gate996(.a(s_16), .O(gate380inter3));
  inv1  gate997(.a(s_17), .O(gate380inter4));
  nand2 gate998(.a(gate380inter4), .b(gate380inter3), .O(gate380inter5));
  nor2  gate999(.a(gate380inter5), .b(gate380inter2), .O(gate380inter6));
  inv1  gate1000(.a(N1379), .O(gate380inter7));
  inv1  gate1001(.a(N1157), .O(gate380inter8));
  nand2 gate1002(.a(gate380inter8), .b(gate380inter7), .O(gate380inter9));
  nand2 gate1003(.a(s_17), .b(gate380inter3), .O(gate380inter10));
  nor2  gate1004(.a(gate380inter10), .b(gate380inter9), .O(gate380inter11));
  nor2  gate1005(.a(gate380inter11), .b(gate380inter6), .O(gate380inter12));
  nand2 gate1006(.a(gate380inter12), .b(gate380inter1), .O(N1459));
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate1133(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate1134(.a(gate383inter0), .b(s_36), .O(gate383inter1));
  and2  gate1135(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate1136(.a(s_36), .O(gate383inter3));
  inv1  gate1137(.a(s_37), .O(gate383inter4));
  nand2 gate1138(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate1139(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate1140(.a(N1393), .O(gate383inter7));
  inv1  gate1141(.a(N1161), .O(gate383inter8));
  nand2 gate1142(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate1143(.a(s_37), .b(gate383inter3), .O(gate383inter10));
  nor2  gate1144(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate1145(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate1146(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );

  xor2  gate1273(.a(N1433), .b(N1387), .O(gate390inter0));
  nand2 gate1274(.a(gate390inter0), .b(s_56), .O(gate390inter1));
  and2  gate1275(.a(N1433), .b(N1387), .O(gate390inter2));
  inv1  gate1276(.a(s_56), .O(gate390inter3));
  inv1  gate1277(.a(s_57), .O(gate390inter4));
  nand2 gate1278(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1279(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1280(.a(N1387), .O(gate390inter7));
  inv1  gate1281(.a(N1433), .O(gate390inter8));
  nand2 gate1282(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1283(.a(s_57), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1284(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1285(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1286(.a(gate390inter12), .b(gate390inter1), .O(N1472));
inv1 gate391( .a(N1390), .O(N1475) );

  xor2  gate1665(.a(N1240), .b(N1390), .O(gate392inter0));
  nand2 gate1666(.a(gate392inter0), .b(s_112), .O(gate392inter1));
  and2  gate1667(.a(N1240), .b(N1390), .O(gate392inter2));
  inv1  gate1668(.a(s_112), .O(gate392inter3));
  inv1  gate1669(.a(s_113), .O(gate392inter4));
  nand2 gate1670(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1671(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1672(.a(N1390), .O(gate392inter7));
  inv1  gate1673(.a(N1240), .O(gate392inter8));
  nand2 gate1674(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1675(.a(s_113), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1676(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1677(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1678(.a(gate392inter12), .b(gate392inter1), .O(N1476));

  xor2  gate965(.a(N1434), .b(N1389), .O(gate393inter0));
  nand2 gate966(.a(gate393inter0), .b(s_12), .O(gate393inter1));
  and2  gate967(.a(N1434), .b(N1389), .O(gate393inter2));
  inv1  gate968(.a(s_12), .O(gate393inter3));
  inv1  gate969(.a(s_13), .O(gate393inter4));
  nand2 gate970(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate971(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate972(.a(N1389), .O(gate393inter7));
  inv1  gate973(.a(N1434), .O(gate393inter8));
  nand2 gate974(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate975(.a(s_13), .b(gate393inter3), .O(gate393inter10));
  nor2  gate976(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate977(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate978(.a(gate393inter12), .b(gate393inter1), .O(N1478));

  xor2  gate1511(.a(N1439), .b(N1399), .O(gate394inter0));
  nand2 gate1512(.a(gate394inter0), .b(s_90), .O(gate394inter1));
  and2  gate1513(.a(N1439), .b(N1399), .O(gate394inter2));
  inv1  gate1514(.a(s_90), .O(gate394inter3));
  inv1  gate1515(.a(s_91), .O(gate394inter4));
  nand2 gate1516(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1517(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1518(.a(N1399), .O(gate394inter7));
  inv1  gate1519(.a(N1439), .O(gate394inter8));
  nand2 gate1520(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1521(.a(s_91), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1522(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1523(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1524(.a(gate394inter12), .b(gate394inter1), .O(N1481));
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );

  xor2  gate2323(.a(N1444), .b(N939), .O(gate396inter0));
  nand2 gate2324(.a(gate396inter0), .b(s_206), .O(gate396inter1));
  and2  gate2325(.a(N1444), .b(N939), .O(gate396inter2));
  inv1  gate2326(.a(s_206), .O(gate396inter3));
  inv1  gate2327(.a(s_207), .O(gate396inter4));
  nand2 gate2328(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2329(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2330(.a(N939), .O(gate396inter7));
  inv1  gate2331(.a(N1444), .O(gate396inter8));
  nand2 gate2332(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2333(.a(s_207), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2334(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2335(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2336(.a(gate396inter12), .b(gate396inter1), .O(N1487));

  xor2  gate1301(.a(N1446), .b(N935), .O(gate397inter0));
  nand2 gate1302(.a(gate397inter0), .b(s_60), .O(gate397inter1));
  and2  gate1303(.a(N1446), .b(N935), .O(gate397inter2));
  inv1  gate1304(.a(s_60), .O(gate397inter3));
  inv1  gate1305(.a(s_61), .O(gate397inter4));
  nand2 gate1306(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1307(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1308(.a(N935), .O(gate397inter7));
  inv1  gate1309(.a(N1446), .O(gate397inter8));
  nand2 gate1310(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1311(.a(s_61), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1312(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1313(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1314(.a(gate397inter12), .b(gate397inter1), .O(N1488));

  xor2  gate1721(.a(N1448), .b(N943), .O(gate398inter0));
  nand2 gate1722(.a(gate398inter0), .b(s_120), .O(gate398inter1));
  and2  gate1723(.a(N1448), .b(N943), .O(gate398inter2));
  inv1  gate1724(.a(s_120), .O(gate398inter3));
  inv1  gate1725(.a(s_121), .O(gate398inter4));
  nand2 gate1726(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1727(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1728(.a(N943), .O(gate398inter7));
  inv1  gate1729(.a(N1448), .O(gate398inter8));
  nand2 gate1730(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1731(.a(s_121), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1732(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1733(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1734(.a(gate398inter12), .b(gate398inter1), .O(N1489));
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );

  xor2  gate1875(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate1876(.a(gate402inter0), .b(s_142), .O(gate402inter1));
  and2  gate1877(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate1878(.a(s_142), .O(gate402inter3));
  inv1  gate1879(.a(s_143), .O(gate402inter4));
  nand2 gate1880(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1881(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1882(.a(N955), .O(gate402inter7));
  inv1  gate1883(.a(N1454), .O(gate402inter8));
  nand2 gate1884(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1885(.a(s_143), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1886(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1887(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1888(.a(gate402inter12), .b(gate402inter1), .O(N1493));
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );

  xor2  gate2113(.a(N1468), .b(N965), .O(gate408inter0));
  nand2 gate2114(.a(gate408inter0), .b(s_176), .O(gate408inter1));
  and2  gate2115(.a(N1468), .b(N965), .O(gate408inter2));
  inv1  gate2116(.a(s_176), .O(gate408inter3));
  inv1  gate2117(.a(s_177), .O(gate408inter4));
  nand2 gate2118(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2119(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2120(.a(N965), .O(gate408inter7));
  inv1  gate2121(.a(N1468), .O(gate408inter8));
  nand2 gate2122(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2123(.a(s_177), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2124(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2125(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2126(.a(gate408inter12), .b(gate408inter1), .O(N1500));

  xor2  gate1931(.a(N1470), .b(N973), .O(gate409inter0));
  nand2 gate1932(.a(gate409inter0), .b(s_150), .O(gate409inter1));
  and2  gate1933(.a(N1470), .b(N973), .O(gate409inter2));
  inv1  gate1934(.a(s_150), .O(gate409inter3));
  inv1  gate1935(.a(s_151), .O(gate409inter4));
  nand2 gate1936(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1937(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1938(.a(N973), .O(gate409inter7));
  inv1  gate1939(.a(N1470), .O(gate409inter8));
  nand2 gate1940(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1941(.a(s_151), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1942(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1943(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1944(.a(gate409inter12), .b(gate409inter1), .O(N1501));

  xor2  gate1595(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate1596(.a(gate410inter0), .b(s_102), .O(gate410inter1));
  and2  gate1597(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate1598(.a(s_102), .O(gate410inter3));
  inv1  gate1599(.a(s_103), .O(gate410inter4));
  nand2 gate1600(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1601(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1602(.a(N994), .O(gate410inter7));
  inv1  gate1603(.a(N1475), .O(gate410inter8));
  nand2 gate1604(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1605(.a(s_103), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1606(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1607(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1608(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );

  xor2  gate1413(.a(N1489), .b(N1447), .O(gate414inter0));
  nand2 gate1414(.a(gate414inter0), .b(s_76), .O(gate414inter1));
  and2  gate1415(.a(N1489), .b(N1447), .O(gate414inter2));
  inv1  gate1416(.a(s_76), .O(gate414inter3));
  inv1  gate1417(.a(s_77), .O(gate414inter4));
  nand2 gate1418(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1419(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1420(.a(N1447), .O(gate414inter7));
  inv1  gate1421(.a(N1489), .O(gate414inter8));
  nand2 gate1422(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1423(.a(s_77), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1424(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1425(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1426(.a(gate414inter12), .b(gate414inter1), .O(N1517));
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );

  xor2  gate2337(.a(N1495), .b(N1457), .O(gate418inter0));
  nand2 gate2338(.a(gate418inter0), .b(s_208), .O(gate418inter1));
  and2  gate2339(.a(N1495), .b(N1457), .O(gate418inter2));
  inv1  gate2340(.a(s_208), .O(gate418inter3));
  inv1  gate2341(.a(s_209), .O(gate418inter4));
  nand2 gate2342(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2343(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2344(.a(N1457), .O(gate418inter7));
  inv1  gate2345(.a(N1495), .O(gate418inter8));
  nand2 gate2346(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2347(.a(s_209), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2348(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2349(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2350(.a(gate418inter12), .b(gate418inter1), .O(N1526));

  xor2  gate2407(.a(N1496), .b(N1459), .O(gate419inter0));
  nand2 gate2408(.a(gate419inter0), .b(s_218), .O(gate419inter1));
  and2  gate2409(.a(N1496), .b(N1459), .O(gate419inter2));
  inv1  gate2410(.a(s_218), .O(gate419inter3));
  inv1  gate2411(.a(s_219), .O(gate419inter4));
  nand2 gate2412(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2413(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2414(.a(N1459), .O(gate419inter7));
  inv1  gate2415(.a(N1496), .O(gate419inter8));
  nand2 gate2416(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2417(.a(s_219), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2418(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2419(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2420(.a(gate419inter12), .b(gate419inter1), .O(N1527));
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate881(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate882(.a(gate421inter0), .b(s_0), .O(gate421inter1));
  and2  gate883(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate884(.a(s_0), .O(gate421inter3));
  inv1  gate885(.a(s_1), .O(gate421inter4));
  nand2 gate886(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate887(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate888(.a(N1462), .O(gate421inter7));
  inv1  gate889(.a(N1498), .O(gate421inter8));
  nand2 gate890(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate891(.a(s_1), .b(gate421inter3), .O(gate421inter10));
  nor2  gate892(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate893(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate894(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );

  xor2  gate1105(.a(N1501), .b(N1471), .O(gate425inter0));
  nand2 gate1106(.a(gate425inter0), .b(s_32), .O(gate425inter1));
  and2  gate1107(.a(N1501), .b(N1471), .O(gate425inter2));
  inv1  gate1108(.a(s_32), .O(gate425inter3));
  inv1  gate1109(.a(s_33), .O(gate425inter4));
  nand2 gate1110(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1111(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1112(.a(N1471), .O(gate425inter7));
  inv1  gate1113(.a(N1501), .O(gate425inter8));
  nand2 gate1114(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1115(.a(s_33), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1116(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1117(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1118(.a(gate425inter12), .b(gate425inter1), .O(N1534));
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );

  xor2  gate2085(.a(N1531), .b(N1484), .O(gate432inter0));
  nand2 gate2086(.a(gate432inter0), .b(s_172), .O(gate432inter1));
  and2  gate2087(.a(N1531), .b(N1484), .O(gate432inter2));
  inv1  gate2088(.a(s_172), .O(gate432inter3));
  inv1  gate2089(.a(s_173), .O(gate432inter4));
  nand2 gate2090(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2091(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2092(.a(N1484), .O(gate432inter7));
  inv1  gate2093(.a(N1531), .O(gate432inter8));
  nand2 gate2094(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2095(.a(s_173), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2096(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2097(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2098(.a(gate432inter12), .b(gate432inter1), .O(N1567));

  xor2  gate1749(.a(N1532), .b(N1481), .O(gate433inter0));
  nand2 gate1750(.a(gate433inter0), .b(s_124), .O(gate433inter1));
  and2  gate1751(.a(N1532), .b(N1481), .O(gate433inter2));
  inv1  gate1752(.a(s_124), .O(gate433inter3));
  inv1  gate1753(.a(s_125), .O(gate433inter4));
  nand2 gate1754(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1755(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1756(.a(N1481), .O(gate433inter7));
  inv1  gate1757(.a(N1532), .O(gate433inter8));
  nand2 gate1758(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1759(.a(s_125), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1760(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1761(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1762(.a(gate433inter12), .b(gate433inter1), .O(N1568));
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );

  xor2  gate1469(.a(N1568), .b(N1567), .O(gate442inter0));
  nand2 gate1470(.a(gate442inter0), .b(s_84), .O(gate442inter1));
  and2  gate1471(.a(N1568), .b(N1567), .O(gate442inter2));
  inv1  gate1472(.a(s_84), .O(gate442inter3));
  inv1  gate1473(.a(s_85), .O(gate442inter4));
  nand2 gate1474(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1475(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1476(.a(N1567), .O(gate442inter7));
  inv1  gate1477(.a(N1568), .O(gate442inter8));
  nand2 gate1478(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1479(.a(s_85), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1480(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1481(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1482(.a(gate442inter12), .b(gate442inter1), .O(N1596));
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );

  xor2  gate2911(.a(N1217), .b(N1606), .O(gate466inter0));
  nand2 gate2912(.a(gate466inter0), .b(s_290), .O(gate466inter1));
  and2  gate2913(.a(N1217), .b(N1606), .O(gate466inter2));
  inv1  gate2914(.a(s_290), .O(gate466inter3));
  inv1  gate2915(.a(s_291), .O(gate466inter4));
  nand2 gate2916(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2917(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2918(.a(N1606), .O(gate466inter7));
  inv1  gate2919(.a(N1217), .O(gate466inter8));
  nand2 gate2920(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2921(.a(s_291), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2922(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2923(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2924(.a(gate466inter12), .b(gate466inter1), .O(N1678));
inv1 gate467( .a(N1606), .O(N1679) );

  xor2  gate1539(.a(N1219), .b(N1609), .O(gate468inter0));
  nand2 gate1540(.a(gate468inter0), .b(s_94), .O(gate468inter1));
  and2  gate1541(.a(N1219), .b(N1609), .O(gate468inter2));
  inv1  gate1542(.a(s_94), .O(gate468inter3));
  inv1  gate1543(.a(s_95), .O(gate468inter4));
  nand2 gate1544(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1545(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1546(.a(N1609), .O(gate468inter7));
  inv1  gate1547(.a(N1219), .O(gate468inter8));
  nand2 gate1548(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1549(.a(s_95), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1550(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1551(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1552(.a(gate468inter12), .b(gate468inter1), .O(N1680));
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );

  xor2  gate2869(.a(N1672), .b(N643), .O(gate476inter0));
  nand2 gate2870(.a(gate476inter0), .b(s_284), .O(gate476inter1));
  and2  gate2871(.a(N1672), .b(N643), .O(gate476inter2));
  inv1  gate2872(.a(s_284), .O(gate476inter3));
  inv1  gate2873(.a(s_285), .O(gate476inter4));
  nand2 gate2874(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2875(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2876(.a(N643), .O(gate476inter7));
  inv1  gate2877(.a(N1672), .O(gate476inter8));
  nand2 gate2878(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2879(.a(s_285), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2880(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2881(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2882(.a(gate476inter12), .b(gate476inter1), .O(N1706));
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );

  xor2  gate2491(.a(N1677), .b(N1651), .O(gate480inter0));
  nand2 gate2492(.a(gate480inter0), .b(s_230), .O(gate480inter1));
  and2  gate2493(.a(N1677), .b(N1651), .O(gate480inter2));
  inv1  gate2494(.a(s_230), .O(gate480inter3));
  inv1  gate2495(.a(s_231), .O(gate480inter4));
  nand2 gate2496(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2497(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2498(.a(N1651), .O(gate480inter7));
  inv1  gate2499(.a(N1677), .O(gate480inter8));
  nand2 gate2500(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2501(.a(s_231), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2502(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2503(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2504(.a(gate480inter12), .b(gate480inter1), .O(N1710));
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );

  xor2  gate1525(.a(N1688), .b(N1638), .O(gate488inter0));
  nand2 gate1526(.a(gate488inter0), .b(s_92), .O(gate488inter1));
  and2  gate1527(.a(N1688), .b(N1638), .O(gate488inter2));
  inv1  gate1528(.a(s_92), .O(gate488inter3));
  inv1  gate1529(.a(s_93), .O(gate488inter4));
  nand2 gate1530(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1531(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1532(.a(N1638), .O(gate488inter7));
  inv1  gate1533(.a(N1688), .O(gate488inter8));
  nand2 gate1534(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1535(.a(s_93), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1536(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1537(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1538(.a(gate488inter12), .b(gate488inter1), .O(N1723));
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );

  xor2  gate895(.a(N1528), .b(N1685), .O(gate494inter0));
  nand2 gate896(.a(gate494inter0), .b(s_2), .O(gate494inter1));
  and2  gate897(.a(N1528), .b(N1685), .O(gate494inter2));
  inv1  gate898(.a(s_2), .O(gate494inter3));
  inv1  gate899(.a(s_3), .O(gate494inter4));
  nand2 gate900(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate901(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate902(.a(N1685), .O(gate494inter7));
  inv1  gate903(.a(N1528), .O(gate494inter8));
  nand2 gate904(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate905(.a(s_3), .b(gate494inter3), .O(gate494inter10));
  nor2  gate906(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate907(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate908(.a(gate494inter12), .b(gate494inter1), .O(N1740));
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );

  xor2  gate1973(.a(N1730), .b(N1701), .O(gate505inter0));
  nand2 gate1974(.a(gate505inter0), .b(s_156), .O(gate505inter1));
  and2  gate1975(.a(N1730), .b(N1701), .O(gate505inter2));
  inv1  gate1976(.a(s_156), .O(gate505inter3));
  inv1  gate1977(.a(s_157), .O(gate505inter4));
  nand2 gate1978(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1979(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1980(.a(N1701), .O(gate505inter7));
  inv1  gate1981(.a(N1730), .O(gate505inter8));
  nand2 gate1982(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1983(.a(s_157), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1984(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1985(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1986(.a(gate505inter12), .b(gate505inter1), .O(N1764));
inv1 gate506( .a(N1717), .O(N1768) );

  xor2  gate1231(.a(N1741), .b(N1472), .O(gate507inter0));
  nand2 gate1232(.a(gate507inter0), .b(s_50), .O(gate507inter1));
  and2  gate1233(.a(N1741), .b(N1472), .O(gate507inter2));
  inv1  gate1234(.a(s_50), .O(gate507inter3));
  inv1  gate1235(.a(s_51), .O(gate507inter4));
  nand2 gate1236(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1237(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1238(.a(N1472), .O(gate507inter7));
  inv1  gate1239(.a(N1741), .O(gate507inter8));
  nand2 gate1240(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1241(.a(s_51), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1242(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1243(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1244(.a(gate507inter12), .b(gate507inter1), .O(N1769));

  xor2  gate2141(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate2142(.a(gate508inter0), .b(s_180), .O(gate508inter1));
  and2  gate2143(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate2144(.a(s_180), .O(gate508inter3));
  inv1  gate2145(.a(s_181), .O(gate508inter4));
  nand2 gate2146(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2147(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2148(.a(N1723), .O(gate508inter7));
  inv1  gate2149(.a(N1413), .O(gate508inter8));
  nand2 gate2150(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2151(.a(s_181), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2152(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2153(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2154(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate2379(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate2380(.a(gate513inter0), .b(s_214), .O(gate513inter1));
  and2  gate2381(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate2382(.a(s_214), .O(gate513inter3));
  inv1  gate2383(.a(s_215), .O(gate513inter4));
  nand2 gate2384(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2385(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2386(.a(N1731), .O(gate513inter7));
  inv1  gate2387(.a(N1682), .O(gate513inter8));
  nand2 gate2388(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2389(.a(s_215), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2390(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2391(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2392(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );

  xor2  gate1819(.a(N1683), .b(N1734), .O(gate516inter0));
  nand2 gate1820(.a(gate516inter0), .b(s_134), .O(gate516inter1));
  and2  gate1821(.a(N1683), .b(N1734), .O(gate516inter2));
  inv1  gate1822(.a(s_134), .O(gate516inter3));
  inv1  gate1823(.a(s_135), .O(gate516inter4));
  nand2 gate1824(.a(gate516inter4), .b(gate516inter3), .O(gate516inter5));
  nor2  gate1825(.a(gate516inter5), .b(gate516inter2), .O(gate516inter6));
  inv1  gate1826(.a(N1734), .O(gate516inter7));
  inv1  gate1827(.a(N1683), .O(gate516inter8));
  nand2 gate1828(.a(gate516inter8), .b(gate516inter7), .O(gate516inter9));
  nand2 gate1829(.a(s_135), .b(gate516inter3), .O(gate516inter10));
  nor2  gate1830(.a(gate516inter10), .b(gate516inter9), .O(gate516inter11));
  nor2  gate1831(.a(gate516inter11), .b(gate516inter6), .O(gate516inter12));
  nand2 gate1832(.a(gate516inter12), .b(gate516inter1), .O(N1787));
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );

  xor2  gate2127(.a(N1763), .b(N1664), .O(gate519inter0));
  nand2 gate2128(.a(gate519inter0), .b(s_178), .O(gate519inter1));
  and2  gate2129(.a(N1763), .b(N1664), .O(gate519inter2));
  inv1  gate2130(.a(s_178), .O(gate519inter3));
  inv1  gate2131(.a(s_179), .O(gate519inter4));
  nand2 gate2132(.a(gate519inter4), .b(gate519inter3), .O(gate519inter5));
  nor2  gate2133(.a(gate519inter5), .b(gate519inter2), .O(gate519inter6));
  inv1  gate2134(.a(N1664), .O(gate519inter7));
  inv1  gate2135(.a(N1763), .O(gate519inter8));
  nand2 gate2136(.a(gate519inter8), .b(gate519inter7), .O(gate519inter9));
  nand2 gate2137(.a(s_179), .b(gate519inter3), .O(gate519inter10));
  nor2  gate2138(.a(gate519inter10), .b(gate519inter9), .O(gate519inter11));
  nor2  gate2139(.a(gate519inter11), .b(gate519inter6), .O(gate519inter12));
  nand2 gate2140(.a(gate519inter12), .b(gate519inter1), .O(N1792));
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate2239(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate2240(.a(gate522inter0), .b(s_194), .O(gate522inter1));
  and2  gate2241(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate2242(.a(s_194), .O(gate522inter3));
  inv1  gate2243(.a(s_195), .O(gate522inter4));
  nand2 gate2244(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate2245(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate2246(.a(N1740), .O(gate522inter7));
  inv1  gate2247(.a(N1769), .O(gate522inter8));
  nand2 gate2248(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate2249(.a(s_195), .b(gate522inter3), .O(gate522inter10));
  nor2  gate2250(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate2251(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate2252(.a(gate522inter12), .b(gate522inter1), .O(N1798));
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );

  xor2  gate1427(.a(N290), .b(N1742), .O(gate524inter0));
  nand2 gate1428(.a(gate524inter0), .b(s_78), .O(gate524inter1));
  and2  gate1429(.a(N290), .b(N1742), .O(gate524inter2));
  inv1  gate1430(.a(s_78), .O(gate524inter3));
  inv1  gate1431(.a(s_79), .O(gate524inter4));
  nand2 gate1432(.a(gate524inter4), .b(gate524inter3), .O(gate524inter5));
  nor2  gate1433(.a(gate524inter5), .b(gate524inter2), .O(gate524inter6));
  inv1  gate1434(.a(N1742), .O(gate524inter7));
  inv1  gate1435(.a(N290), .O(gate524inter8));
  nand2 gate1436(.a(gate524inter8), .b(gate524inter7), .O(gate524inter9));
  nand2 gate1437(.a(s_79), .b(gate524inter3), .O(gate524inter10));
  nor2  gate1438(.a(gate524inter10), .b(gate524inter9), .O(gate524inter11));
  nor2  gate1439(.a(gate524inter11), .b(gate524inter6), .O(gate524inter12));
  nand2 gate1440(.a(gate524inter12), .b(gate524inter1), .O(N1802));
inv1 gate525( .a(N1748), .O(N1807) );

  xor2  gate2295(.a(N1218), .b(N1748), .O(gate526inter0));
  nand2 gate2296(.a(gate526inter0), .b(s_202), .O(gate526inter1));
  and2  gate2297(.a(N1218), .b(N1748), .O(gate526inter2));
  inv1  gate2298(.a(s_202), .O(gate526inter3));
  inv1  gate2299(.a(s_203), .O(gate526inter4));
  nand2 gate2300(.a(gate526inter4), .b(gate526inter3), .O(gate526inter5));
  nor2  gate2301(.a(gate526inter5), .b(gate526inter2), .O(gate526inter6));
  inv1  gate2302(.a(N1748), .O(gate526inter7));
  inv1  gate2303(.a(N1218), .O(gate526inter8));
  nand2 gate2304(.a(gate526inter8), .b(gate526inter7), .O(gate526inter9));
  nand2 gate2305(.a(s_203), .b(gate526inter3), .O(gate526inter10));
  nor2  gate2306(.a(gate526inter10), .b(gate526inter9), .O(gate526inter11));
  nor2  gate2307(.a(gate526inter11), .b(gate526inter6), .O(gate526inter12));
  nand2 gate2308(.a(gate526inter12), .b(gate526inter1), .O(N1808));
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );

  xor2  gate2197(.a(N1786), .b(N1615), .O(gate528inter0));
  nand2 gate2198(.a(gate528inter0), .b(s_188), .O(gate528inter1));
  and2  gate2199(.a(N1786), .b(N1615), .O(gate528inter2));
  inv1  gate2200(.a(s_188), .O(gate528inter3));
  inv1  gate2201(.a(s_189), .O(gate528inter4));
  nand2 gate2202(.a(gate528inter4), .b(gate528inter3), .O(gate528inter5));
  nor2  gate2203(.a(gate528inter5), .b(gate528inter2), .O(gate528inter6));
  inv1  gate2204(.a(N1615), .O(gate528inter7));
  inv1  gate2205(.a(N1786), .O(gate528inter8));
  nand2 gate2206(.a(gate528inter8), .b(gate528inter7), .O(gate528inter9));
  nand2 gate2207(.a(s_189), .b(gate528inter3), .O(gate528inter10));
  nor2  gate2208(.a(gate528inter10), .b(gate528inter9), .O(gate528inter11));
  nor2  gate2209(.a(gate528inter11), .b(gate528inter6), .O(gate528inter12));
  nand2 gate2210(.a(gate528inter12), .b(gate528inter1), .O(N1810));
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );

  xor2  gate2701(.a(N1764), .b(N1792), .O(gate530inter0));
  nand2 gate2702(.a(gate530inter0), .b(s_260), .O(gate530inter1));
  and2  gate2703(.a(N1764), .b(N1792), .O(gate530inter2));
  inv1  gate2704(.a(s_260), .O(gate530inter3));
  inv1  gate2705(.a(s_261), .O(gate530inter4));
  nand2 gate2706(.a(gate530inter4), .b(gate530inter3), .O(gate530inter5));
  nor2  gate2707(.a(gate530inter5), .b(gate530inter2), .O(gate530inter6));
  inv1  gate2708(.a(N1792), .O(gate530inter7));
  inv1  gate2709(.a(N1764), .O(gate530inter8));
  nand2 gate2710(.a(gate530inter8), .b(gate530inter7), .O(gate530inter9));
  nand2 gate2711(.a(s_261), .b(gate530inter3), .O(gate530inter10));
  nor2  gate2712(.a(gate530inter10), .b(gate530inter9), .O(gate530inter11));
  nor2  gate2713(.a(gate530inter11), .b(gate530inter6), .O(gate530inter12));
  nand2 gate2714(.a(gate530inter12), .b(gate530inter1), .O(N1815));
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate2225(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate2226(.a(gate532inter0), .b(s_192), .O(gate532inter1));
  and2  gate2227(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate2228(.a(s_192), .O(gate532inter3));
  inv1  gate2229(.a(s_193), .O(gate532inter4));
  nand2 gate2230(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate2231(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate2232(.a(N1777), .O(gate532inter7));
  inv1  gate2233(.a(N1490), .O(gate532inter8));
  nand2 gate2234(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate2235(.a(s_193), .b(gate532inter3), .O(gate532inter10));
  nor2  gate2236(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate2237(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate2238(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );

  xor2  gate979(.a(N1801), .b(N1772), .O(gate539inter0));
  nand2 gate980(.a(gate539inter0), .b(s_14), .O(gate539inter1));
  and2  gate981(.a(N1801), .b(N1772), .O(gate539inter2));
  inv1  gate982(.a(s_14), .O(gate539inter3));
  inv1  gate983(.a(s_15), .O(gate539inter4));
  nand2 gate984(.a(gate539inter4), .b(gate539inter3), .O(gate539inter5));
  nor2  gate985(.a(gate539inter5), .b(gate539inter2), .O(gate539inter6));
  inv1  gate986(.a(N1772), .O(gate539inter7));
  inv1  gate987(.a(N1801), .O(gate539inter8));
  nand2 gate988(.a(gate539inter8), .b(gate539inter7), .O(gate539inter9));
  nand2 gate989(.a(s_15), .b(gate539inter3), .O(gate539inter10));
  nor2  gate990(.a(gate539inter10), .b(gate539inter9), .O(gate539inter11));
  nor2  gate991(.a(gate539inter11), .b(gate539inter6), .O(gate539inter12));
  nand2 gate992(.a(gate539inter12), .b(gate539inter1), .O(N1830));

  xor2  gate1203(.a(N1807), .b(N959), .O(gate540inter0));
  nand2 gate1204(.a(gate540inter0), .b(s_46), .O(gate540inter1));
  and2  gate1205(.a(N1807), .b(N959), .O(gate540inter2));
  inv1  gate1206(.a(s_46), .O(gate540inter3));
  inv1  gate1207(.a(s_47), .O(gate540inter4));
  nand2 gate1208(.a(gate540inter4), .b(gate540inter3), .O(gate540inter5));
  nor2  gate1209(.a(gate540inter5), .b(gate540inter2), .O(gate540inter6));
  inv1  gate1210(.a(N959), .O(gate540inter7));
  inv1  gate1211(.a(N1807), .O(gate540inter8));
  nand2 gate1212(.a(gate540inter8), .b(gate540inter7), .O(gate540inter9));
  nand2 gate1213(.a(s_47), .b(gate540inter3), .O(gate540inter10));
  nor2  gate1214(.a(gate540inter10), .b(gate540inter9), .O(gate540inter11));
  nor2  gate1215(.a(gate540inter11), .b(gate540inter6), .O(gate540inter12));
  nand2 gate1216(.a(gate540inter12), .b(gate540inter1), .O(N1837));

  xor2  gate1707(.a(N1784), .b(N1809), .O(gate541inter0));
  nand2 gate1708(.a(gate541inter0), .b(s_118), .O(gate541inter1));
  and2  gate1709(.a(N1784), .b(N1809), .O(gate541inter2));
  inv1  gate1710(.a(s_118), .O(gate541inter3));
  inv1  gate1711(.a(s_119), .O(gate541inter4));
  nand2 gate1712(.a(gate541inter4), .b(gate541inter3), .O(gate541inter5));
  nor2  gate1713(.a(gate541inter5), .b(gate541inter2), .O(gate541inter6));
  inv1  gate1714(.a(N1809), .O(gate541inter7));
  inv1  gate1715(.a(N1784), .O(gate541inter8));
  nand2 gate1716(.a(gate541inter8), .b(gate541inter7), .O(gate541inter9));
  nand2 gate1717(.a(s_119), .b(gate541inter3), .O(gate541inter10));
  nor2  gate1718(.a(gate541inter10), .b(gate541inter9), .O(gate541inter11));
  nor2  gate1719(.a(gate541inter11), .b(gate541inter6), .O(gate541inter12));
  nand2 gate1720(.a(gate541inter12), .b(gate541inter1), .O(N1838));
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );

  xor2  gate1861(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate1862(.a(gate544inter0), .b(s_140), .O(gate544inter1));
  and2  gate1863(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate1864(.a(s_140), .O(gate544inter3));
  inv1  gate1865(.a(s_141), .O(gate544inter4));
  nand2 gate1866(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate1867(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate1868(.a(N1416), .O(gate544inter7));
  inv1  gate1869(.a(N1824), .O(gate544inter8));
  nand2 gate1870(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate1871(.a(s_141), .b(gate544inter3), .O(gate544inter10));
  nor2  gate1872(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate1873(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate1874(.a(gate544inter12), .b(gate544inter1), .O(N1849));
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );

  xor2  gate2309(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate2310(.a(gate546inter0), .b(s_204), .O(gate546inter1));
  and2  gate2311(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate2312(.a(s_204), .O(gate546inter3));
  inv1  gate2313(.a(s_205), .O(gate546inter4));
  nand2 gate2314(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate2315(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate2316(.a(N1319), .O(gate546inter7));
  inv1  gate2317(.a(N1827), .O(gate546inter8));
  nand2 gate2318(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate2319(.a(s_205), .b(gate546inter3), .O(gate546inter10));
  nor2  gate2320(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate2321(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate2322(.a(gate546inter12), .b(gate546inter1), .O(N1852));
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );

  xor2  gate937(.a(N1837), .b(N1808), .O(gate556inter0));
  nand2 gate938(.a(gate556inter0), .b(s_8), .O(gate556inter1));
  and2  gate939(.a(N1837), .b(N1808), .O(gate556inter2));
  inv1  gate940(.a(s_8), .O(gate556inter3));
  inv1  gate941(.a(s_9), .O(gate556inter4));
  nand2 gate942(.a(gate556inter4), .b(gate556inter3), .O(gate556inter5));
  nor2  gate943(.a(gate556inter5), .b(gate556inter2), .O(gate556inter6));
  inv1  gate944(.a(N1808), .O(gate556inter7));
  inv1  gate945(.a(N1837), .O(gate556inter8));
  nand2 gate946(.a(gate556inter8), .b(gate556inter7), .O(gate556inter9));
  nand2 gate947(.a(s_9), .b(gate556inter3), .O(gate556inter10));
  nor2  gate948(.a(gate556inter10), .b(gate556inter9), .O(gate556inter11));
  nor2  gate949(.a(gate556inter11), .b(gate556inter6), .O(gate556inter12));
  nand2 gate950(.a(gate556inter12), .b(gate556inter1), .O(N1875));
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );

  xor2  gate2841(.a(N1768), .b(N1841), .O(gate559inter0));
  nand2 gate2842(.a(gate559inter0), .b(s_280), .O(gate559inter1));
  and2  gate2843(.a(N1768), .b(N1841), .O(gate559inter2));
  inv1  gate2844(.a(s_280), .O(gate559inter3));
  inv1  gate2845(.a(s_281), .O(gate559inter4));
  nand2 gate2846(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate2847(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate2848(.a(N1841), .O(gate559inter7));
  inv1  gate2849(.a(N1768), .O(gate559inter8));
  nand2 gate2850(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate2851(.a(s_281), .b(gate559inter3), .O(gate559inter10));
  nor2  gate2852(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate2853(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate2854(.a(gate559inter12), .b(gate559inter1), .O(N1882));
inv1 gate560( .a(N1841), .O(N1883) );

  xor2  gate1021(.a(N1852), .b(N1826), .O(gate561inter0));
  nand2 gate1022(.a(gate561inter0), .b(s_20), .O(gate561inter1));
  and2  gate1023(.a(N1852), .b(N1826), .O(gate561inter2));
  inv1  gate1024(.a(s_20), .O(gate561inter3));
  inv1  gate1025(.a(s_21), .O(gate561inter4));
  nand2 gate1026(.a(gate561inter4), .b(gate561inter3), .O(gate561inter5));
  nor2  gate1027(.a(gate561inter5), .b(gate561inter2), .O(gate561inter6));
  inv1  gate1028(.a(N1826), .O(gate561inter7));
  inv1  gate1029(.a(N1852), .O(gate561inter8));
  nand2 gate1030(.a(gate561inter8), .b(gate561inter7), .O(gate561inter9));
  nand2 gate1031(.a(s_21), .b(gate561inter3), .O(gate561inter10));
  nor2  gate1032(.a(gate561inter10), .b(gate561inter9), .O(gate561inter11));
  nor2  gate1033(.a(gate561inter11), .b(gate561inter6), .O(gate561inter12));
  nand2 gate1034(.a(gate561inter12), .b(gate561inter1), .O(N1884));
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );

  xor2  gate1007(.a(N1883), .b(N1717), .O(gate570inter0));
  nand2 gate1008(.a(gate570inter0), .b(s_18), .O(gate570inter1));
  and2  gate1009(.a(N1883), .b(N1717), .O(gate570inter2));
  inv1  gate1010(.a(s_18), .O(gate570inter3));
  inv1  gate1011(.a(s_19), .O(gate570inter4));
  nand2 gate1012(.a(gate570inter4), .b(gate570inter3), .O(gate570inter5));
  nor2  gate1013(.a(gate570inter5), .b(gate570inter2), .O(gate570inter6));
  inv1  gate1014(.a(N1717), .O(gate570inter7));
  inv1  gate1015(.a(N1883), .O(gate570inter8));
  nand2 gate1016(.a(gate570inter8), .b(gate570inter7), .O(gate570inter9));
  nand2 gate1017(.a(s_19), .b(gate570inter3), .O(gate570inter10));
  nor2  gate1018(.a(gate570inter10), .b(gate570inter9), .O(gate570inter11));
  nor2  gate1019(.a(gate570inter11), .b(gate570inter6), .O(gate570inter12));
  nand2 gate1020(.a(gate570inter12), .b(gate570inter1), .O(N1911));
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate2449(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate2450(.a(gate574inter0), .b(s_224), .O(gate574inter1));
  and2  gate2451(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate2452(.a(s_224), .O(gate574inter3));
  inv1  gate2453(.a(s_225), .O(gate574inter4));
  nand2 gate2454(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate2455(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate2456(.a(N1872), .O(gate574inter7));
  inv1  gate2457(.a(N919), .O(gate574inter8));
  nand2 gate2458(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate2459(.a(s_225), .b(gate574inter3), .O(gate574inter10));
  nor2  gate2460(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate2461(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate2462(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );

  xor2  gate2547(.a(N920), .b(N1869), .O(gate576inter0));
  nand2 gate2548(.a(gate576inter0), .b(s_238), .O(gate576inter1));
  and2  gate2549(.a(N920), .b(N1869), .O(gate576inter2));
  inv1  gate2550(.a(s_238), .O(gate576inter3));
  inv1  gate2551(.a(s_239), .O(gate576inter4));
  nand2 gate2552(.a(gate576inter4), .b(gate576inter3), .O(gate576inter5));
  nor2  gate2553(.a(gate576inter5), .b(gate576inter2), .O(gate576inter6));
  inv1  gate2554(.a(N1869), .O(gate576inter7));
  inv1  gate2555(.a(N920), .O(gate576inter8));
  nand2 gate2556(.a(gate576inter8), .b(gate576inter7), .O(gate576inter9));
  nand2 gate2557(.a(s_239), .b(gate576inter3), .O(gate576inter10));
  nor2  gate2558(.a(gate576inter10), .b(gate576inter9), .O(gate576inter11));
  nor2  gate2559(.a(gate576inter11), .b(gate576inter6), .O(gate576inter12));
  nand2 gate2560(.a(gate576inter12), .b(gate576inter1), .O(N1921));
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );

  xor2  gate1959(.a(N1920), .b(N679), .O(gate586inter0));
  nand2 gate1960(.a(gate586inter0), .b(s_154), .O(gate586inter1));
  and2  gate1961(.a(N1920), .b(N679), .O(gate586inter2));
  inv1  gate1962(.a(s_154), .O(gate586inter3));
  inv1  gate1963(.a(s_155), .O(gate586inter4));
  nand2 gate1964(.a(gate586inter4), .b(gate586inter3), .O(gate586inter5));
  nor2  gate1965(.a(gate586inter5), .b(gate586inter2), .O(gate586inter6));
  inv1  gate1966(.a(N679), .O(gate586inter7));
  inv1  gate1967(.a(N1920), .O(gate586inter8));
  nand2 gate1968(.a(gate586inter8), .b(gate586inter7), .O(gate586inter9));
  nand2 gate1969(.a(s_155), .b(gate586inter3), .O(gate586inter10));
  nor2  gate1970(.a(gate586inter10), .b(gate586inter9), .O(gate586inter11));
  nor2  gate1971(.a(gate586inter11), .b(gate586inter6), .O(gate586inter12));
  nand2 gate1972(.a(gate586inter12), .b(gate586inter1), .O(N1941));

  xor2  gate1805(.a(N1922), .b(N676), .O(gate587inter0));
  nand2 gate1806(.a(gate587inter0), .b(s_132), .O(gate587inter1));
  and2  gate1807(.a(N1922), .b(N676), .O(gate587inter2));
  inv1  gate1808(.a(s_132), .O(gate587inter3));
  inv1  gate1809(.a(s_133), .O(gate587inter4));
  nand2 gate1810(.a(gate587inter4), .b(gate587inter3), .O(gate587inter5));
  nor2  gate1811(.a(gate587inter5), .b(gate587inter2), .O(gate587inter6));
  inv1  gate1812(.a(N676), .O(gate587inter7));
  inv1  gate1813(.a(N1922), .O(gate587inter8));
  nand2 gate1814(.a(gate587inter8), .b(gate587inter7), .O(gate587inter9));
  nand2 gate1815(.a(s_133), .b(gate587inter3), .O(gate587inter10));
  nor2  gate1816(.a(gate587inter10), .b(gate587inter9), .O(gate587inter11));
  nor2  gate1817(.a(gate587inter11), .b(gate587inter6), .O(gate587inter12));
  nand2 gate1818(.a(gate587inter12), .b(gate587inter1), .O(N1942));
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );

  xor2  gate2757(.a(N1941), .b(N1919), .O(gate600inter0));
  nand2 gate2758(.a(gate600inter0), .b(s_268), .O(gate600inter1));
  and2  gate2759(.a(N1941), .b(N1919), .O(gate600inter2));
  inv1  gate2760(.a(s_268), .O(gate600inter3));
  inv1  gate2761(.a(s_269), .O(gate600inter4));
  nand2 gate2762(.a(gate600inter4), .b(gate600inter3), .O(gate600inter5));
  nor2  gate2763(.a(gate600inter5), .b(gate600inter2), .O(gate600inter6));
  inv1  gate2764(.a(N1919), .O(gate600inter7));
  inv1  gate2765(.a(N1941), .O(gate600inter8));
  nand2 gate2766(.a(gate600inter8), .b(gate600inter7), .O(gate600inter9));
  nand2 gate2767(.a(s_269), .b(gate600inter3), .O(gate600inter10));
  nor2  gate2768(.a(gate600inter10), .b(gate600inter9), .O(gate600inter11));
  nor2  gate2769(.a(gate600inter11), .b(gate600inter6), .O(gate600inter12));
  nand2 gate2770(.a(gate600inter12), .b(gate600inter1), .O(N1979));

  xor2  gate1889(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate1890(.a(gate601inter0), .b(s_144), .O(gate601inter1));
  and2  gate1891(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate1892(.a(s_144), .O(gate601inter3));
  inv1  gate1893(.a(s_145), .O(gate601inter4));
  nand2 gate1894(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate1895(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate1896(.a(N1921), .O(gate601inter7));
  inv1  gate1897(.a(N1942), .O(gate601inter8));
  nand2 gate1898(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate1899(.a(s_145), .b(gate601inter3), .O(gate601inter10));
  nor2  gate1900(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate1901(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate1902(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );

  xor2  gate2785(.a(N1937), .b(N1944), .O(gate605inter0));
  nand2 gate2786(.a(gate605inter0), .b(s_272), .O(gate605inter1));
  and2  gate2787(.a(N1937), .b(N1944), .O(gate605inter2));
  inv1  gate2788(.a(s_272), .O(gate605inter3));
  inv1  gate2789(.a(s_273), .O(gate605inter4));
  nand2 gate2790(.a(gate605inter4), .b(gate605inter3), .O(gate605inter5));
  nor2  gate2791(.a(gate605inter5), .b(gate605inter2), .O(gate605inter6));
  inv1  gate2792(.a(N1944), .O(gate605inter7));
  inv1  gate2793(.a(N1937), .O(gate605inter8));
  nand2 gate2794(.a(gate605inter8), .b(gate605inter7), .O(gate605inter9));
  nand2 gate2795(.a(s_273), .b(gate605inter3), .O(gate605inter10));
  nor2  gate2796(.a(gate605inter10), .b(gate605inter9), .O(gate605inter11));
  nor2  gate2797(.a(gate605inter11), .b(gate605inter6), .O(gate605inter12));
  nand2 gate2798(.a(gate605inter12), .b(gate605inter1), .O(N2000));
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );

  xor2  gate1063(.a(N1350), .b(N1953), .O(gate608inter0));
  nand2 gate1064(.a(gate608inter0), .b(s_26), .O(gate608inter1));
  and2  gate1065(.a(N1350), .b(N1953), .O(gate608inter2));
  inv1  gate1066(.a(s_26), .O(gate608inter3));
  inv1  gate1067(.a(s_27), .O(gate608inter4));
  nand2 gate1068(.a(gate608inter4), .b(gate608inter3), .O(gate608inter5));
  nor2  gate1069(.a(gate608inter5), .b(gate608inter2), .O(gate608inter6));
  inv1  gate1070(.a(N1953), .O(gate608inter7));
  inv1  gate1071(.a(N1350), .O(gate608inter8));
  nand2 gate1072(.a(gate608inter8), .b(gate608inter7), .O(gate608inter9));
  nand2 gate1073(.a(s_27), .b(gate608inter3), .O(gate608inter10));
  nor2  gate1074(.a(gate608inter10), .b(gate608inter9), .O(gate608inter11));
  nor2  gate1075(.a(gate608inter11), .b(gate608inter6), .O(gate608inter12));
  nand2 gate1076(.a(gate608inter12), .b(gate608inter1), .O(N2004));
inv1 gate609( .a(N1953), .O(N2005) );

  xor2  gate1693(.a(N1351), .b(N1950), .O(gate610inter0));
  nand2 gate1694(.a(gate610inter0), .b(s_116), .O(gate610inter1));
  and2  gate1695(.a(N1351), .b(N1950), .O(gate610inter2));
  inv1  gate1696(.a(s_116), .O(gate610inter3));
  inv1  gate1697(.a(s_117), .O(gate610inter4));
  nand2 gate1698(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate1699(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate1700(.a(N1950), .O(gate610inter7));
  inv1  gate1701(.a(N1351), .O(gate610inter8));
  nand2 gate1702(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate1703(.a(s_117), .b(gate610inter3), .O(gate610inter10));
  nor2  gate1704(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate1705(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate1706(.a(gate610inter12), .b(gate610inter1), .O(N2006));
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate1441(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate1442(.a(gate612inter0), .b(s_80), .O(gate612inter1));
  and2  gate1443(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate1444(.a(s_80), .O(gate612inter3));
  inv1  gate1445(.a(s_81), .O(gate612inter4));
  nand2 gate1446(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate1447(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate1448(.a(N673), .O(gate612inter7));
  inv1  gate1449(.a(N1976), .O(gate612inter8));
  nand2 gate1450(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate1451(.a(s_81), .b(gate612inter3), .O(gate612inter10));
  nor2  gate1452(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate1453(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate1454(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );

  xor2  gate1259(.a(N1923), .b(N1958), .O(gate616inter0));
  nand2 gate1260(.a(gate616inter0), .b(s_54), .O(gate616inter1));
  and2  gate1261(.a(N1923), .b(N1958), .O(gate616inter2));
  inv1  gate1262(.a(s_54), .O(gate616inter3));
  inv1  gate1263(.a(s_55), .O(gate616inter4));
  nand2 gate1264(.a(gate616inter4), .b(gate616inter3), .O(gate616inter5));
  nor2  gate1265(.a(gate616inter5), .b(gate616inter2), .O(gate616inter6));
  inv1  gate1266(.a(N1958), .O(gate616inter7));
  inv1  gate1267(.a(N1923), .O(gate616inter8));
  nand2 gate1268(.a(gate616inter8), .b(gate616inter7), .O(gate616inter9));
  nand2 gate1269(.a(s_55), .b(gate616inter3), .O(gate616inter10));
  nor2  gate1270(.a(gate616inter10), .b(gate616inter9), .O(gate616inter11));
  nor2  gate1271(.a(gate616inter11), .b(gate616inter6), .O(gate616inter12));
  nand2 gate1272(.a(gate616inter12), .b(gate616inter1), .O(N2014));
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );

  xor2  gate1455(.a(N2007), .b(N1258), .O(gate626inter0));
  nand2 gate1456(.a(gate626inter0), .b(s_82), .O(gate626inter1));
  and2  gate1457(.a(N2007), .b(N1258), .O(gate626inter2));
  inv1  gate1458(.a(s_82), .O(gate626inter3));
  inv1  gate1459(.a(s_83), .O(gate626inter4));
  nand2 gate1460(.a(gate626inter4), .b(gate626inter3), .O(gate626inter5));
  nor2  gate1461(.a(gate626inter5), .b(gate626inter2), .O(gate626inter6));
  inv1  gate1462(.a(N1258), .O(gate626inter7));
  inv1  gate1463(.a(N2007), .O(gate626inter8));
  nand2 gate1464(.a(gate626inter8), .b(gate626inter7), .O(gate626inter9));
  nand2 gate1465(.a(s_83), .b(gate626inter3), .O(gate626inter10));
  nor2  gate1466(.a(gate626inter10), .b(gate626inter9), .O(gate626inter11));
  nor2  gate1467(.a(gate626inter11), .b(gate626inter6), .O(gate626inter12));
  nand2 gate1468(.a(gate626inter12), .b(gate626inter1), .O(N2025));

  xor2  gate1119(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate1120(.a(gate627inter0), .b(s_34), .O(gate627inter1));
  and2  gate1121(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate1122(.a(s_34), .O(gate627inter3));
  inv1  gate1123(.a(s_35), .O(gate627inter4));
  nand2 gate1124(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate1125(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate1126(.a(N1975), .O(gate627inter7));
  inv1  gate1127(.a(N2008), .O(gate627inter8));
  nand2 gate1128(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate1129(.a(s_35), .b(gate627inter3), .O(gate627inter10));
  nor2  gate1130(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate1131(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate1132(.a(gate627inter12), .b(gate627inter1), .O(N2026));
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate2589(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate2590(.a(gate633inter0), .b(s_244), .O(gate633inter1));
  and2  gate2591(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate2592(.a(s_244), .O(gate633inter3));
  inv1  gate2593(.a(s_245), .O(gate633inter4));
  nand2 gate2594(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate2595(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate2596(.a(N2020), .O(gate633inter7));
  inv1  gate2597(.a(N2000), .O(gate633inter8));
  nand2 gate2598(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate2599(.a(s_245), .b(gate633inter3), .O(gate633inter10));
  nor2  gate2600(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate2601(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate2602(.a(gate633inter12), .b(gate633inter1), .O(N2038));

  xor2  gate2211(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate2212(.a(gate634inter0), .b(s_190), .O(gate634inter1));
  and2  gate2213(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate2214(.a(s_190), .O(gate634inter3));
  inv1  gate2215(.a(s_191), .O(gate634inter4));
  nand2 gate2216(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate2217(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate2218(.a(N1534), .O(gate634inter7));
  inv1  gate2219(.a(N2021), .O(gate634inter8));
  nand2 gate2220(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate2221(.a(s_191), .b(gate634inter3), .O(gate634inter10));
  nor2  gate2222(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate2223(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate2224(.a(gate634inter12), .b(gate634inter1), .O(N2039));
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );

  xor2  gate1077(.a(N290), .b(N2061), .O(gate650inter0));
  nand2 gate1078(.a(gate650inter0), .b(s_28), .O(gate650inter1));
  and2  gate1079(.a(N290), .b(N2061), .O(gate650inter2));
  inv1  gate1080(.a(s_28), .O(gate650inter3));
  inv1  gate1081(.a(s_29), .O(gate650inter4));
  nand2 gate1082(.a(gate650inter4), .b(gate650inter3), .O(gate650inter5));
  nor2  gate1083(.a(gate650inter5), .b(gate650inter2), .O(gate650inter6));
  inv1  gate1084(.a(N2061), .O(gate650inter7));
  inv1  gate1085(.a(N290), .O(gate650inter8));
  nand2 gate1086(.a(gate650inter8), .b(gate650inter7), .O(gate650inter9));
  nand2 gate1087(.a(s_29), .b(gate650inter3), .O(gate650inter10));
  nor2  gate1088(.a(gate650inter10), .b(gate650inter9), .O(gate650inter11));
  nor2  gate1089(.a(gate650inter11), .b(gate650inter6), .O(gate650inter12));
  nand2 gate1090(.a(gate650inter12), .b(gate650inter1), .O(N2081));
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate2421(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate2422(.a(gate667inter0), .b(s_220), .O(gate667inter1));
  and2  gate2423(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate2424(.a(s_220), .O(gate667inter3));
  inv1  gate2425(.a(s_221), .O(gate667inter4));
  nand2 gate2426(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate2427(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate2428(.a(N2199), .O(gate667inter7));
  inv1  gate2429(.a(N1348), .O(gate667inter8));
  nand2 gate2430(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate2431(.a(s_221), .b(gate667inter3), .O(gate667inter10));
  nor2  gate2432(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate2433(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate2434(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate1791(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate1792(.a(gate671inter0), .b(s_130), .O(gate671inter1));
  and2  gate1793(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate1794(.a(s_130), .O(gate671inter3));
  inv1  gate1795(.a(s_131), .O(gate671inter4));
  nand2 gate1796(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate1797(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate1798(.a(N2205), .O(gate671inter7));
  inv1  gate1799(.a(N913), .O(gate671inter8));
  nand2 gate1800(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate1801(.a(s_131), .b(gate671inter3), .O(gate671inter10));
  nor2  gate1802(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate1803(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate1804(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );

  xor2  gate2015(.a(N2223), .b(N1255), .O(gate677inter0));
  nand2 gate2016(.a(gate677inter0), .b(s_162), .O(gate677inter1));
  and2  gate2017(.a(N2223), .b(N1255), .O(gate677inter2));
  inv1  gate2018(.a(s_162), .O(gate677inter3));
  inv1  gate2019(.a(s_163), .O(gate677inter4));
  nand2 gate2020(.a(gate677inter4), .b(gate677inter3), .O(gate677inter5));
  nor2  gate2021(.a(gate677inter5), .b(gate677inter2), .O(gate677inter6));
  inv1  gate2022(.a(N1255), .O(gate677inter7));
  inv1  gate2023(.a(N2223), .O(gate677inter8));
  nand2 gate2024(.a(gate677inter8), .b(gate677inter7), .O(gate677inter9));
  nand2 gate2025(.a(s_163), .b(gate677inter3), .O(gate677inter10));
  nor2  gate2026(.a(gate677inter10), .b(gate677inter9), .O(gate677inter11));
  nor2  gate2027(.a(gate677inter11), .b(gate677inter6), .O(gate677inter12));
  nand2 gate2028(.a(gate677inter12), .b(gate677inter1), .O(N2232));

  xor2  gate2687(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate2688(.a(gate678inter0), .b(s_258), .O(gate678inter1));
  and2  gate2689(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate2690(.a(s_258), .O(gate678inter3));
  inv1  gate2691(.a(s_259), .O(gate678inter4));
  nand2 gate2692(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate2693(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate2694(.a(N1252), .O(gate678inter7));
  inv1  gate2695(.a(N2225), .O(gate678inter8));
  nand2 gate2696(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate2697(.a(s_259), .b(gate678inter3), .O(gate678inter10));
  nor2  gate2698(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate2699(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate2700(.a(gate678inter12), .b(gate678inter1), .O(N2233));
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );

  xor2  gate1917(.a(N2231), .b(N2216), .O(gate682inter0));
  nand2 gate1918(.a(gate682inter0), .b(s_148), .O(gate682inter1));
  and2  gate1919(.a(N2231), .b(N2216), .O(gate682inter2));
  inv1  gate1920(.a(s_148), .O(gate682inter3));
  inv1  gate1921(.a(s_149), .O(gate682inter4));
  nand2 gate1922(.a(gate682inter4), .b(gate682inter3), .O(gate682inter5));
  nor2  gate1923(.a(gate682inter5), .b(gate682inter2), .O(gate682inter6));
  inv1  gate1924(.a(N2216), .O(gate682inter7));
  inv1  gate1925(.a(N2231), .O(gate682inter8));
  nand2 gate1926(.a(gate682inter8), .b(gate682inter7), .O(gate682inter9));
  nand2 gate1927(.a(s_149), .b(gate682inter3), .O(gate682inter10));
  nor2  gate1928(.a(gate682inter10), .b(gate682inter9), .O(gate682inter11));
  nor2  gate1929(.a(gate682inter11), .b(gate682inter6), .O(gate682inter12));
  nand2 gate1930(.a(gate682inter12), .b(gate682inter1), .O(N2237));

  xor2  gate2575(.a(N2232), .b(N2222), .O(gate683inter0));
  nand2 gate2576(.a(gate683inter0), .b(s_242), .O(gate683inter1));
  and2  gate2577(.a(N2232), .b(N2222), .O(gate683inter2));
  inv1  gate2578(.a(s_242), .O(gate683inter3));
  inv1  gate2579(.a(s_243), .O(gate683inter4));
  nand2 gate2580(.a(gate683inter4), .b(gate683inter3), .O(gate683inter5));
  nor2  gate2581(.a(gate683inter5), .b(gate683inter2), .O(gate683inter6));
  inv1  gate2582(.a(N2222), .O(gate683inter7));
  inv1  gate2583(.a(N2232), .O(gate683inter8));
  nand2 gate2584(.a(gate683inter8), .b(gate683inter7), .O(gate683inter9));
  nand2 gate2585(.a(s_243), .b(gate683inter3), .O(gate683inter10));
  nor2  gate2586(.a(gate683inter10), .b(gate683inter9), .O(gate683inter11));
  nor2  gate2587(.a(gate683inter11), .b(gate683inter6), .O(gate683inter12));
  nand2 gate2588(.a(gate683inter12), .b(gate683inter1), .O(N2240));
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate1679(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate1680(.a(gate754inter0), .b(s_114), .O(gate754inter1));
  and2  gate1681(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate1682(.a(s_114), .O(gate754inter3));
  inv1  gate1683(.a(s_115), .O(gate754inter4));
  nand2 gate1684(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1685(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1686(.a(N2564), .O(gate754inter7));
  inv1  gate1687(.a(N536), .O(gate754inter8));
  nand2 gate1688(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1689(.a(s_115), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1690(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1691(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1692(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );

  xor2  gate1245(.a(N543), .b(N2570), .O(gate758inter0));
  nand2 gate1246(.a(gate758inter0), .b(s_52), .O(gate758inter1));
  and2  gate1247(.a(N543), .b(N2570), .O(gate758inter2));
  inv1  gate1248(.a(s_52), .O(gate758inter3));
  inv1  gate1249(.a(s_53), .O(gate758inter4));
  nand2 gate1250(.a(gate758inter4), .b(gate758inter3), .O(gate758inter5));
  nor2  gate1251(.a(gate758inter5), .b(gate758inter2), .O(gate758inter6));
  inv1  gate1252(.a(N2570), .O(gate758inter7));
  inv1  gate1253(.a(N543), .O(gate758inter8));
  nand2 gate1254(.a(gate758inter8), .b(gate758inter7), .O(gate758inter9));
  nand2 gate1255(.a(s_53), .b(gate758inter3), .O(gate758inter10));
  nor2  gate1256(.a(gate758inter10), .b(gate758inter9), .O(gate758inter11));
  nor2  gate1257(.a(gate758inter11), .b(gate758inter6), .O(gate758inter12));
  nand2 gate1258(.a(gate758inter12), .b(gate758inter1), .O(N2682));
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );

  xor2  gate1217(.a(N2670), .b(N343), .O(gate765inter0));
  nand2 gate1218(.a(gate765inter0), .b(s_48), .O(gate765inter1));
  and2  gate1219(.a(N2670), .b(N343), .O(gate765inter2));
  inv1  gate1220(.a(s_48), .O(gate765inter3));
  inv1  gate1221(.a(s_49), .O(gate765inter4));
  nand2 gate1222(.a(gate765inter4), .b(gate765inter3), .O(gate765inter5));
  nor2  gate1223(.a(gate765inter5), .b(gate765inter2), .O(gate765inter6));
  inv1  gate1224(.a(N343), .O(gate765inter7));
  inv1  gate1225(.a(N2670), .O(gate765inter8));
  nand2 gate1226(.a(gate765inter8), .b(gate765inter7), .O(gate765inter9));
  nand2 gate1227(.a(s_49), .b(gate765inter3), .O(gate765inter10));
  nor2  gate1228(.a(gate765inter10), .b(gate765inter9), .O(gate765inter11));
  nor2  gate1229(.a(gate765inter11), .b(gate765inter6), .O(gate765inter12));
  nand2 gate1230(.a(gate765inter12), .b(gate765inter1), .O(N2720));
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );

  xor2  gate2519(.a(N538), .b(N2639), .O(gate769inter0));
  nand2 gate2520(.a(gate769inter0), .b(s_234), .O(gate769inter1));
  and2  gate2521(.a(N538), .b(N2639), .O(gate769inter2));
  inv1  gate2522(.a(s_234), .O(gate769inter3));
  inv1  gate2523(.a(s_235), .O(gate769inter4));
  nand2 gate2524(.a(gate769inter4), .b(gate769inter3), .O(gate769inter5));
  nor2  gate2525(.a(gate769inter5), .b(gate769inter2), .O(gate769inter6));
  inv1  gate2526(.a(N2639), .O(gate769inter7));
  inv1  gate2527(.a(N538), .O(gate769inter8));
  nand2 gate2528(.a(gate769inter8), .b(gate769inter7), .O(gate769inter9));
  nand2 gate2529(.a(s_235), .b(gate769inter3), .O(gate769inter10));
  nor2  gate2530(.a(gate769inter10), .b(gate769inter9), .O(gate769inter11));
  nor2  gate2531(.a(gate769inter11), .b(gate769inter6), .O(gate769inter12));
  nand2 gate2532(.a(gate769inter12), .b(gate769inter1), .O(N2724));
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate1161(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate1162(.a(gate773inter0), .b(s_40), .O(gate773inter1));
  and2  gate1163(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate1164(.a(s_40), .O(gate773inter3));
  inv1  gate1165(.a(s_41), .O(gate773inter4));
  nand2 gate1166(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate1167(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate1168(.a(N2645), .O(gate773inter7));
  inv1  gate1169(.a(N540), .O(gate773inter8));
  nand2 gate1170(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate1171(.a(s_41), .b(gate773inter3), .O(gate773inter10));
  nor2  gate1172(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate1173(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate1174(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );

  xor2  gate1847(.a(N542), .b(N2651), .O(gate777inter0));
  nand2 gate1848(.a(gate777inter0), .b(s_138), .O(gate777inter1));
  and2  gate1849(.a(N542), .b(N2651), .O(gate777inter2));
  inv1  gate1850(.a(s_138), .O(gate777inter3));
  inv1  gate1851(.a(s_139), .O(gate777inter4));
  nand2 gate1852(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate1853(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate1854(.a(N2651), .O(gate777inter7));
  inv1  gate1855(.a(N542), .O(gate777inter8));
  nand2 gate1856(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate1857(.a(s_139), .b(gate777inter3), .O(gate777inter10));
  nor2  gate1858(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate1859(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate1860(.a(gate777inter12), .b(gate777inter1), .O(N2732));
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );

  xor2  gate1623(.a(N546), .b(N2661), .O(gate784inter0));
  nand2 gate1624(.a(gate784inter0), .b(s_106), .O(gate784inter1));
  and2  gate1625(.a(N546), .b(N2661), .O(gate784inter2));
  inv1  gate1626(.a(s_106), .O(gate784inter3));
  inv1  gate1627(.a(s_107), .O(gate784inter4));
  nand2 gate1628(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate1629(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate1630(.a(N2661), .O(gate784inter7));
  inv1  gate1631(.a(N546), .O(gate784inter8));
  nand2 gate1632(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate1633(.a(s_107), .b(gate784inter3), .O(gate784inter10));
  nor2  gate1634(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate1635(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate1636(.a(gate784inter12), .b(gate784inter1), .O(N2739));
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );

  xor2  gate2393(.a(N2720), .b(N2669), .O(gate794inter0));
  nand2 gate2394(.a(gate794inter0), .b(s_216), .O(gate794inter1));
  and2  gate2395(.a(N2720), .b(N2669), .O(gate794inter2));
  inv1  gate2396(.a(s_216), .O(gate794inter3));
  inv1  gate2397(.a(s_217), .O(gate794inter4));
  nand2 gate2398(.a(gate794inter4), .b(gate794inter3), .O(gate794inter5));
  nor2  gate2399(.a(gate794inter5), .b(gate794inter2), .O(gate794inter6));
  inv1  gate2400(.a(N2669), .O(gate794inter7));
  inv1  gate2401(.a(N2720), .O(gate794inter8));
  nand2 gate2402(.a(gate794inter8), .b(gate794inter7), .O(gate794inter9));
  nand2 gate2403(.a(s_217), .b(gate794inter3), .O(gate794inter10));
  nor2  gate2404(.a(gate794inter10), .b(gate794inter9), .O(gate794inter11));
  nor2  gate2405(.a(gate794inter11), .b(gate794inter6), .O(gate794inter12));
  nand2 gate2406(.a(gate794inter12), .b(gate794inter1), .O(N2753));
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );

  xor2  gate1483(.a(N2723), .b(N2675), .O(gate797inter0));
  nand2 gate1484(.a(gate797inter0), .b(s_86), .O(gate797inter1));
  and2  gate1485(.a(N2723), .b(N2675), .O(gate797inter2));
  inv1  gate1486(.a(s_86), .O(gate797inter3));
  inv1  gate1487(.a(s_87), .O(gate797inter4));
  nand2 gate1488(.a(gate797inter4), .b(gate797inter3), .O(gate797inter5));
  nor2  gate1489(.a(gate797inter5), .b(gate797inter2), .O(gate797inter6));
  inv1  gate1490(.a(N2675), .O(gate797inter7));
  inv1  gate1491(.a(N2723), .O(gate797inter8));
  nand2 gate1492(.a(gate797inter8), .b(gate797inter7), .O(gate797inter9));
  nand2 gate1493(.a(s_87), .b(gate797inter3), .O(gate797inter10));
  nor2  gate1494(.a(gate797inter10), .b(gate797inter9), .O(gate797inter11));
  nor2  gate1495(.a(gate797inter11), .b(gate797inter6), .O(gate797inter12));
  nand2 gate1496(.a(gate797inter12), .b(gate797inter1), .O(N2756));
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );

  xor2  gate1833(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate1834(.a(gate799inter0), .b(s_136), .O(gate799inter1));
  and2  gate1835(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate1836(.a(s_136), .O(gate799inter3));
  inv1  gate1837(.a(s_137), .O(gate799inter4));
  nand2 gate1838(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate1839(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate1840(.a(N358), .O(gate799inter7));
  inv1  gate1841(.a(N2727), .O(gate799inter8));
  nand2 gate1842(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate1843(.a(s_137), .b(gate799inter3), .O(gate799inter10));
  nor2  gate1844(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate1845(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate1846(.a(gate799inter12), .b(gate799inter1), .O(N2758));

  xor2  gate1287(.a(N2729), .b(N361), .O(gate800inter0));
  nand2 gate1288(.a(gate800inter0), .b(s_58), .O(gate800inter1));
  and2  gate1289(.a(N2729), .b(N361), .O(gate800inter2));
  inv1  gate1290(.a(s_58), .O(gate800inter3));
  inv1  gate1291(.a(s_59), .O(gate800inter4));
  nand2 gate1292(.a(gate800inter4), .b(gate800inter3), .O(gate800inter5));
  nor2  gate1293(.a(gate800inter5), .b(gate800inter2), .O(gate800inter6));
  inv1  gate1294(.a(N361), .O(gate800inter7));
  inv1  gate1295(.a(N2729), .O(gate800inter8));
  nand2 gate1296(.a(gate800inter8), .b(gate800inter7), .O(gate800inter9));
  nand2 gate1297(.a(s_59), .b(gate800inter3), .O(gate800inter10));
  nor2  gate1298(.a(gate800inter10), .b(gate800inter9), .O(gate800inter11));
  nor2  gate1299(.a(gate800inter11), .b(gate800inter6), .O(gate800inter12));
  nand2 gate1300(.a(gate800inter12), .b(gate800inter1), .O(N2759));

  xor2  gate2799(.a(N2731), .b(N364), .O(gate801inter0));
  nand2 gate2800(.a(gate801inter0), .b(s_274), .O(gate801inter1));
  and2  gate2801(.a(N2731), .b(N364), .O(gate801inter2));
  inv1  gate2802(.a(s_274), .O(gate801inter3));
  inv1  gate2803(.a(s_275), .O(gate801inter4));
  nand2 gate2804(.a(gate801inter4), .b(gate801inter3), .O(gate801inter5));
  nor2  gate2805(.a(gate801inter5), .b(gate801inter2), .O(gate801inter6));
  inv1  gate2806(.a(N364), .O(gate801inter7));
  inv1  gate2807(.a(N2731), .O(gate801inter8));
  nand2 gate2808(.a(gate801inter8), .b(gate801inter7), .O(gate801inter9));
  nand2 gate2809(.a(s_275), .b(gate801inter3), .O(gate801inter10));
  nor2  gate2810(.a(gate801inter10), .b(gate801inter9), .O(gate801inter11));
  nor2  gate2811(.a(gate801inter11), .b(gate801inter6), .O(gate801inter12));
  nand2 gate2812(.a(gate801inter12), .b(gate801inter1), .O(N2760));
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );

  xor2  gate1777(.a(N2736), .b(N373), .O(gate804inter0));
  nand2 gate1778(.a(gate804inter0), .b(s_128), .O(gate804inter1));
  and2  gate1779(.a(N2736), .b(N373), .O(gate804inter2));
  inv1  gate1780(.a(s_128), .O(gate804inter3));
  inv1  gate1781(.a(s_129), .O(gate804inter4));
  nand2 gate1782(.a(gate804inter4), .b(gate804inter3), .O(gate804inter5));
  nor2  gate1783(.a(gate804inter5), .b(gate804inter2), .O(gate804inter6));
  inv1  gate1784(.a(N373), .O(gate804inter7));
  inv1  gate1785(.a(N2736), .O(gate804inter8));
  nand2 gate1786(.a(gate804inter8), .b(gate804inter7), .O(gate804inter9));
  nand2 gate1787(.a(s_129), .b(gate804inter3), .O(gate804inter10));
  nor2  gate1788(.a(gate804inter10), .b(gate804inter9), .O(gate804inter11));
  nor2  gate1789(.a(gate804inter11), .b(gate804inter6), .O(gate804inter12));
  nand2 gate1790(.a(gate804inter12), .b(gate804inter1), .O(N2763));
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );

  xor2  gate1637(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate1638(.a(gate806inter0), .b(s_108), .O(gate806inter1));
  and2  gate1639(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate1640(.a(s_108), .O(gate806inter3));
  inv1  gate1641(.a(s_109), .O(gate806inter4));
  nand2 gate1642(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate1643(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate1644(.a(N379), .O(gate806inter7));
  inv1  gate1645(.a(N2740), .O(gate806inter8));
  nand2 gate1646(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate1647(.a(s_109), .b(gate806inter3), .O(gate806inter10));
  nor2  gate1648(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate1649(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate1650(.a(gate806inter12), .b(gate806inter1), .O(N2765));

  xor2  gate2631(.a(N2742), .b(N382), .O(gate807inter0));
  nand2 gate2632(.a(gate807inter0), .b(s_250), .O(gate807inter1));
  and2  gate2633(.a(N2742), .b(N382), .O(gate807inter2));
  inv1  gate2634(.a(s_250), .O(gate807inter3));
  inv1  gate2635(.a(s_251), .O(gate807inter4));
  nand2 gate2636(.a(gate807inter4), .b(gate807inter3), .O(gate807inter5));
  nor2  gate2637(.a(gate807inter5), .b(gate807inter2), .O(gate807inter6));
  inv1  gate2638(.a(N382), .O(gate807inter7));
  inv1  gate2639(.a(N2742), .O(gate807inter8));
  nand2 gate2640(.a(gate807inter8), .b(gate807inter7), .O(gate807inter9));
  nand2 gate2641(.a(s_251), .b(gate807inter3), .O(gate807inter10));
  nor2  gate2642(.a(gate807inter10), .b(gate807inter9), .O(gate807inter11));
  nor2  gate2643(.a(gate807inter11), .b(gate807inter6), .O(gate807inter12));
  nand2 gate2644(.a(gate807inter12), .b(gate807inter1), .O(N2766));

  xor2  gate1945(.a(N2743), .b(N2688), .O(gate808inter0));
  nand2 gate1946(.a(gate808inter0), .b(s_152), .O(gate808inter1));
  and2  gate1947(.a(N2743), .b(N2688), .O(gate808inter2));
  inv1  gate1948(.a(s_152), .O(gate808inter3));
  inv1  gate1949(.a(s_153), .O(gate808inter4));
  nand2 gate1950(.a(gate808inter4), .b(gate808inter3), .O(gate808inter5));
  nor2  gate1951(.a(gate808inter5), .b(gate808inter2), .O(gate808inter6));
  inv1  gate1952(.a(N2688), .O(gate808inter7));
  inv1  gate1953(.a(N2743), .O(gate808inter8));
  nand2 gate1954(.a(gate808inter8), .b(gate808inter7), .O(gate808inter9));
  nand2 gate1955(.a(s_153), .b(gate808inter3), .O(gate808inter10));
  nor2  gate1956(.a(gate808inter10), .b(gate808inter9), .O(gate808inter11));
  nor2  gate1957(.a(gate808inter11), .b(gate808inter6), .O(gate808inter12));
  nand2 gate1958(.a(gate808inter12), .b(gate808inter1), .O(N2767));
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );

  xor2  gate1399(.a(N2759), .b(N2728), .O(gate814inter0));
  nand2 gate1400(.a(gate814inter0), .b(s_74), .O(gate814inter1));
  and2  gate1401(.a(N2759), .b(N2728), .O(gate814inter2));
  inv1  gate1402(.a(s_74), .O(gate814inter3));
  inv1  gate1403(.a(s_75), .O(gate814inter4));
  nand2 gate1404(.a(gate814inter4), .b(gate814inter3), .O(gate814inter5));
  nor2  gate1405(.a(gate814inter5), .b(gate814inter2), .O(gate814inter6));
  inv1  gate1406(.a(N2728), .O(gate814inter7));
  inv1  gate1407(.a(N2759), .O(gate814inter8));
  nand2 gate1408(.a(gate814inter8), .b(gate814inter7), .O(gate814inter9));
  nand2 gate1409(.a(s_75), .b(gate814inter3), .O(gate814inter10));
  nor2  gate1410(.a(gate814inter10), .b(gate814inter9), .O(gate814inter11));
  nor2  gate1411(.a(gate814inter11), .b(gate814inter6), .O(gate814inter12));
  nand2 gate1412(.a(gate814inter12), .b(gate814inter1), .O(N2781));
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );

  xor2  gate2365(.a(N2761), .b(N2732), .O(gate816inter0));
  nand2 gate2366(.a(gate816inter0), .b(s_212), .O(gate816inter1));
  and2  gate2367(.a(N2761), .b(N2732), .O(gate816inter2));
  inv1  gate2368(.a(s_212), .O(gate816inter3));
  inv1  gate2369(.a(s_213), .O(gate816inter4));
  nand2 gate2370(.a(gate816inter4), .b(gate816inter3), .O(gate816inter5));
  nor2  gate2371(.a(gate816inter5), .b(gate816inter2), .O(gate816inter6));
  inv1  gate2372(.a(N2732), .O(gate816inter7));
  inv1  gate2373(.a(N2761), .O(gate816inter8));
  nand2 gate2374(.a(gate816inter8), .b(gate816inter7), .O(gate816inter9));
  nand2 gate2375(.a(s_213), .b(gate816inter3), .O(gate816inter10));
  nor2  gate2376(.a(gate816inter10), .b(gate816inter9), .O(gate816inter11));
  nor2  gate2377(.a(gate816inter11), .b(gate816inter6), .O(gate816inter12));
  nand2 gate2378(.a(gate816inter12), .b(gate816inter1), .O(N2783));

  xor2  gate1735(.a(N2763), .b(N2735), .O(gate817inter0));
  nand2 gate1736(.a(gate817inter0), .b(s_122), .O(gate817inter1));
  and2  gate1737(.a(N2763), .b(N2735), .O(gate817inter2));
  inv1  gate1738(.a(s_122), .O(gate817inter3));
  inv1  gate1739(.a(s_123), .O(gate817inter4));
  nand2 gate1740(.a(gate817inter4), .b(gate817inter3), .O(gate817inter5));
  nor2  gate1741(.a(gate817inter5), .b(gate817inter2), .O(gate817inter6));
  inv1  gate1742(.a(N2735), .O(gate817inter7));
  inv1  gate1743(.a(N2763), .O(gate817inter8));
  nand2 gate1744(.a(gate817inter8), .b(gate817inter7), .O(gate817inter9));
  nand2 gate1745(.a(s_123), .b(gate817inter3), .O(gate817inter10));
  nor2  gate1746(.a(gate817inter10), .b(gate817inter9), .O(gate817inter11));
  nor2  gate1747(.a(gate817inter11), .b(gate817inter6), .O(gate817inter12));
  nand2 gate1748(.a(gate817inter12), .b(gate817inter1), .O(N2784));

  xor2  gate1343(.a(N2764), .b(N2737), .O(gate818inter0));
  nand2 gate1344(.a(gate818inter0), .b(s_66), .O(gate818inter1));
  and2  gate1345(.a(N2764), .b(N2737), .O(gate818inter2));
  inv1  gate1346(.a(s_66), .O(gate818inter3));
  inv1  gate1347(.a(s_67), .O(gate818inter4));
  nand2 gate1348(.a(gate818inter4), .b(gate818inter3), .O(gate818inter5));
  nor2  gate1349(.a(gate818inter5), .b(gate818inter2), .O(gate818inter6));
  inv1  gate1350(.a(N2737), .O(gate818inter7));
  inv1  gate1351(.a(N2764), .O(gate818inter8));
  nand2 gate1352(.a(gate818inter8), .b(gate818inter7), .O(gate818inter9));
  nand2 gate1353(.a(s_67), .b(gate818inter3), .O(gate818inter10));
  nor2  gate1354(.a(gate818inter10), .b(gate818inter9), .O(gate818inter11));
  nor2  gate1355(.a(gate818inter11), .b(gate818inter6), .O(gate818inter12));
  nand2 gate1356(.a(gate818inter12), .b(gate818inter1), .O(N2785));

  xor2  gate1357(.a(N2765), .b(N2739), .O(gate819inter0));
  nand2 gate1358(.a(gate819inter0), .b(s_68), .O(gate819inter1));
  and2  gate1359(.a(N2765), .b(N2739), .O(gate819inter2));
  inv1  gate1360(.a(s_68), .O(gate819inter3));
  inv1  gate1361(.a(s_69), .O(gate819inter4));
  nand2 gate1362(.a(gate819inter4), .b(gate819inter3), .O(gate819inter5));
  nor2  gate1363(.a(gate819inter5), .b(gate819inter2), .O(gate819inter6));
  inv1  gate1364(.a(N2739), .O(gate819inter7));
  inv1  gate1365(.a(N2765), .O(gate819inter8));
  nand2 gate1366(.a(gate819inter8), .b(gate819inter7), .O(gate819inter9));
  nand2 gate1367(.a(s_69), .b(gate819inter3), .O(gate819inter10));
  nor2  gate1368(.a(gate819inter10), .b(gate819inter9), .O(gate819inter11));
  nor2  gate1369(.a(gate819inter11), .b(gate819inter6), .O(gate819inter12));
  nand2 gate1370(.a(gate819inter12), .b(gate819inter1), .O(N2786));
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );

  xor2  gate1049(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate1050(.a(gate839inter0), .b(s_24), .O(gate839inter1));
  and2  gate1051(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate1052(.a(s_24), .O(gate839inter3));
  inv1  gate1053(.a(s_25), .O(gate839inter4));
  nand2 gate1054(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate1055(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate1056(.a(N2812), .O(gate839inter7));
  inv1  gate1057(.a(N2076), .O(gate839inter8));
  nand2 gate1058(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate1059(.a(s_25), .b(gate839inter3), .O(gate839inter10));
  nor2  gate1060(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate1061(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate1062(.a(gate839inter12), .b(gate839inter1), .O(N2850));

  xor2  gate909(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate910(.a(gate840inter0), .b(s_4), .O(gate840inter1));
  and2  gate911(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate912(.a(s_4), .O(gate840inter3));
  inv1  gate913(.a(s_5), .O(gate840inter4));
  nand2 gate914(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate915(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate916(.a(N2815), .O(gate840inter7));
  inv1  gate917(.a(N2077), .O(gate840inter8));
  nand2 gate918(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate919(.a(s_5), .b(gate840inter3), .O(gate840inter10));
  nor2  gate920(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate921(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate922(.a(gate840inter12), .b(gate840inter1), .O(N2851));
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );

  xor2  gate1315(.a(N1938), .b(N2824), .O(gate843inter0));
  nand2 gate1316(.a(gate843inter0), .b(s_62), .O(gate843inter1));
  and2  gate1317(.a(N1938), .b(N2824), .O(gate843inter2));
  inv1  gate1318(.a(s_62), .O(gate843inter3));
  inv1  gate1319(.a(s_63), .O(gate843inter4));
  nand2 gate1320(.a(gate843inter4), .b(gate843inter3), .O(gate843inter5));
  nor2  gate1321(.a(gate843inter5), .b(gate843inter2), .O(gate843inter6));
  inv1  gate1322(.a(N2824), .O(gate843inter7));
  inv1  gate1323(.a(N1938), .O(gate843inter8));
  nand2 gate1324(.a(gate843inter8), .b(gate843inter7), .O(gate843inter9));
  nand2 gate1325(.a(s_63), .b(gate843inter3), .O(gate843inter10));
  nor2  gate1326(.a(gate843inter10), .b(gate843inter9), .O(gate843inter11));
  nor2  gate1327(.a(gate843inter11), .b(gate843inter6), .O(gate843inter12));
  nand2 gate1328(.a(gate843inter12), .b(gate843inter1), .O(N2854));
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );

  xor2  gate923(.a(N2857), .b(N2052), .O(gate851inter0));
  nand2 gate924(.a(gate851inter0), .b(s_6), .O(gate851inter1));
  and2  gate925(.a(N2857), .b(N2052), .O(gate851inter2));
  inv1  gate926(.a(s_6), .O(gate851inter3));
  inv1  gate927(.a(s_7), .O(gate851inter4));
  nand2 gate928(.a(gate851inter4), .b(gate851inter3), .O(gate851inter5));
  nor2  gate929(.a(gate851inter5), .b(gate851inter2), .O(gate851inter6));
  inv1  gate930(.a(N2052), .O(gate851inter7));
  inv1  gate931(.a(N2857), .O(gate851inter8));
  nand2 gate932(.a(gate851inter8), .b(gate851inter7), .O(gate851inter9));
  nand2 gate933(.a(s_7), .b(gate851inter3), .O(gate851inter10));
  nor2  gate934(.a(gate851inter10), .b(gate851inter9), .O(gate851inter11));
  nor2  gate935(.a(gate851inter11), .b(gate851inter6), .O(gate851inter12));
  nand2 gate936(.a(gate851inter12), .b(gate851inter1), .O(N2866));
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate2477(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate2478(.a(gate860inter0), .b(s_228), .O(gate860inter1));
  and2  gate2479(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate2480(.a(s_228), .O(gate860inter3));
  inv1  gate2481(.a(s_229), .O(gate860inter4));
  nand2 gate2482(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate2483(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate2484(.a(N1933), .O(gate860inter7));
  inv1  gate2485(.a(N2862), .O(gate860inter8));
  nand2 gate2486(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate2487(.a(s_229), .b(gate860inter3), .O(gate860inter10));
  nor2  gate2488(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate2489(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate2490(.a(gate860inter12), .b(gate860inter1), .O(N2875));
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );

  xor2  gate2267(.a(N2853), .b(N2869), .O(gate864inter0));
  nand2 gate2268(.a(gate864inter0), .b(s_198), .O(gate864inter1));
  and2  gate2269(.a(N2853), .b(N2869), .O(gate864inter2));
  inv1  gate2270(.a(s_198), .O(gate864inter3));
  inv1  gate2271(.a(s_199), .O(gate864inter4));
  nand2 gate2272(.a(gate864inter4), .b(gate864inter3), .O(gate864inter5));
  nor2  gate2273(.a(gate864inter5), .b(gate864inter2), .O(gate864inter6));
  inv1  gate2274(.a(N2869), .O(gate864inter7));
  inv1  gate2275(.a(N2853), .O(gate864inter8));
  nand2 gate2276(.a(gate864inter8), .b(gate864inter7), .O(gate864inter9));
  nand2 gate2277(.a(s_199), .b(gate864inter3), .O(gate864inter10));
  nor2  gate2278(.a(gate864inter10), .b(gate864inter9), .O(gate864inter11));
  nor2  gate2279(.a(gate864inter11), .b(gate864inter6), .O(gate864inter12));
  nand2 gate2280(.a(gate864inter12), .b(gate864inter1), .O(N2879));
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );

  xor2  gate2855(.a(N2874), .b(N685), .O(gate867inter0));
  nand2 gate2856(.a(gate867inter0), .b(s_282), .O(gate867inter1));
  and2  gate2857(.a(N2874), .b(N685), .O(gate867inter2));
  inv1  gate2858(.a(s_282), .O(gate867inter3));
  inv1  gate2859(.a(s_283), .O(gate867inter4));
  nand2 gate2860(.a(gate867inter4), .b(gate867inter3), .O(gate867inter5));
  nor2  gate2861(.a(gate867inter5), .b(gate867inter2), .O(gate867inter6));
  inv1  gate2862(.a(N685), .O(gate867inter7));
  inv1  gate2863(.a(N2874), .O(gate867inter8));
  nand2 gate2864(.a(gate867inter8), .b(gate867inter7), .O(gate867inter9));
  nand2 gate2865(.a(s_283), .b(gate867inter3), .O(gate867inter10));
  nor2  gate2866(.a(gate867inter10), .b(gate867inter9), .O(gate867inter11));
  nor2  gate2867(.a(gate867inter11), .b(gate867inter6), .O(gate867inter12));
  nand2 gate2868(.a(gate867inter12), .b(gate867inter1), .O(N2882));

  xor2  gate1385(.a(N2863), .b(N2875), .O(gate868inter0));
  nand2 gate1386(.a(gate868inter0), .b(s_72), .O(gate868inter1));
  and2  gate1387(.a(N2863), .b(N2875), .O(gate868inter2));
  inv1  gate1388(.a(s_72), .O(gate868inter3));
  inv1  gate1389(.a(s_73), .O(gate868inter4));
  nand2 gate1390(.a(gate868inter4), .b(gate868inter3), .O(gate868inter5));
  nor2  gate1391(.a(gate868inter5), .b(gate868inter2), .O(gate868inter6));
  inv1  gate1392(.a(N2875), .O(gate868inter7));
  inv1  gate1393(.a(N2863), .O(gate868inter8));
  nand2 gate1394(.a(gate868inter8), .b(gate868inter7), .O(gate868inter9));
  nand2 gate1395(.a(s_73), .b(gate868inter3), .O(gate868inter10));
  nor2  gate1396(.a(gate868inter10), .b(gate868inter9), .O(gate868inter11));
  nor2  gate1397(.a(gate868inter11), .b(gate868inter6), .O(gate868inter12));
  nand2 gate1398(.a(gate868inter12), .b(gate868inter1), .O(N2883));
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate2743(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate2744(.a(gate874inter0), .b(s_266), .O(gate874inter1));
  and2  gate2745(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate2746(.a(s_266), .O(gate874inter3));
  inv1  gate2747(.a(s_267), .O(gate874inter4));
  nand2 gate2748(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate2749(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate2750(.a(N2871), .O(gate874inter7));
  inv1  gate2751(.a(N2881), .O(gate874inter8));
  nand2 gate2752(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate2753(.a(s_267), .b(gate874inter3), .O(gate874inter10));
  nor2  gate2754(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate2755(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate2756(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );

  xor2  gate2435(.a(N2897), .b(N2895), .O(gate879inter0));
  nand2 gate2436(.a(gate879inter0), .b(s_222), .O(gate879inter1));
  and2  gate2437(.a(N2897), .b(N2895), .O(gate879inter2));
  inv1  gate2438(.a(s_222), .O(gate879inter3));
  inv1  gate2439(.a(s_223), .O(gate879inter4));
  nand2 gate2440(.a(gate879inter4), .b(gate879inter3), .O(gate879inter5));
  nor2  gate2441(.a(gate879inter5), .b(gate879inter2), .O(gate879inter6));
  inv1  gate2442(.a(N2895), .O(gate879inter7));
  inv1  gate2443(.a(N2897), .O(gate879inter8));
  nand2 gate2444(.a(gate879inter8), .b(gate879inter7), .O(gate879inter9));
  nand2 gate2445(.a(s_223), .b(gate879inter3), .O(gate879inter10));
  nor2  gate2446(.a(gate879inter10), .b(gate879inter9), .O(gate879inter11));
  nor2  gate2447(.a(gate879inter11), .b(gate879inter6), .O(gate879inter12));
  nand2 gate2448(.a(gate879inter12), .b(gate879inter1), .O(N2898));
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule