module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1471(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1472(.a(gate9inter0), .b(s_132), .O(gate9inter1));
  and2  gate1473(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1474(.a(s_132), .O(gate9inter3));
  inv1  gate1475(.a(s_133), .O(gate9inter4));
  nand2 gate1476(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1477(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1478(.a(G1), .O(gate9inter7));
  inv1  gate1479(.a(G2), .O(gate9inter8));
  nand2 gate1480(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1481(.a(s_133), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1482(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1483(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1484(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1793(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1794(.a(gate12inter0), .b(s_178), .O(gate12inter1));
  and2  gate1795(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1796(.a(s_178), .O(gate12inter3));
  inv1  gate1797(.a(s_179), .O(gate12inter4));
  nand2 gate1798(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1799(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1800(.a(G7), .O(gate12inter7));
  inv1  gate1801(.a(G8), .O(gate12inter8));
  nand2 gate1802(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1803(.a(s_179), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1804(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1805(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1806(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2619(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2620(.a(gate13inter0), .b(s_296), .O(gate13inter1));
  and2  gate2621(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2622(.a(s_296), .O(gate13inter3));
  inv1  gate2623(.a(s_297), .O(gate13inter4));
  nand2 gate2624(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2625(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2626(.a(G9), .O(gate13inter7));
  inv1  gate2627(.a(G10), .O(gate13inter8));
  nand2 gate2628(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2629(.a(s_297), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2630(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2631(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2632(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2675(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2676(.a(gate15inter0), .b(s_304), .O(gate15inter1));
  and2  gate2677(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2678(.a(s_304), .O(gate15inter3));
  inv1  gate2679(.a(s_305), .O(gate15inter4));
  nand2 gate2680(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2681(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2682(.a(G13), .O(gate15inter7));
  inv1  gate2683(.a(G14), .O(gate15inter8));
  nand2 gate2684(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2685(.a(s_305), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2686(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2687(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2688(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2143(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2144(.a(gate17inter0), .b(s_228), .O(gate17inter1));
  and2  gate2145(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2146(.a(s_228), .O(gate17inter3));
  inv1  gate2147(.a(s_229), .O(gate17inter4));
  nand2 gate2148(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2149(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2150(.a(G17), .O(gate17inter7));
  inv1  gate2151(.a(G18), .O(gate17inter8));
  nand2 gate2152(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2153(.a(s_229), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2154(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2155(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2156(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2563(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2564(.a(gate19inter0), .b(s_288), .O(gate19inter1));
  and2  gate2565(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2566(.a(s_288), .O(gate19inter3));
  inv1  gate2567(.a(s_289), .O(gate19inter4));
  nand2 gate2568(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2569(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2570(.a(G21), .O(gate19inter7));
  inv1  gate2571(.a(G22), .O(gate19inter8));
  nand2 gate2572(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2573(.a(s_289), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2574(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2575(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2576(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate673(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate674(.a(gate23inter0), .b(s_18), .O(gate23inter1));
  and2  gate675(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate676(.a(s_18), .O(gate23inter3));
  inv1  gate677(.a(s_19), .O(gate23inter4));
  nand2 gate678(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate679(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate680(.a(G29), .O(gate23inter7));
  inv1  gate681(.a(G30), .O(gate23inter8));
  nand2 gate682(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate683(.a(s_19), .b(gate23inter3), .O(gate23inter10));
  nor2  gate684(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate685(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate686(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2857(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2858(.a(gate25inter0), .b(s_330), .O(gate25inter1));
  and2  gate2859(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2860(.a(s_330), .O(gate25inter3));
  inv1  gate2861(.a(s_331), .O(gate25inter4));
  nand2 gate2862(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2863(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2864(.a(G1), .O(gate25inter7));
  inv1  gate2865(.a(G5), .O(gate25inter8));
  nand2 gate2866(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2867(.a(s_331), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2868(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2869(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2870(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate701(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate702(.a(gate33inter0), .b(s_22), .O(gate33inter1));
  and2  gate703(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate704(.a(s_22), .O(gate33inter3));
  inv1  gate705(.a(s_23), .O(gate33inter4));
  nand2 gate706(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate707(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate708(.a(G17), .O(gate33inter7));
  inv1  gate709(.a(G21), .O(gate33inter8));
  nand2 gate710(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate711(.a(s_23), .b(gate33inter3), .O(gate33inter10));
  nor2  gate712(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate713(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate714(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2101(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2102(.a(gate35inter0), .b(s_222), .O(gate35inter1));
  and2  gate2103(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2104(.a(s_222), .O(gate35inter3));
  inv1  gate2105(.a(s_223), .O(gate35inter4));
  nand2 gate2106(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2107(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2108(.a(G18), .O(gate35inter7));
  inv1  gate2109(.a(G22), .O(gate35inter8));
  nand2 gate2110(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2111(.a(s_223), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2112(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2113(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2114(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2339(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2340(.a(gate36inter0), .b(s_256), .O(gate36inter1));
  and2  gate2341(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2342(.a(s_256), .O(gate36inter3));
  inv1  gate2343(.a(s_257), .O(gate36inter4));
  nand2 gate2344(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2345(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2346(.a(G26), .O(gate36inter7));
  inv1  gate2347(.a(G30), .O(gate36inter8));
  nand2 gate2348(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2349(.a(s_257), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2350(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2351(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2352(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate757(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate758(.a(gate38inter0), .b(s_30), .O(gate38inter1));
  and2  gate759(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate760(.a(s_30), .O(gate38inter3));
  inv1  gate761(.a(s_31), .O(gate38inter4));
  nand2 gate762(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate763(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate764(.a(G27), .O(gate38inter7));
  inv1  gate765(.a(G31), .O(gate38inter8));
  nand2 gate766(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate767(.a(s_31), .b(gate38inter3), .O(gate38inter10));
  nor2  gate768(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate769(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate770(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1681(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1682(.a(gate41inter0), .b(s_162), .O(gate41inter1));
  and2  gate1683(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1684(.a(s_162), .O(gate41inter3));
  inv1  gate1685(.a(s_163), .O(gate41inter4));
  nand2 gate1686(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1687(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1688(.a(G1), .O(gate41inter7));
  inv1  gate1689(.a(G266), .O(gate41inter8));
  nand2 gate1690(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1691(.a(s_163), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1692(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1693(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1694(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2059(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2060(.a(gate42inter0), .b(s_216), .O(gate42inter1));
  and2  gate2061(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2062(.a(s_216), .O(gate42inter3));
  inv1  gate2063(.a(s_217), .O(gate42inter4));
  nand2 gate2064(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2065(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2066(.a(G2), .O(gate42inter7));
  inv1  gate2067(.a(G266), .O(gate42inter8));
  nand2 gate2068(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2069(.a(s_217), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2070(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2071(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2072(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2605(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2606(.a(gate47inter0), .b(s_294), .O(gate47inter1));
  and2  gate2607(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2608(.a(s_294), .O(gate47inter3));
  inv1  gate2609(.a(s_295), .O(gate47inter4));
  nand2 gate2610(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2611(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2612(.a(G7), .O(gate47inter7));
  inv1  gate2613(.a(G275), .O(gate47inter8));
  nand2 gate2614(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2615(.a(s_295), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2616(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2617(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2618(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate827(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate828(.a(gate49inter0), .b(s_40), .O(gate49inter1));
  and2  gate829(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate830(.a(s_40), .O(gate49inter3));
  inv1  gate831(.a(s_41), .O(gate49inter4));
  nand2 gate832(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate833(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate834(.a(G9), .O(gate49inter7));
  inv1  gate835(.a(G278), .O(gate49inter8));
  nand2 gate836(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate837(.a(s_41), .b(gate49inter3), .O(gate49inter10));
  nor2  gate838(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate839(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate840(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2423(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2424(.a(gate52inter0), .b(s_268), .O(gate52inter1));
  and2  gate2425(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2426(.a(s_268), .O(gate52inter3));
  inv1  gate2427(.a(s_269), .O(gate52inter4));
  nand2 gate2428(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2429(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2430(.a(G12), .O(gate52inter7));
  inv1  gate2431(.a(G281), .O(gate52inter8));
  nand2 gate2432(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2433(.a(s_269), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2434(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2435(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2436(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1107(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1108(.a(gate53inter0), .b(s_80), .O(gate53inter1));
  and2  gate1109(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1110(.a(s_80), .O(gate53inter3));
  inv1  gate1111(.a(s_81), .O(gate53inter4));
  nand2 gate1112(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1113(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1114(.a(G13), .O(gate53inter7));
  inv1  gate1115(.a(G284), .O(gate53inter8));
  nand2 gate1116(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1117(.a(s_81), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1118(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1119(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1120(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1919(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1920(.a(gate55inter0), .b(s_196), .O(gate55inter1));
  and2  gate1921(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1922(.a(s_196), .O(gate55inter3));
  inv1  gate1923(.a(s_197), .O(gate55inter4));
  nand2 gate1924(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1925(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1926(.a(G15), .O(gate55inter7));
  inv1  gate1927(.a(G287), .O(gate55inter8));
  nand2 gate1928(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1929(.a(s_197), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1930(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1931(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1932(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2717(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2718(.a(gate56inter0), .b(s_310), .O(gate56inter1));
  and2  gate2719(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2720(.a(s_310), .O(gate56inter3));
  inv1  gate2721(.a(s_311), .O(gate56inter4));
  nand2 gate2722(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2723(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2724(.a(G16), .O(gate56inter7));
  inv1  gate2725(.a(G287), .O(gate56inter8));
  nand2 gate2726(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2727(.a(s_311), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2728(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2729(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2730(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2451(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2452(.a(gate58inter0), .b(s_272), .O(gate58inter1));
  and2  gate2453(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2454(.a(s_272), .O(gate58inter3));
  inv1  gate2455(.a(s_273), .O(gate58inter4));
  nand2 gate2456(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2457(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2458(.a(G18), .O(gate58inter7));
  inv1  gate2459(.a(G290), .O(gate58inter8));
  nand2 gate2460(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2461(.a(s_273), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2462(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2463(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2464(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1947(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1948(.a(gate59inter0), .b(s_200), .O(gate59inter1));
  and2  gate1949(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1950(.a(s_200), .O(gate59inter3));
  inv1  gate1951(.a(s_201), .O(gate59inter4));
  nand2 gate1952(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1953(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1954(.a(G19), .O(gate59inter7));
  inv1  gate1955(.a(G293), .O(gate59inter8));
  nand2 gate1956(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1957(.a(s_201), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1958(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1959(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1960(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate911(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate912(.a(gate63inter0), .b(s_52), .O(gate63inter1));
  and2  gate913(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate914(.a(s_52), .O(gate63inter3));
  inv1  gate915(.a(s_53), .O(gate63inter4));
  nand2 gate916(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate917(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate918(.a(G23), .O(gate63inter7));
  inv1  gate919(.a(G299), .O(gate63inter8));
  nand2 gate920(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate921(.a(s_53), .b(gate63inter3), .O(gate63inter10));
  nor2  gate922(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate923(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate924(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1331(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1332(.a(gate64inter0), .b(s_112), .O(gate64inter1));
  and2  gate1333(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1334(.a(s_112), .O(gate64inter3));
  inv1  gate1335(.a(s_113), .O(gate64inter4));
  nand2 gate1336(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1337(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1338(.a(G24), .O(gate64inter7));
  inv1  gate1339(.a(G299), .O(gate64inter8));
  nand2 gate1340(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1341(.a(s_113), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1342(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1343(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1344(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate2213(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2214(.a(gate65inter0), .b(s_238), .O(gate65inter1));
  and2  gate2215(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2216(.a(s_238), .O(gate65inter3));
  inv1  gate2217(.a(s_239), .O(gate65inter4));
  nand2 gate2218(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2219(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2220(.a(G25), .O(gate65inter7));
  inv1  gate2221(.a(G302), .O(gate65inter8));
  nand2 gate2222(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2223(.a(s_239), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2224(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2225(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2226(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1275(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1276(.a(gate68inter0), .b(s_104), .O(gate68inter1));
  and2  gate1277(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1278(.a(s_104), .O(gate68inter3));
  inv1  gate1279(.a(s_105), .O(gate68inter4));
  nand2 gate1280(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1281(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1282(.a(G28), .O(gate68inter7));
  inv1  gate1283(.a(G305), .O(gate68inter8));
  nand2 gate1284(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1285(.a(s_105), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1286(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1287(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1288(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1849(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1850(.a(gate70inter0), .b(s_186), .O(gate70inter1));
  and2  gate1851(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1852(.a(s_186), .O(gate70inter3));
  inv1  gate1853(.a(s_187), .O(gate70inter4));
  nand2 gate1854(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1855(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1856(.a(G30), .O(gate70inter7));
  inv1  gate1857(.a(G308), .O(gate70inter8));
  nand2 gate1858(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1859(.a(s_187), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1860(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1861(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1862(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1135(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1136(.a(gate73inter0), .b(s_84), .O(gate73inter1));
  and2  gate1137(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1138(.a(s_84), .O(gate73inter3));
  inv1  gate1139(.a(s_85), .O(gate73inter4));
  nand2 gate1140(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1141(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1142(.a(G1), .O(gate73inter7));
  inv1  gate1143(.a(G314), .O(gate73inter8));
  nand2 gate1144(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1145(.a(s_85), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1146(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1147(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1148(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2661(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2662(.a(gate76inter0), .b(s_302), .O(gate76inter1));
  and2  gate2663(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2664(.a(s_302), .O(gate76inter3));
  inv1  gate2665(.a(s_303), .O(gate76inter4));
  nand2 gate2666(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2667(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2668(.a(G13), .O(gate76inter7));
  inv1  gate2669(.a(G317), .O(gate76inter8));
  nand2 gate2670(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2671(.a(s_303), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2672(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2673(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2674(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1037(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1038(.a(gate78inter0), .b(s_70), .O(gate78inter1));
  and2  gate1039(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1040(.a(s_70), .O(gate78inter3));
  inv1  gate1041(.a(s_71), .O(gate78inter4));
  nand2 gate1042(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1043(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1044(.a(G6), .O(gate78inter7));
  inv1  gate1045(.a(G320), .O(gate78inter8));
  nand2 gate1046(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1047(.a(s_71), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1048(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1049(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1050(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1835(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1836(.a(gate84inter0), .b(s_184), .O(gate84inter1));
  and2  gate1837(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1838(.a(s_184), .O(gate84inter3));
  inv1  gate1839(.a(s_185), .O(gate84inter4));
  nand2 gate1840(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1841(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1842(.a(G15), .O(gate84inter7));
  inv1  gate1843(.a(G329), .O(gate84inter8));
  nand2 gate1844(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1845(.a(s_185), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1846(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1847(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1848(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1821(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1822(.a(gate87inter0), .b(s_182), .O(gate87inter1));
  and2  gate1823(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1824(.a(s_182), .O(gate87inter3));
  inv1  gate1825(.a(s_183), .O(gate87inter4));
  nand2 gate1826(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1827(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1828(.a(G12), .O(gate87inter7));
  inv1  gate1829(.a(G335), .O(gate87inter8));
  nand2 gate1830(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1831(.a(s_183), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1832(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1833(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1834(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate841(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate842(.a(gate88inter0), .b(s_42), .O(gate88inter1));
  and2  gate843(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate844(.a(s_42), .O(gate88inter3));
  inv1  gate845(.a(s_43), .O(gate88inter4));
  nand2 gate846(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate847(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate848(.a(G16), .O(gate88inter7));
  inv1  gate849(.a(G335), .O(gate88inter8));
  nand2 gate850(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate851(.a(s_43), .b(gate88inter3), .O(gate88inter10));
  nor2  gate852(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate853(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate854(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2227(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2228(.a(gate89inter0), .b(s_240), .O(gate89inter1));
  and2  gate2229(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2230(.a(s_240), .O(gate89inter3));
  inv1  gate2231(.a(s_241), .O(gate89inter4));
  nand2 gate2232(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2233(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2234(.a(G17), .O(gate89inter7));
  inv1  gate2235(.a(G338), .O(gate89inter8));
  nand2 gate2236(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2237(.a(s_241), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2238(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2239(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2240(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2731(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2732(.a(gate91inter0), .b(s_312), .O(gate91inter1));
  and2  gate2733(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2734(.a(s_312), .O(gate91inter3));
  inv1  gate2735(.a(s_313), .O(gate91inter4));
  nand2 gate2736(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2737(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2738(.a(G25), .O(gate91inter7));
  inv1  gate2739(.a(G341), .O(gate91inter8));
  nand2 gate2740(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2741(.a(s_313), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2742(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2743(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2744(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1905(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1906(.a(gate95inter0), .b(s_194), .O(gate95inter1));
  and2  gate1907(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1908(.a(s_194), .O(gate95inter3));
  inv1  gate1909(.a(s_195), .O(gate95inter4));
  nand2 gate1910(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1911(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1912(.a(G26), .O(gate95inter7));
  inv1  gate1913(.a(G347), .O(gate95inter8));
  nand2 gate1914(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1915(.a(s_195), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1916(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1917(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1918(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2507(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2508(.a(gate97inter0), .b(s_280), .O(gate97inter1));
  and2  gate2509(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2510(.a(s_280), .O(gate97inter3));
  inv1  gate2511(.a(s_281), .O(gate97inter4));
  nand2 gate2512(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2513(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2514(.a(G19), .O(gate97inter7));
  inv1  gate2515(.a(G350), .O(gate97inter8));
  nand2 gate2516(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2517(.a(s_281), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2518(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2519(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2520(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1611(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1612(.a(gate98inter0), .b(s_152), .O(gate98inter1));
  and2  gate1613(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1614(.a(s_152), .O(gate98inter3));
  inv1  gate1615(.a(s_153), .O(gate98inter4));
  nand2 gate1616(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1617(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1618(.a(G23), .O(gate98inter7));
  inv1  gate1619(.a(G350), .O(gate98inter8));
  nand2 gate1620(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1621(.a(s_153), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1622(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1623(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1624(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2815(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2816(.a(gate99inter0), .b(s_324), .O(gate99inter1));
  and2  gate2817(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2818(.a(s_324), .O(gate99inter3));
  inv1  gate2819(.a(s_325), .O(gate99inter4));
  nand2 gate2820(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2821(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2822(.a(G27), .O(gate99inter7));
  inv1  gate2823(.a(G353), .O(gate99inter8));
  nand2 gate2824(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2825(.a(s_325), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2826(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2827(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2828(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate2185(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2186(.a(gate100inter0), .b(s_234), .O(gate100inter1));
  and2  gate2187(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2188(.a(s_234), .O(gate100inter3));
  inv1  gate2189(.a(s_235), .O(gate100inter4));
  nand2 gate2190(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2191(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2192(.a(G31), .O(gate100inter7));
  inv1  gate2193(.a(G353), .O(gate100inter8));
  nand2 gate2194(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2195(.a(s_235), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2196(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2197(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2198(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1527(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1528(.a(gate104inter0), .b(s_140), .O(gate104inter1));
  and2  gate1529(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1530(.a(s_140), .O(gate104inter3));
  inv1  gate1531(.a(s_141), .O(gate104inter4));
  nand2 gate1532(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1533(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1534(.a(G32), .O(gate104inter7));
  inv1  gate1535(.a(G359), .O(gate104inter8));
  nand2 gate1536(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1537(.a(s_141), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1538(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1539(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1540(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1261(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1262(.a(gate105inter0), .b(s_102), .O(gate105inter1));
  and2  gate1263(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1264(.a(s_102), .O(gate105inter3));
  inv1  gate1265(.a(s_103), .O(gate105inter4));
  nand2 gate1266(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1267(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1268(.a(G362), .O(gate105inter7));
  inv1  gate1269(.a(G363), .O(gate105inter8));
  nand2 gate1270(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1271(.a(s_103), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1272(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1273(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1274(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1485(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1486(.a(gate111inter0), .b(s_134), .O(gate111inter1));
  and2  gate1487(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1488(.a(s_134), .O(gate111inter3));
  inv1  gate1489(.a(s_135), .O(gate111inter4));
  nand2 gate1490(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1491(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1492(.a(G374), .O(gate111inter7));
  inv1  gate1493(.a(G375), .O(gate111inter8));
  nand2 gate1494(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1495(.a(s_135), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1496(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1497(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1498(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1051(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1052(.a(gate113inter0), .b(s_72), .O(gate113inter1));
  and2  gate1053(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1054(.a(s_72), .O(gate113inter3));
  inv1  gate1055(.a(s_73), .O(gate113inter4));
  nand2 gate1056(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1057(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1058(.a(G378), .O(gate113inter7));
  inv1  gate1059(.a(G379), .O(gate113inter8));
  nand2 gate1060(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1061(.a(s_73), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1062(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1063(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1064(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1569(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1570(.a(gate115inter0), .b(s_146), .O(gate115inter1));
  and2  gate1571(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1572(.a(s_146), .O(gate115inter3));
  inv1  gate1573(.a(s_147), .O(gate115inter4));
  nand2 gate1574(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1575(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1576(.a(G382), .O(gate115inter7));
  inv1  gate1577(.a(G383), .O(gate115inter8));
  nand2 gate1578(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1579(.a(s_147), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1580(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1581(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1582(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate645(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate646(.a(gate116inter0), .b(s_14), .O(gate116inter1));
  and2  gate647(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate648(.a(s_14), .O(gate116inter3));
  inv1  gate649(.a(s_15), .O(gate116inter4));
  nand2 gate650(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate651(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate652(.a(G384), .O(gate116inter7));
  inv1  gate653(.a(G385), .O(gate116inter8));
  nand2 gate654(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate655(.a(s_15), .b(gate116inter3), .O(gate116inter10));
  nor2  gate656(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate657(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate658(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate2493(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2494(.a(gate117inter0), .b(s_278), .O(gate117inter1));
  and2  gate2495(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2496(.a(s_278), .O(gate117inter3));
  inv1  gate2497(.a(s_279), .O(gate117inter4));
  nand2 gate2498(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2499(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2500(.a(G386), .O(gate117inter7));
  inv1  gate2501(.a(G387), .O(gate117inter8));
  nand2 gate2502(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2503(.a(s_279), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2504(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2505(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2506(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate2787(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2788(.a(gate118inter0), .b(s_320), .O(gate118inter1));
  and2  gate2789(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2790(.a(s_320), .O(gate118inter3));
  inv1  gate2791(.a(s_321), .O(gate118inter4));
  nand2 gate2792(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2793(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2794(.a(G388), .O(gate118inter7));
  inv1  gate2795(.a(G389), .O(gate118inter8));
  nand2 gate2796(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2797(.a(s_321), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2798(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2799(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2800(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate589(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate590(.a(gate120inter0), .b(s_6), .O(gate120inter1));
  and2  gate591(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate592(.a(s_6), .O(gate120inter3));
  inv1  gate593(.a(s_7), .O(gate120inter4));
  nand2 gate594(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate595(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate596(.a(G392), .O(gate120inter7));
  inv1  gate597(.a(G393), .O(gate120inter8));
  nand2 gate598(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate599(.a(s_7), .b(gate120inter3), .O(gate120inter10));
  nor2  gate600(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate601(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate602(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1009(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1010(.a(gate123inter0), .b(s_66), .O(gate123inter1));
  and2  gate1011(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1012(.a(s_66), .O(gate123inter3));
  inv1  gate1013(.a(s_67), .O(gate123inter4));
  nand2 gate1014(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1015(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1016(.a(G398), .O(gate123inter7));
  inv1  gate1017(.a(G399), .O(gate123inter8));
  nand2 gate1018(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1019(.a(s_67), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1020(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1021(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1022(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1499(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1500(.a(gate125inter0), .b(s_136), .O(gate125inter1));
  and2  gate1501(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1502(.a(s_136), .O(gate125inter3));
  inv1  gate1503(.a(s_137), .O(gate125inter4));
  nand2 gate1504(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1505(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1506(.a(G402), .O(gate125inter7));
  inv1  gate1507(.a(G403), .O(gate125inter8));
  nand2 gate1508(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1509(.a(s_137), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1510(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1511(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1512(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate2689(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2690(.a(gate126inter0), .b(s_306), .O(gate126inter1));
  and2  gate2691(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2692(.a(s_306), .O(gate126inter3));
  inv1  gate2693(.a(s_307), .O(gate126inter4));
  nand2 gate2694(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2695(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2696(.a(G404), .O(gate126inter7));
  inv1  gate2697(.a(G405), .O(gate126inter8));
  nand2 gate2698(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2699(.a(s_307), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2700(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2701(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2702(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1877(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1878(.a(gate134inter0), .b(s_190), .O(gate134inter1));
  and2  gate1879(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1880(.a(s_190), .O(gate134inter3));
  inv1  gate1881(.a(s_191), .O(gate134inter4));
  nand2 gate1882(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1883(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1884(.a(G420), .O(gate134inter7));
  inv1  gate1885(.a(G421), .O(gate134inter8));
  nand2 gate1886(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1887(.a(s_191), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1888(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1889(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1890(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2745(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2746(.a(gate136inter0), .b(s_314), .O(gate136inter1));
  and2  gate2747(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2748(.a(s_314), .O(gate136inter3));
  inv1  gate2749(.a(s_315), .O(gate136inter4));
  nand2 gate2750(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2751(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2752(.a(G424), .O(gate136inter7));
  inv1  gate2753(.a(G425), .O(gate136inter8));
  nand2 gate2754(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2755(.a(s_315), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2756(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2757(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2758(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2535(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2536(.a(gate137inter0), .b(s_284), .O(gate137inter1));
  and2  gate2537(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2538(.a(s_284), .O(gate137inter3));
  inv1  gate2539(.a(s_285), .O(gate137inter4));
  nand2 gate2540(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2541(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2542(.a(G426), .O(gate137inter7));
  inv1  gate2543(.a(G429), .O(gate137inter8));
  nand2 gate2544(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2545(.a(s_285), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2546(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2547(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2548(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1765(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1766(.a(gate139inter0), .b(s_174), .O(gate139inter1));
  and2  gate1767(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1768(.a(s_174), .O(gate139inter3));
  inv1  gate1769(.a(s_175), .O(gate139inter4));
  nand2 gate1770(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1771(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1772(.a(G438), .O(gate139inter7));
  inv1  gate1773(.a(G441), .O(gate139inter8));
  nand2 gate1774(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1775(.a(s_175), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1776(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1777(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1778(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1933(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1934(.a(gate140inter0), .b(s_198), .O(gate140inter1));
  and2  gate1935(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1936(.a(s_198), .O(gate140inter3));
  inv1  gate1937(.a(s_199), .O(gate140inter4));
  nand2 gate1938(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1939(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1940(.a(G444), .O(gate140inter7));
  inv1  gate1941(.a(G447), .O(gate140inter8));
  nand2 gate1942(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1943(.a(s_199), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1944(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1945(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1946(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate953(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate954(.a(gate146inter0), .b(s_58), .O(gate146inter1));
  and2  gate955(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate956(.a(s_58), .O(gate146inter3));
  inv1  gate957(.a(s_59), .O(gate146inter4));
  nand2 gate958(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate959(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate960(.a(G480), .O(gate146inter7));
  inv1  gate961(.a(G483), .O(gate146inter8));
  nand2 gate962(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate963(.a(s_59), .b(gate146inter3), .O(gate146inter10));
  nor2  gate964(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate965(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate966(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1807(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1808(.a(gate147inter0), .b(s_180), .O(gate147inter1));
  and2  gate1809(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1810(.a(s_180), .O(gate147inter3));
  inv1  gate1811(.a(s_181), .O(gate147inter4));
  nand2 gate1812(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1813(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1814(.a(G486), .O(gate147inter7));
  inv1  gate1815(.a(G489), .O(gate147inter8));
  nand2 gate1816(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1817(.a(s_181), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1818(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1819(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1820(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate925(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate926(.a(gate149inter0), .b(s_54), .O(gate149inter1));
  and2  gate927(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate928(.a(s_54), .O(gate149inter3));
  inv1  gate929(.a(s_55), .O(gate149inter4));
  nand2 gate930(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate931(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate932(.a(G498), .O(gate149inter7));
  inv1  gate933(.a(G501), .O(gate149inter8));
  nand2 gate934(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate935(.a(s_55), .b(gate149inter3), .O(gate149inter10));
  nor2  gate936(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate937(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate938(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2255(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2256(.a(gate153inter0), .b(s_244), .O(gate153inter1));
  and2  gate2257(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2258(.a(s_244), .O(gate153inter3));
  inv1  gate2259(.a(s_245), .O(gate153inter4));
  nand2 gate2260(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2261(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2262(.a(G426), .O(gate153inter7));
  inv1  gate2263(.a(G522), .O(gate153inter8));
  nand2 gate2264(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2265(.a(s_245), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2266(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2267(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2268(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate603(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate604(.a(gate154inter0), .b(s_8), .O(gate154inter1));
  and2  gate605(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate606(.a(s_8), .O(gate154inter3));
  inv1  gate607(.a(s_9), .O(gate154inter4));
  nand2 gate608(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate609(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate610(.a(G429), .O(gate154inter7));
  inv1  gate611(.a(G522), .O(gate154inter8));
  nand2 gate612(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate613(.a(s_9), .b(gate154inter3), .O(gate154inter10));
  nor2  gate614(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate615(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate616(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2073(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2074(.a(gate156inter0), .b(s_218), .O(gate156inter1));
  and2  gate2075(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2076(.a(s_218), .O(gate156inter3));
  inv1  gate2077(.a(s_219), .O(gate156inter4));
  nand2 gate2078(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2079(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2080(.a(G435), .O(gate156inter7));
  inv1  gate2081(.a(G525), .O(gate156inter8));
  nand2 gate2082(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2083(.a(s_219), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2084(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2085(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2086(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate2311(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2312(.a(gate158inter0), .b(s_252), .O(gate158inter1));
  and2  gate2313(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2314(.a(s_252), .O(gate158inter3));
  inv1  gate2315(.a(s_253), .O(gate158inter4));
  nand2 gate2316(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2317(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2318(.a(G441), .O(gate158inter7));
  inv1  gate2319(.a(G528), .O(gate158inter8));
  nand2 gate2320(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2321(.a(s_253), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2322(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2323(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2324(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1961(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1962(.a(gate165inter0), .b(s_202), .O(gate165inter1));
  and2  gate1963(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1964(.a(s_202), .O(gate165inter3));
  inv1  gate1965(.a(s_203), .O(gate165inter4));
  nand2 gate1966(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1967(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1968(.a(G462), .O(gate165inter7));
  inv1  gate1969(.a(G540), .O(gate165inter8));
  nand2 gate1970(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1971(.a(s_203), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1972(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1973(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1974(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate995(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate996(.a(gate167inter0), .b(s_64), .O(gate167inter1));
  and2  gate997(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate998(.a(s_64), .O(gate167inter3));
  inv1  gate999(.a(s_65), .O(gate167inter4));
  nand2 gate1000(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1001(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1002(.a(G468), .O(gate167inter7));
  inv1  gate1003(.a(G543), .O(gate167inter8));
  nand2 gate1004(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1005(.a(s_65), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1006(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1007(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1008(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1751(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1752(.a(gate174inter0), .b(s_172), .O(gate174inter1));
  and2  gate1753(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1754(.a(s_172), .O(gate174inter3));
  inv1  gate1755(.a(s_173), .O(gate174inter4));
  nand2 gate1756(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1757(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1758(.a(G489), .O(gate174inter7));
  inv1  gate1759(.a(G552), .O(gate174inter8));
  nand2 gate1760(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1761(.a(s_173), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1762(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1763(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1764(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate687(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate688(.a(gate175inter0), .b(s_20), .O(gate175inter1));
  and2  gate689(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate690(.a(s_20), .O(gate175inter3));
  inv1  gate691(.a(s_21), .O(gate175inter4));
  nand2 gate692(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate693(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate694(.a(G492), .O(gate175inter7));
  inv1  gate695(.a(G555), .O(gate175inter8));
  nand2 gate696(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate697(.a(s_21), .b(gate175inter3), .O(gate175inter10));
  nor2  gate698(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate699(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate700(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2381(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2382(.a(gate180inter0), .b(s_262), .O(gate180inter1));
  and2  gate2383(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2384(.a(s_262), .O(gate180inter3));
  inv1  gate2385(.a(s_263), .O(gate180inter4));
  nand2 gate2386(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2387(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2388(.a(G507), .O(gate180inter7));
  inv1  gate2389(.a(G561), .O(gate180inter8));
  nand2 gate2390(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2391(.a(s_263), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2392(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2393(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2394(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1247(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1248(.a(gate181inter0), .b(s_100), .O(gate181inter1));
  and2  gate1249(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1250(.a(s_100), .O(gate181inter3));
  inv1  gate1251(.a(s_101), .O(gate181inter4));
  nand2 gate1252(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1253(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1254(.a(G510), .O(gate181inter7));
  inv1  gate1255(.a(G564), .O(gate181inter8));
  nand2 gate1256(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1257(.a(s_101), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1258(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1259(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1260(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2577(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2578(.a(gate184inter0), .b(s_290), .O(gate184inter1));
  and2  gate2579(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2580(.a(s_290), .O(gate184inter3));
  inv1  gate2581(.a(s_291), .O(gate184inter4));
  nand2 gate2582(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2583(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2584(.a(G519), .O(gate184inter7));
  inv1  gate2585(.a(G567), .O(gate184inter8));
  nand2 gate2586(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2587(.a(s_291), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2588(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2589(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2590(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2353(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2354(.a(gate185inter0), .b(s_258), .O(gate185inter1));
  and2  gate2355(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2356(.a(s_258), .O(gate185inter3));
  inv1  gate2357(.a(s_259), .O(gate185inter4));
  nand2 gate2358(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2359(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2360(.a(G570), .O(gate185inter7));
  inv1  gate2361(.a(G571), .O(gate185inter8));
  nand2 gate2362(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2363(.a(s_259), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2364(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2365(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2366(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2773(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2774(.a(gate186inter0), .b(s_318), .O(gate186inter1));
  and2  gate2775(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2776(.a(s_318), .O(gate186inter3));
  inv1  gate2777(.a(s_319), .O(gate186inter4));
  nand2 gate2778(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2779(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2780(.a(G572), .O(gate186inter7));
  inv1  gate2781(.a(G573), .O(gate186inter8));
  nand2 gate2782(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2783(.a(s_319), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2784(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2785(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2786(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1163(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1164(.a(gate188inter0), .b(s_88), .O(gate188inter1));
  and2  gate1165(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1166(.a(s_88), .O(gate188inter3));
  inv1  gate1167(.a(s_89), .O(gate188inter4));
  nand2 gate1168(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1169(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1170(.a(G576), .O(gate188inter7));
  inv1  gate1171(.a(G577), .O(gate188inter8));
  nand2 gate1172(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1173(.a(s_89), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1174(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1175(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1176(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2437(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2438(.a(gate190inter0), .b(s_270), .O(gate190inter1));
  and2  gate2439(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2440(.a(s_270), .O(gate190inter3));
  inv1  gate2441(.a(s_271), .O(gate190inter4));
  nand2 gate2442(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2443(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2444(.a(G580), .O(gate190inter7));
  inv1  gate2445(.a(G581), .O(gate190inter8));
  nand2 gate2446(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2447(.a(s_271), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2448(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2449(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2450(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1191(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1192(.a(gate195inter0), .b(s_92), .O(gate195inter1));
  and2  gate1193(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1194(.a(s_92), .O(gate195inter3));
  inv1  gate1195(.a(s_93), .O(gate195inter4));
  nand2 gate1196(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1197(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1198(.a(G590), .O(gate195inter7));
  inv1  gate1199(.a(G591), .O(gate195inter8));
  nand2 gate1200(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1201(.a(s_93), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1202(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1203(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1204(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1541(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1542(.a(gate197inter0), .b(s_142), .O(gate197inter1));
  and2  gate1543(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1544(.a(s_142), .O(gate197inter3));
  inv1  gate1545(.a(s_143), .O(gate197inter4));
  nand2 gate1546(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1547(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1548(.a(G594), .O(gate197inter7));
  inv1  gate1549(.a(G595), .O(gate197inter8));
  nand2 gate1550(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1551(.a(s_143), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1552(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1553(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1554(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1723(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1724(.a(gate199inter0), .b(s_168), .O(gate199inter1));
  and2  gate1725(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1726(.a(s_168), .O(gate199inter3));
  inv1  gate1727(.a(s_169), .O(gate199inter4));
  nand2 gate1728(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1729(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1730(.a(G598), .O(gate199inter7));
  inv1  gate1731(.a(G599), .O(gate199inter8));
  nand2 gate1732(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1733(.a(s_169), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1734(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1735(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1736(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1359(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1360(.a(gate204inter0), .b(s_116), .O(gate204inter1));
  and2  gate1361(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1362(.a(s_116), .O(gate204inter3));
  inv1  gate1363(.a(s_117), .O(gate204inter4));
  nand2 gate1364(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1365(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1366(.a(G607), .O(gate204inter7));
  inv1  gate1367(.a(G617), .O(gate204inter8));
  nand2 gate1368(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1369(.a(s_117), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1370(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1371(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1372(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate2633(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2634(.a(gate205inter0), .b(s_298), .O(gate205inter1));
  and2  gate2635(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2636(.a(s_298), .O(gate205inter3));
  inv1  gate2637(.a(s_299), .O(gate205inter4));
  nand2 gate2638(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2639(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2640(.a(G622), .O(gate205inter7));
  inv1  gate2641(.a(G627), .O(gate205inter8));
  nand2 gate2642(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2643(.a(s_299), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2644(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2645(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2646(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2479(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2480(.a(gate206inter0), .b(s_276), .O(gate206inter1));
  and2  gate2481(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2482(.a(s_276), .O(gate206inter3));
  inv1  gate2483(.a(s_277), .O(gate206inter4));
  nand2 gate2484(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2485(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2486(.a(G632), .O(gate206inter7));
  inv1  gate2487(.a(G637), .O(gate206inter8));
  nand2 gate2488(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2489(.a(s_277), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2490(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2491(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2492(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1863(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1864(.a(gate210inter0), .b(s_188), .O(gate210inter1));
  and2  gate1865(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1866(.a(s_188), .O(gate210inter3));
  inv1  gate1867(.a(s_189), .O(gate210inter4));
  nand2 gate1868(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1869(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1870(.a(G607), .O(gate210inter7));
  inv1  gate1871(.a(G666), .O(gate210inter8));
  nand2 gate1872(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1873(.a(s_189), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1874(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1875(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1876(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1317(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1318(.a(gate214inter0), .b(s_110), .O(gate214inter1));
  and2  gate1319(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1320(.a(s_110), .O(gate214inter3));
  inv1  gate1321(.a(s_111), .O(gate214inter4));
  nand2 gate1322(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1323(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1324(.a(G612), .O(gate214inter7));
  inv1  gate1325(.a(G672), .O(gate214inter8));
  nand2 gate1326(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1327(.a(s_111), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1328(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1329(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1330(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2129(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2130(.a(gate215inter0), .b(s_226), .O(gate215inter1));
  and2  gate2131(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2132(.a(s_226), .O(gate215inter3));
  inv1  gate2133(.a(s_227), .O(gate215inter4));
  nand2 gate2134(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2135(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2136(.a(G607), .O(gate215inter7));
  inv1  gate2137(.a(G675), .O(gate215inter8));
  nand2 gate2138(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2139(.a(s_227), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2140(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2141(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2142(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate785(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate786(.a(gate216inter0), .b(s_34), .O(gate216inter1));
  and2  gate787(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate788(.a(s_34), .O(gate216inter3));
  inv1  gate789(.a(s_35), .O(gate216inter4));
  nand2 gate790(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate791(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate792(.a(G617), .O(gate216inter7));
  inv1  gate793(.a(G675), .O(gate216inter8));
  nand2 gate794(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate795(.a(s_35), .b(gate216inter3), .O(gate216inter10));
  nor2  gate796(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate797(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate798(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2843(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2844(.a(gate217inter0), .b(s_328), .O(gate217inter1));
  and2  gate2845(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2846(.a(s_328), .O(gate217inter3));
  inv1  gate2847(.a(s_329), .O(gate217inter4));
  nand2 gate2848(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2849(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2850(.a(G622), .O(gate217inter7));
  inv1  gate2851(.a(G678), .O(gate217inter8));
  nand2 gate2852(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2853(.a(s_329), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2854(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2855(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2856(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1667(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1668(.a(gate223inter0), .b(s_160), .O(gate223inter1));
  and2  gate1669(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1670(.a(s_160), .O(gate223inter3));
  inv1  gate1671(.a(s_161), .O(gate223inter4));
  nand2 gate1672(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1673(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1674(.a(G627), .O(gate223inter7));
  inv1  gate1675(.a(G687), .O(gate223inter8));
  nand2 gate1676(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1677(.a(s_161), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1678(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1679(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1680(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1093(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1094(.a(gate225inter0), .b(s_78), .O(gate225inter1));
  and2  gate1095(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1096(.a(s_78), .O(gate225inter3));
  inv1  gate1097(.a(s_79), .O(gate225inter4));
  nand2 gate1098(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1099(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1100(.a(G690), .O(gate225inter7));
  inv1  gate1101(.a(G691), .O(gate225inter8));
  nand2 gate1102(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1103(.a(s_79), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1104(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1105(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1106(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate743(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate744(.a(gate226inter0), .b(s_28), .O(gate226inter1));
  and2  gate745(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate746(.a(s_28), .O(gate226inter3));
  inv1  gate747(.a(s_29), .O(gate226inter4));
  nand2 gate748(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate749(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate750(.a(G692), .O(gate226inter7));
  inv1  gate751(.a(G693), .O(gate226inter8));
  nand2 gate752(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate753(.a(s_29), .b(gate226inter3), .O(gate226inter10));
  nor2  gate754(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate755(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate756(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1779(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1780(.a(gate227inter0), .b(s_176), .O(gate227inter1));
  and2  gate1781(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1782(.a(s_176), .O(gate227inter3));
  inv1  gate1783(.a(s_177), .O(gate227inter4));
  nand2 gate1784(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1785(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1786(.a(G694), .O(gate227inter7));
  inv1  gate1787(.a(G695), .O(gate227inter8));
  nand2 gate1788(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1789(.a(s_177), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1790(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1791(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1792(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2703(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2704(.a(gate229inter0), .b(s_308), .O(gate229inter1));
  and2  gate2705(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2706(.a(s_308), .O(gate229inter3));
  inv1  gate2707(.a(s_309), .O(gate229inter4));
  nand2 gate2708(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2709(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2710(.a(G698), .O(gate229inter7));
  inv1  gate2711(.a(G699), .O(gate229inter8));
  nand2 gate2712(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2713(.a(s_309), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2714(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2715(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2716(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1289(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1290(.a(gate230inter0), .b(s_106), .O(gate230inter1));
  and2  gate1291(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1292(.a(s_106), .O(gate230inter3));
  inv1  gate1293(.a(s_107), .O(gate230inter4));
  nand2 gate1294(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1295(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1296(.a(G700), .O(gate230inter7));
  inv1  gate1297(.a(G701), .O(gate230inter8));
  nand2 gate1298(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1299(.a(s_107), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1300(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1301(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1302(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate897(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate898(.a(gate231inter0), .b(s_50), .O(gate231inter1));
  and2  gate899(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate900(.a(s_50), .O(gate231inter3));
  inv1  gate901(.a(s_51), .O(gate231inter4));
  nand2 gate902(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate903(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate904(.a(G702), .O(gate231inter7));
  inv1  gate905(.a(G703), .O(gate231inter8));
  nand2 gate906(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate907(.a(s_51), .b(gate231inter3), .O(gate231inter10));
  nor2  gate908(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate909(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate910(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate855(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate856(.a(gate232inter0), .b(s_44), .O(gate232inter1));
  and2  gate857(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate858(.a(s_44), .O(gate232inter3));
  inv1  gate859(.a(s_45), .O(gate232inter4));
  nand2 gate860(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate861(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate862(.a(G704), .O(gate232inter7));
  inv1  gate863(.a(G705), .O(gate232inter8));
  nand2 gate864(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate865(.a(s_45), .b(gate232inter3), .O(gate232inter10));
  nor2  gate866(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate867(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate868(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1121(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1122(.a(gate233inter0), .b(s_82), .O(gate233inter1));
  and2  gate1123(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1124(.a(s_82), .O(gate233inter3));
  inv1  gate1125(.a(s_83), .O(gate233inter4));
  nand2 gate1126(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1127(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1128(.a(G242), .O(gate233inter7));
  inv1  gate1129(.a(G718), .O(gate233inter8));
  nand2 gate1130(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1131(.a(s_83), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1132(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1133(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1134(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2171(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2172(.a(gate240inter0), .b(s_232), .O(gate240inter1));
  and2  gate2173(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2174(.a(s_232), .O(gate240inter3));
  inv1  gate2175(.a(s_233), .O(gate240inter4));
  nand2 gate2176(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2177(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2178(.a(G263), .O(gate240inter7));
  inv1  gate2179(.a(G715), .O(gate240inter8));
  nand2 gate2180(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2181(.a(s_233), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2182(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2183(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2184(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate771(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate772(.a(gate243inter0), .b(s_32), .O(gate243inter1));
  and2  gate773(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate774(.a(s_32), .O(gate243inter3));
  inv1  gate775(.a(s_33), .O(gate243inter4));
  nand2 gate776(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate777(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate778(.a(G245), .O(gate243inter7));
  inv1  gate779(.a(G733), .O(gate243inter8));
  nand2 gate780(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate781(.a(s_33), .b(gate243inter3), .O(gate243inter10));
  nor2  gate782(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate783(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate784(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2017(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2018(.a(gate250inter0), .b(s_210), .O(gate250inter1));
  and2  gate2019(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2020(.a(s_210), .O(gate250inter3));
  inv1  gate2021(.a(s_211), .O(gate250inter4));
  nand2 gate2022(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2023(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2024(.a(G706), .O(gate250inter7));
  inv1  gate2025(.a(G742), .O(gate250inter8));
  nand2 gate2026(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2027(.a(s_211), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2028(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2029(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2030(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2241(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2242(.a(gate251inter0), .b(s_242), .O(gate251inter1));
  and2  gate2243(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2244(.a(s_242), .O(gate251inter3));
  inv1  gate2245(.a(s_243), .O(gate251inter4));
  nand2 gate2246(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2247(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2248(.a(G257), .O(gate251inter7));
  inv1  gate2249(.a(G745), .O(gate251inter8));
  nand2 gate2250(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2251(.a(s_243), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2252(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2253(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2254(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate617(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate618(.a(gate253inter0), .b(s_10), .O(gate253inter1));
  and2  gate619(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate620(.a(s_10), .O(gate253inter3));
  inv1  gate621(.a(s_11), .O(gate253inter4));
  nand2 gate622(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate623(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate624(.a(G260), .O(gate253inter7));
  inv1  gate625(.a(G748), .O(gate253inter8));
  nand2 gate626(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate627(.a(s_11), .b(gate253inter3), .O(gate253inter10));
  nor2  gate628(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate629(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate630(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1373(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1374(.a(gate254inter0), .b(s_118), .O(gate254inter1));
  and2  gate1375(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1376(.a(s_118), .O(gate254inter3));
  inv1  gate1377(.a(s_119), .O(gate254inter4));
  nand2 gate1378(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1379(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1380(.a(G712), .O(gate254inter7));
  inv1  gate1381(.a(G748), .O(gate254inter8));
  nand2 gate1382(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1383(.a(s_119), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1384(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1385(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1386(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1989(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1990(.a(gate256inter0), .b(s_206), .O(gate256inter1));
  and2  gate1991(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1992(.a(s_206), .O(gate256inter3));
  inv1  gate1993(.a(s_207), .O(gate256inter4));
  nand2 gate1994(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1995(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1996(.a(G715), .O(gate256inter7));
  inv1  gate1997(.a(G751), .O(gate256inter8));
  nand2 gate1998(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1999(.a(s_207), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2000(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2001(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2002(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2283(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2284(.a(gate258inter0), .b(s_248), .O(gate258inter1));
  and2  gate2285(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2286(.a(s_248), .O(gate258inter3));
  inv1  gate2287(.a(s_249), .O(gate258inter4));
  nand2 gate2288(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2289(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2290(.a(G756), .O(gate258inter7));
  inv1  gate2291(.a(G757), .O(gate258inter8));
  nand2 gate2292(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2293(.a(s_249), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2294(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2295(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2296(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1429(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1430(.a(gate262inter0), .b(s_126), .O(gate262inter1));
  and2  gate1431(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1432(.a(s_126), .O(gate262inter3));
  inv1  gate1433(.a(s_127), .O(gate262inter4));
  nand2 gate1434(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1435(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1436(.a(G764), .O(gate262inter7));
  inv1  gate1437(.a(G765), .O(gate262inter8));
  nand2 gate1438(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1439(.a(s_127), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1440(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1441(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1442(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1597(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1598(.a(gate264inter0), .b(s_150), .O(gate264inter1));
  and2  gate1599(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1600(.a(s_150), .O(gate264inter3));
  inv1  gate1601(.a(s_151), .O(gate264inter4));
  nand2 gate1602(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1603(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1604(.a(G768), .O(gate264inter7));
  inv1  gate1605(.a(G769), .O(gate264inter8));
  nand2 gate1606(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1607(.a(s_151), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1608(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1609(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1610(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate631(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate632(.a(gate266inter0), .b(s_12), .O(gate266inter1));
  and2  gate633(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate634(.a(s_12), .O(gate266inter3));
  inv1  gate635(.a(s_13), .O(gate266inter4));
  nand2 gate636(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate637(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate638(.a(G645), .O(gate266inter7));
  inv1  gate639(.a(G773), .O(gate266inter8));
  nand2 gate640(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate641(.a(s_13), .b(gate266inter3), .O(gate266inter10));
  nor2  gate642(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate643(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate644(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2759(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2760(.a(gate267inter0), .b(s_316), .O(gate267inter1));
  and2  gate2761(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2762(.a(s_316), .O(gate267inter3));
  inv1  gate2763(.a(s_317), .O(gate267inter4));
  nand2 gate2764(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2765(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2766(.a(G648), .O(gate267inter7));
  inv1  gate2767(.a(G776), .O(gate267inter8));
  nand2 gate2768(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2769(.a(s_317), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2770(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2771(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2772(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1219(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1220(.a(gate271inter0), .b(s_96), .O(gate271inter1));
  and2  gate1221(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1222(.a(s_96), .O(gate271inter3));
  inv1  gate1223(.a(s_97), .O(gate271inter4));
  nand2 gate1224(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1225(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1226(.a(G660), .O(gate271inter7));
  inv1  gate1227(.a(G788), .O(gate271inter8));
  nand2 gate1228(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1229(.a(s_97), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1230(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1231(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1232(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2269(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2270(.a(gate272inter0), .b(s_246), .O(gate272inter1));
  and2  gate2271(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2272(.a(s_246), .O(gate272inter3));
  inv1  gate2273(.a(s_247), .O(gate272inter4));
  nand2 gate2274(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2275(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2276(.a(G663), .O(gate272inter7));
  inv1  gate2277(.a(G791), .O(gate272inter8));
  nand2 gate2278(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2279(.a(s_247), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2280(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2281(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2282(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1401(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1402(.a(gate275inter0), .b(s_122), .O(gate275inter1));
  and2  gate1403(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1404(.a(s_122), .O(gate275inter3));
  inv1  gate1405(.a(s_123), .O(gate275inter4));
  nand2 gate1406(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1407(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1408(.a(G645), .O(gate275inter7));
  inv1  gate1409(.a(G797), .O(gate275inter8));
  nand2 gate1410(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1411(.a(s_123), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1412(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1413(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1414(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2367(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2368(.a(gate278inter0), .b(s_260), .O(gate278inter1));
  and2  gate2369(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2370(.a(s_260), .O(gate278inter3));
  inv1  gate2371(.a(s_261), .O(gate278inter4));
  nand2 gate2372(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2373(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2374(.a(G776), .O(gate278inter7));
  inv1  gate2375(.a(G800), .O(gate278inter8));
  nand2 gate2376(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2377(.a(s_261), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2378(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2379(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2380(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1625(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1626(.a(gate282inter0), .b(s_154), .O(gate282inter1));
  and2  gate1627(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1628(.a(s_154), .O(gate282inter3));
  inv1  gate1629(.a(s_155), .O(gate282inter4));
  nand2 gate1630(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1631(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1632(.a(G782), .O(gate282inter7));
  inv1  gate1633(.a(G806), .O(gate282inter8));
  nand2 gate1634(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1635(.a(s_155), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1636(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1637(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1638(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1177(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1178(.a(gate283inter0), .b(s_90), .O(gate283inter1));
  and2  gate1179(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1180(.a(s_90), .O(gate283inter3));
  inv1  gate1181(.a(s_91), .O(gate283inter4));
  nand2 gate1182(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1183(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1184(.a(G657), .O(gate283inter7));
  inv1  gate1185(.a(G809), .O(gate283inter8));
  nand2 gate1186(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1187(.a(s_91), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1188(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1189(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1190(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate715(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate716(.a(gate284inter0), .b(s_24), .O(gate284inter1));
  and2  gate717(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate718(.a(s_24), .O(gate284inter3));
  inv1  gate719(.a(s_25), .O(gate284inter4));
  nand2 gate720(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate721(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate722(.a(G785), .O(gate284inter7));
  inv1  gate723(.a(G809), .O(gate284inter8));
  nand2 gate724(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate725(.a(s_25), .b(gate284inter3), .O(gate284inter10));
  nor2  gate726(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate727(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate728(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1065(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1066(.a(gate287inter0), .b(s_74), .O(gate287inter1));
  and2  gate1067(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1068(.a(s_74), .O(gate287inter3));
  inv1  gate1069(.a(s_75), .O(gate287inter4));
  nand2 gate1070(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1071(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1072(.a(G663), .O(gate287inter7));
  inv1  gate1073(.a(G815), .O(gate287inter8));
  nand2 gate1074(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1075(.a(s_75), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1076(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1077(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1078(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1653(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1654(.a(gate295inter0), .b(s_158), .O(gate295inter1));
  and2  gate1655(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1656(.a(s_158), .O(gate295inter3));
  inv1  gate1657(.a(s_159), .O(gate295inter4));
  nand2 gate1658(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1659(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1660(.a(G830), .O(gate295inter7));
  inv1  gate1661(.a(G831), .O(gate295inter8));
  nand2 gate1662(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1663(.a(s_159), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1664(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1665(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1666(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1695(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1696(.a(gate389inter0), .b(s_164), .O(gate389inter1));
  and2  gate1697(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1698(.a(s_164), .O(gate389inter3));
  inv1  gate1699(.a(s_165), .O(gate389inter4));
  nand2 gate1700(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1701(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1702(.a(G3), .O(gate389inter7));
  inv1  gate1703(.a(G1042), .O(gate389inter8));
  nand2 gate1704(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1705(.a(s_165), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1706(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1707(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1708(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate981(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate982(.a(gate390inter0), .b(s_62), .O(gate390inter1));
  and2  gate983(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate984(.a(s_62), .O(gate390inter3));
  inv1  gate985(.a(s_63), .O(gate390inter4));
  nand2 gate986(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate987(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate988(.a(G4), .O(gate390inter7));
  inv1  gate989(.a(G1045), .O(gate390inter8));
  nand2 gate990(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate991(.a(s_63), .b(gate390inter3), .O(gate390inter10));
  nor2  gate992(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate993(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate994(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1513(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1514(.a(gate391inter0), .b(s_138), .O(gate391inter1));
  and2  gate1515(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1516(.a(s_138), .O(gate391inter3));
  inv1  gate1517(.a(s_139), .O(gate391inter4));
  nand2 gate1518(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1519(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1520(.a(G5), .O(gate391inter7));
  inv1  gate1521(.a(G1048), .O(gate391inter8));
  nand2 gate1522(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1523(.a(s_139), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1524(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1525(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1526(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2521(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2522(.a(gate394inter0), .b(s_282), .O(gate394inter1));
  and2  gate2523(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2524(.a(s_282), .O(gate394inter3));
  inv1  gate2525(.a(s_283), .O(gate394inter4));
  nand2 gate2526(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2527(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2528(.a(G8), .O(gate394inter7));
  inv1  gate2529(.a(G1057), .O(gate394inter8));
  nand2 gate2530(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2531(.a(s_283), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2532(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2533(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2534(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1149(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1150(.a(gate397inter0), .b(s_86), .O(gate397inter1));
  and2  gate1151(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1152(.a(s_86), .O(gate397inter3));
  inv1  gate1153(.a(s_87), .O(gate397inter4));
  nand2 gate1154(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1155(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1156(.a(G11), .O(gate397inter7));
  inv1  gate1157(.a(G1066), .O(gate397inter8));
  nand2 gate1158(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1159(.a(s_87), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1160(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1161(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1162(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1709(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1710(.a(gate399inter0), .b(s_166), .O(gate399inter1));
  and2  gate1711(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1712(.a(s_166), .O(gate399inter3));
  inv1  gate1713(.a(s_167), .O(gate399inter4));
  nand2 gate1714(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1715(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1716(.a(G13), .O(gate399inter7));
  inv1  gate1717(.a(G1072), .O(gate399inter8));
  nand2 gate1718(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1719(.a(s_167), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1720(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1721(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1722(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1345(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1346(.a(gate403inter0), .b(s_114), .O(gate403inter1));
  and2  gate1347(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1348(.a(s_114), .O(gate403inter3));
  inv1  gate1349(.a(s_115), .O(gate403inter4));
  nand2 gate1350(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1351(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1352(.a(G17), .O(gate403inter7));
  inv1  gate1353(.a(G1084), .O(gate403inter8));
  nand2 gate1354(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1355(.a(s_115), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1356(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1357(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1358(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate659(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate660(.a(gate405inter0), .b(s_16), .O(gate405inter1));
  and2  gate661(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate662(.a(s_16), .O(gate405inter3));
  inv1  gate663(.a(s_17), .O(gate405inter4));
  nand2 gate664(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate665(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate666(.a(G19), .O(gate405inter7));
  inv1  gate667(.a(G1090), .O(gate405inter8));
  nand2 gate668(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate669(.a(s_17), .b(gate405inter3), .O(gate405inter10));
  nor2  gate670(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate671(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate672(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate547(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate548(.a(gate407inter0), .b(s_0), .O(gate407inter1));
  and2  gate549(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate550(.a(s_0), .O(gate407inter3));
  inv1  gate551(.a(s_1), .O(gate407inter4));
  nand2 gate552(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate553(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate554(.a(G21), .O(gate407inter7));
  inv1  gate555(.a(G1096), .O(gate407inter8));
  nand2 gate556(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate557(.a(s_1), .b(gate407inter3), .O(gate407inter10));
  nor2  gate558(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate559(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate560(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate2801(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2802(.a(gate408inter0), .b(s_322), .O(gate408inter1));
  and2  gate2803(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2804(.a(s_322), .O(gate408inter3));
  inv1  gate2805(.a(s_323), .O(gate408inter4));
  nand2 gate2806(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2807(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2808(.a(G22), .O(gate408inter7));
  inv1  gate2809(.a(G1099), .O(gate408inter8));
  nand2 gate2810(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2811(.a(s_323), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2812(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2813(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2814(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate799(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate800(.a(gate413inter0), .b(s_36), .O(gate413inter1));
  and2  gate801(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate802(.a(s_36), .O(gate413inter3));
  inv1  gate803(.a(s_37), .O(gate413inter4));
  nand2 gate804(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate805(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate806(.a(G27), .O(gate413inter7));
  inv1  gate807(.a(G1114), .O(gate413inter8));
  nand2 gate808(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate809(.a(s_37), .b(gate413inter3), .O(gate413inter10));
  nor2  gate810(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate811(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate812(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate561(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate562(.a(gate415inter0), .b(s_2), .O(gate415inter1));
  and2  gate563(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate564(.a(s_2), .O(gate415inter3));
  inv1  gate565(.a(s_3), .O(gate415inter4));
  nand2 gate566(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate567(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate568(.a(G29), .O(gate415inter7));
  inv1  gate569(.a(G1120), .O(gate415inter8));
  nand2 gate570(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate571(.a(s_3), .b(gate415inter3), .O(gate415inter10));
  nor2  gate572(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate573(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate574(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1387(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1388(.a(gate418inter0), .b(s_120), .O(gate418inter1));
  and2  gate1389(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1390(.a(s_120), .O(gate418inter3));
  inv1  gate1391(.a(s_121), .O(gate418inter4));
  nand2 gate1392(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1393(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1394(.a(G32), .O(gate418inter7));
  inv1  gate1395(.a(G1129), .O(gate418inter8));
  nand2 gate1396(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1397(.a(s_121), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1398(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1399(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1400(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2199(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2200(.a(gate420inter0), .b(s_236), .O(gate420inter1));
  and2  gate2201(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2202(.a(s_236), .O(gate420inter3));
  inv1  gate2203(.a(s_237), .O(gate420inter4));
  nand2 gate2204(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2205(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2206(.a(G1036), .O(gate420inter7));
  inv1  gate2207(.a(G1132), .O(gate420inter8));
  nand2 gate2208(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2209(.a(s_237), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2210(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2211(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2212(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2003(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2004(.a(gate423inter0), .b(s_208), .O(gate423inter1));
  and2  gate2005(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2006(.a(s_208), .O(gate423inter3));
  inv1  gate2007(.a(s_209), .O(gate423inter4));
  nand2 gate2008(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2009(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2010(.a(G3), .O(gate423inter7));
  inv1  gate2011(.a(G1138), .O(gate423inter8));
  nand2 gate2012(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2013(.a(s_209), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2014(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2015(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2016(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate869(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate870(.a(gate424inter0), .b(s_46), .O(gate424inter1));
  and2  gate871(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate872(.a(s_46), .O(gate424inter3));
  inv1  gate873(.a(s_47), .O(gate424inter4));
  nand2 gate874(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate875(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate876(.a(G1042), .O(gate424inter7));
  inv1  gate877(.a(G1138), .O(gate424inter8));
  nand2 gate878(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate879(.a(s_47), .b(gate424inter3), .O(gate424inter10));
  nor2  gate880(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate881(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate882(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate813(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate814(.a(gate426inter0), .b(s_38), .O(gate426inter1));
  and2  gate815(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate816(.a(s_38), .O(gate426inter3));
  inv1  gate817(.a(s_39), .O(gate426inter4));
  nand2 gate818(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate819(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate820(.a(G1045), .O(gate426inter7));
  inv1  gate821(.a(G1141), .O(gate426inter8));
  nand2 gate822(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate823(.a(s_39), .b(gate426inter3), .O(gate426inter10));
  nor2  gate824(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate825(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate826(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2325(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2326(.a(gate428inter0), .b(s_254), .O(gate428inter1));
  and2  gate2327(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2328(.a(s_254), .O(gate428inter3));
  inv1  gate2329(.a(s_255), .O(gate428inter4));
  nand2 gate2330(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2331(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2332(.a(G1048), .O(gate428inter7));
  inv1  gate2333(.a(G1144), .O(gate428inter8));
  nand2 gate2334(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2335(.a(s_255), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2336(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2337(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2338(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1079(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1080(.a(gate430inter0), .b(s_76), .O(gate430inter1));
  and2  gate1081(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1082(.a(s_76), .O(gate430inter3));
  inv1  gate1083(.a(s_77), .O(gate430inter4));
  nand2 gate1084(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1085(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1086(.a(G1051), .O(gate430inter7));
  inv1  gate1087(.a(G1147), .O(gate430inter8));
  nand2 gate1088(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1089(.a(s_77), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1090(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1091(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1092(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2395(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2396(.a(gate431inter0), .b(s_264), .O(gate431inter1));
  and2  gate2397(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2398(.a(s_264), .O(gate431inter3));
  inv1  gate2399(.a(s_265), .O(gate431inter4));
  nand2 gate2400(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2401(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2402(.a(G7), .O(gate431inter7));
  inv1  gate2403(.a(G1150), .O(gate431inter8));
  nand2 gate2404(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2405(.a(s_265), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2406(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2407(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2408(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate729(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate730(.a(gate432inter0), .b(s_26), .O(gate432inter1));
  and2  gate731(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate732(.a(s_26), .O(gate432inter3));
  inv1  gate733(.a(s_27), .O(gate432inter4));
  nand2 gate734(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate735(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate736(.a(G1054), .O(gate432inter7));
  inv1  gate737(.a(G1150), .O(gate432inter8));
  nand2 gate738(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate739(.a(s_27), .b(gate432inter3), .O(gate432inter10));
  nor2  gate740(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate741(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate742(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1023(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1024(.a(gate435inter0), .b(s_68), .O(gate435inter1));
  and2  gate1025(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1026(.a(s_68), .O(gate435inter3));
  inv1  gate1027(.a(s_69), .O(gate435inter4));
  nand2 gate1028(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1029(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1030(.a(G9), .O(gate435inter7));
  inv1  gate1031(.a(G1156), .O(gate435inter8));
  nand2 gate1032(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1033(.a(s_69), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1034(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1035(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1036(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1303(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1304(.a(gate438inter0), .b(s_108), .O(gate438inter1));
  and2  gate1305(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1306(.a(s_108), .O(gate438inter3));
  inv1  gate1307(.a(s_109), .O(gate438inter4));
  nand2 gate1308(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1309(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1310(.a(G1063), .O(gate438inter7));
  inv1  gate1311(.a(G1159), .O(gate438inter8));
  nand2 gate1312(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1313(.a(s_109), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1314(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1315(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1316(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate575(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate576(.a(gate439inter0), .b(s_4), .O(gate439inter1));
  and2  gate577(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate578(.a(s_4), .O(gate439inter3));
  inv1  gate579(.a(s_5), .O(gate439inter4));
  nand2 gate580(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate581(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate582(.a(G11), .O(gate439inter7));
  inv1  gate583(.a(G1162), .O(gate439inter8));
  nand2 gate584(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate585(.a(s_5), .b(gate439inter3), .O(gate439inter10));
  nor2  gate586(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate587(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate588(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1891(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1892(.a(gate444inter0), .b(s_192), .O(gate444inter1));
  and2  gate1893(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1894(.a(s_192), .O(gate444inter3));
  inv1  gate1895(.a(s_193), .O(gate444inter4));
  nand2 gate1896(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1897(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1898(.a(G1072), .O(gate444inter7));
  inv1  gate1899(.a(G1168), .O(gate444inter8));
  nand2 gate1900(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1901(.a(s_193), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1902(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1903(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1904(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2409(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2410(.a(gate448inter0), .b(s_266), .O(gate448inter1));
  and2  gate2411(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2412(.a(s_266), .O(gate448inter3));
  inv1  gate2413(.a(s_267), .O(gate448inter4));
  nand2 gate2414(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2415(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2416(.a(G1078), .O(gate448inter7));
  inv1  gate2417(.a(G1174), .O(gate448inter8));
  nand2 gate2418(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2419(.a(s_267), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2420(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2421(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2422(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1555(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1556(.a(gate449inter0), .b(s_144), .O(gate449inter1));
  and2  gate1557(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1558(.a(s_144), .O(gate449inter3));
  inv1  gate1559(.a(s_145), .O(gate449inter4));
  nand2 gate1560(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1561(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1562(.a(G16), .O(gate449inter7));
  inv1  gate1563(.a(G1177), .O(gate449inter8));
  nand2 gate1564(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1565(.a(s_145), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1566(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1567(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1568(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate939(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate940(.a(gate450inter0), .b(s_56), .O(gate450inter1));
  and2  gate941(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate942(.a(s_56), .O(gate450inter3));
  inv1  gate943(.a(s_57), .O(gate450inter4));
  nand2 gate944(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate945(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate946(.a(G1081), .O(gate450inter7));
  inv1  gate947(.a(G1177), .O(gate450inter8));
  nand2 gate948(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate949(.a(s_57), .b(gate450inter3), .O(gate450inter10));
  nor2  gate950(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate951(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate952(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1415(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1416(.a(gate451inter0), .b(s_124), .O(gate451inter1));
  and2  gate1417(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1418(.a(s_124), .O(gate451inter3));
  inv1  gate1419(.a(s_125), .O(gate451inter4));
  nand2 gate1420(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1421(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1422(.a(G17), .O(gate451inter7));
  inv1  gate1423(.a(G1180), .O(gate451inter8));
  nand2 gate1424(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1425(.a(s_125), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1426(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1427(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1428(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2115(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2116(.a(gate453inter0), .b(s_224), .O(gate453inter1));
  and2  gate2117(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2118(.a(s_224), .O(gate453inter3));
  inv1  gate2119(.a(s_225), .O(gate453inter4));
  nand2 gate2120(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2121(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2122(.a(G18), .O(gate453inter7));
  inv1  gate2123(.a(G1183), .O(gate453inter8));
  nand2 gate2124(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2125(.a(s_225), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2126(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2127(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2128(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1583(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1584(.a(gate458inter0), .b(s_148), .O(gate458inter1));
  and2  gate1585(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1586(.a(s_148), .O(gate458inter3));
  inv1  gate1587(.a(s_149), .O(gate458inter4));
  nand2 gate1588(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1589(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1590(.a(G1093), .O(gate458inter7));
  inv1  gate1591(.a(G1189), .O(gate458inter8));
  nand2 gate1592(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1593(.a(s_149), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1594(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1595(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1596(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate883(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate884(.a(gate460inter0), .b(s_48), .O(gate460inter1));
  and2  gate885(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate886(.a(s_48), .O(gate460inter3));
  inv1  gate887(.a(s_49), .O(gate460inter4));
  nand2 gate888(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate889(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate890(.a(G1096), .O(gate460inter7));
  inv1  gate891(.a(G1192), .O(gate460inter8));
  nand2 gate892(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate893(.a(s_49), .b(gate460inter3), .O(gate460inter10));
  nor2  gate894(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate895(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate896(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2045(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2046(.a(gate462inter0), .b(s_214), .O(gate462inter1));
  and2  gate2047(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2048(.a(s_214), .O(gate462inter3));
  inv1  gate2049(.a(s_215), .O(gate462inter4));
  nand2 gate2050(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2051(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2052(.a(G1099), .O(gate462inter7));
  inv1  gate2053(.a(G1195), .O(gate462inter8));
  nand2 gate2054(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2055(.a(s_215), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2056(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2057(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2058(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1639(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1640(.a(gate464inter0), .b(s_156), .O(gate464inter1));
  and2  gate1641(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1642(.a(s_156), .O(gate464inter3));
  inv1  gate1643(.a(s_157), .O(gate464inter4));
  nand2 gate1644(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1645(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1646(.a(G1102), .O(gate464inter7));
  inv1  gate1647(.a(G1198), .O(gate464inter8));
  nand2 gate1648(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1649(.a(s_157), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1650(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1651(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1652(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate967(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate968(.a(gate465inter0), .b(s_60), .O(gate465inter1));
  and2  gate969(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate970(.a(s_60), .O(gate465inter3));
  inv1  gate971(.a(s_61), .O(gate465inter4));
  nand2 gate972(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate973(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate974(.a(G24), .O(gate465inter7));
  inv1  gate975(.a(G1201), .O(gate465inter8));
  nand2 gate976(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate977(.a(s_61), .b(gate465inter3), .O(gate465inter10));
  nor2  gate978(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate979(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate980(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2591(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2592(.a(gate466inter0), .b(s_292), .O(gate466inter1));
  and2  gate2593(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2594(.a(s_292), .O(gate466inter3));
  inv1  gate2595(.a(s_293), .O(gate466inter4));
  nand2 gate2596(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2597(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2598(.a(G1105), .O(gate466inter7));
  inv1  gate2599(.a(G1201), .O(gate466inter8));
  nand2 gate2600(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2601(.a(s_293), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2602(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2603(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2604(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2829(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2830(.a(gate470inter0), .b(s_326), .O(gate470inter1));
  and2  gate2831(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2832(.a(s_326), .O(gate470inter3));
  inv1  gate2833(.a(s_327), .O(gate470inter4));
  nand2 gate2834(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2835(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2836(.a(G1111), .O(gate470inter7));
  inv1  gate2837(.a(G1207), .O(gate470inter8));
  nand2 gate2838(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2839(.a(s_327), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2840(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2841(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2842(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2465(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2466(.a(gate475inter0), .b(s_274), .O(gate475inter1));
  and2  gate2467(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2468(.a(s_274), .O(gate475inter3));
  inv1  gate2469(.a(s_275), .O(gate475inter4));
  nand2 gate2470(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2471(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2472(.a(G29), .O(gate475inter7));
  inv1  gate2473(.a(G1216), .O(gate475inter8));
  nand2 gate2474(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2475(.a(s_275), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2476(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2477(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2478(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1975(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1976(.a(gate483inter0), .b(s_204), .O(gate483inter1));
  and2  gate1977(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1978(.a(s_204), .O(gate483inter3));
  inv1  gate1979(.a(s_205), .O(gate483inter4));
  nand2 gate1980(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1981(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1982(.a(G1228), .O(gate483inter7));
  inv1  gate1983(.a(G1229), .O(gate483inter8));
  nand2 gate1984(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1985(.a(s_205), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1986(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1987(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1988(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2031(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2032(.a(gate486inter0), .b(s_212), .O(gate486inter1));
  and2  gate2033(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2034(.a(s_212), .O(gate486inter3));
  inv1  gate2035(.a(s_213), .O(gate486inter4));
  nand2 gate2036(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2037(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2038(.a(G1234), .O(gate486inter7));
  inv1  gate2039(.a(G1235), .O(gate486inter8));
  nand2 gate2040(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2041(.a(s_213), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2042(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2043(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2044(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2549(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2550(.a(gate487inter0), .b(s_286), .O(gate487inter1));
  and2  gate2551(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2552(.a(s_286), .O(gate487inter3));
  inv1  gate2553(.a(s_287), .O(gate487inter4));
  nand2 gate2554(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2555(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2556(.a(G1236), .O(gate487inter7));
  inv1  gate2557(.a(G1237), .O(gate487inter8));
  nand2 gate2558(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2559(.a(s_287), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2560(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2561(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2562(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2647(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2648(.a(gate489inter0), .b(s_300), .O(gate489inter1));
  and2  gate2649(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2650(.a(s_300), .O(gate489inter3));
  inv1  gate2651(.a(s_301), .O(gate489inter4));
  nand2 gate2652(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2653(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2654(.a(G1240), .O(gate489inter7));
  inv1  gate2655(.a(G1241), .O(gate489inter8));
  nand2 gate2656(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2657(.a(s_301), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2658(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2659(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2660(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate2087(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2088(.a(gate490inter0), .b(s_220), .O(gate490inter1));
  and2  gate2089(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2090(.a(s_220), .O(gate490inter3));
  inv1  gate2091(.a(s_221), .O(gate490inter4));
  nand2 gate2092(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2093(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2094(.a(G1242), .O(gate490inter7));
  inv1  gate2095(.a(G1243), .O(gate490inter8));
  nand2 gate2096(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2097(.a(s_221), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2098(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2099(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2100(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1457(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1458(.a(gate492inter0), .b(s_130), .O(gate492inter1));
  and2  gate1459(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1460(.a(s_130), .O(gate492inter3));
  inv1  gate1461(.a(s_131), .O(gate492inter4));
  nand2 gate1462(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1463(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1464(.a(G1246), .O(gate492inter7));
  inv1  gate1465(.a(G1247), .O(gate492inter8));
  nand2 gate1466(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1467(.a(s_131), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1468(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1469(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1470(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2157(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2158(.a(gate493inter0), .b(s_230), .O(gate493inter1));
  and2  gate2159(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2160(.a(s_230), .O(gate493inter3));
  inv1  gate2161(.a(s_231), .O(gate493inter4));
  nand2 gate2162(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2163(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2164(.a(G1248), .O(gate493inter7));
  inv1  gate2165(.a(G1249), .O(gate493inter8));
  nand2 gate2166(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2167(.a(s_231), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2168(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2169(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2170(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1205(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1206(.a(gate496inter0), .b(s_94), .O(gate496inter1));
  and2  gate1207(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1208(.a(s_94), .O(gate496inter3));
  inv1  gate1209(.a(s_95), .O(gate496inter4));
  nand2 gate1210(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1211(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1212(.a(G1254), .O(gate496inter7));
  inv1  gate1213(.a(G1255), .O(gate496inter8));
  nand2 gate1214(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1215(.a(s_95), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1216(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1217(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1218(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1737(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1738(.a(gate497inter0), .b(s_170), .O(gate497inter1));
  and2  gate1739(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1740(.a(s_170), .O(gate497inter3));
  inv1  gate1741(.a(s_171), .O(gate497inter4));
  nand2 gate1742(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1743(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1744(.a(G1256), .O(gate497inter7));
  inv1  gate1745(.a(G1257), .O(gate497inter8));
  nand2 gate1746(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1747(.a(s_171), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1748(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1749(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1750(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2297(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2298(.a(gate503inter0), .b(s_250), .O(gate503inter1));
  and2  gate2299(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2300(.a(s_250), .O(gate503inter3));
  inv1  gate2301(.a(s_251), .O(gate503inter4));
  nand2 gate2302(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2303(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2304(.a(G1268), .O(gate503inter7));
  inv1  gate2305(.a(G1269), .O(gate503inter8));
  nand2 gate2306(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2307(.a(s_251), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2308(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2309(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2310(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1233(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1234(.a(gate506inter0), .b(s_98), .O(gate506inter1));
  and2  gate1235(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1236(.a(s_98), .O(gate506inter3));
  inv1  gate1237(.a(s_99), .O(gate506inter4));
  nand2 gate1238(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1239(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1240(.a(G1274), .O(gate506inter7));
  inv1  gate1241(.a(G1275), .O(gate506inter8));
  nand2 gate1242(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1243(.a(s_99), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1244(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1245(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1246(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1443(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1444(.a(gate508inter0), .b(s_128), .O(gate508inter1));
  and2  gate1445(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1446(.a(s_128), .O(gate508inter3));
  inv1  gate1447(.a(s_129), .O(gate508inter4));
  nand2 gate1448(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1449(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1450(.a(G1278), .O(gate508inter7));
  inv1  gate1451(.a(G1279), .O(gate508inter8));
  nand2 gate1452(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1453(.a(s_129), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1454(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1455(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1456(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule