module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate603(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate604(.a(gate9inter0), .b(s_8), .O(gate9inter1));
  and2  gate605(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate606(.a(s_8), .O(gate9inter3));
  inv1  gate607(.a(s_9), .O(gate9inter4));
  nand2 gate608(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate609(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate610(.a(G1), .O(gate9inter7));
  inv1  gate611(.a(G2), .O(gate9inter8));
  nand2 gate612(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate613(.a(s_9), .b(gate9inter3), .O(gate9inter10));
  nor2  gate614(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate615(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate616(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2017(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2018(.a(gate11inter0), .b(s_210), .O(gate11inter1));
  and2  gate2019(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2020(.a(s_210), .O(gate11inter3));
  inv1  gate2021(.a(s_211), .O(gate11inter4));
  nand2 gate2022(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2023(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2024(.a(G5), .O(gate11inter7));
  inv1  gate2025(.a(G6), .O(gate11inter8));
  nand2 gate2026(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2027(.a(s_211), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2028(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2029(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2030(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate771(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate772(.a(gate13inter0), .b(s_32), .O(gate13inter1));
  and2  gate773(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate774(.a(s_32), .O(gate13inter3));
  inv1  gate775(.a(s_33), .O(gate13inter4));
  nand2 gate776(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate777(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate778(.a(G9), .O(gate13inter7));
  inv1  gate779(.a(G10), .O(gate13inter8));
  nand2 gate780(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate781(.a(s_33), .b(gate13inter3), .O(gate13inter10));
  nor2  gate782(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate783(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate784(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1821(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1822(.a(gate14inter0), .b(s_182), .O(gate14inter1));
  and2  gate1823(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1824(.a(s_182), .O(gate14inter3));
  inv1  gate1825(.a(s_183), .O(gate14inter4));
  nand2 gate1826(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1827(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1828(.a(G11), .O(gate14inter7));
  inv1  gate1829(.a(G12), .O(gate14inter8));
  nand2 gate1830(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1831(.a(s_183), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1832(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1833(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1834(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate3095(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate3096(.a(gate15inter0), .b(s_364), .O(gate15inter1));
  and2  gate3097(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate3098(.a(s_364), .O(gate15inter3));
  inv1  gate3099(.a(s_365), .O(gate15inter4));
  nand2 gate3100(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate3101(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate3102(.a(G13), .O(gate15inter7));
  inv1  gate3103(.a(G14), .O(gate15inter8));
  nand2 gate3104(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate3105(.a(s_365), .b(gate15inter3), .O(gate15inter10));
  nor2  gate3106(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate3107(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate3108(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1079(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1080(.a(gate16inter0), .b(s_76), .O(gate16inter1));
  and2  gate1081(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1082(.a(s_76), .O(gate16inter3));
  inv1  gate1083(.a(s_77), .O(gate16inter4));
  nand2 gate1084(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1085(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1086(.a(G15), .O(gate16inter7));
  inv1  gate1087(.a(G16), .O(gate16inter8));
  nand2 gate1088(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1089(.a(s_77), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1090(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1091(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1092(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2703(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2704(.a(gate18inter0), .b(s_308), .O(gate18inter1));
  and2  gate2705(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2706(.a(s_308), .O(gate18inter3));
  inv1  gate2707(.a(s_309), .O(gate18inter4));
  nand2 gate2708(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2709(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2710(.a(G19), .O(gate18inter7));
  inv1  gate2711(.a(G20), .O(gate18inter8));
  nand2 gate2712(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2713(.a(s_309), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2714(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2715(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2716(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1695(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1696(.a(gate19inter0), .b(s_164), .O(gate19inter1));
  and2  gate1697(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1698(.a(s_164), .O(gate19inter3));
  inv1  gate1699(.a(s_165), .O(gate19inter4));
  nand2 gate1700(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1701(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1702(.a(G21), .O(gate19inter7));
  inv1  gate1703(.a(G22), .O(gate19inter8));
  nand2 gate1704(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1705(.a(s_165), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1706(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1707(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1708(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate855(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate856(.a(gate20inter0), .b(s_44), .O(gate20inter1));
  and2  gate857(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate858(.a(s_44), .O(gate20inter3));
  inv1  gate859(.a(s_45), .O(gate20inter4));
  nand2 gate860(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate861(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate862(.a(G23), .O(gate20inter7));
  inv1  gate863(.a(G24), .O(gate20inter8));
  nand2 gate864(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate865(.a(s_45), .b(gate20inter3), .O(gate20inter10));
  nor2  gate866(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate867(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate868(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1261(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1262(.a(gate22inter0), .b(s_102), .O(gate22inter1));
  and2  gate1263(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1264(.a(s_102), .O(gate22inter3));
  inv1  gate1265(.a(s_103), .O(gate22inter4));
  nand2 gate1266(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1267(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1268(.a(G27), .O(gate22inter7));
  inv1  gate1269(.a(G28), .O(gate22inter8));
  nand2 gate1270(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1271(.a(s_103), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1272(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1273(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1274(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2857(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2858(.a(gate23inter0), .b(s_330), .O(gate23inter1));
  and2  gate2859(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2860(.a(s_330), .O(gate23inter3));
  inv1  gate2861(.a(s_331), .O(gate23inter4));
  nand2 gate2862(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2863(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2864(.a(G29), .O(gate23inter7));
  inv1  gate2865(.a(G30), .O(gate23inter8));
  nand2 gate2866(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2867(.a(s_331), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2868(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2869(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2870(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1219(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1220(.a(gate29inter0), .b(s_96), .O(gate29inter1));
  and2  gate1221(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1222(.a(s_96), .O(gate29inter3));
  inv1  gate1223(.a(s_97), .O(gate29inter4));
  nand2 gate1224(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1225(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1226(.a(G3), .O(gate29inter7));
  inv1  gate1227(.a(G7), .O(gate29inter8));
  nand2 gate1228(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1229(.a(s_97), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1230(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1231(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1232(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate3067(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate3068(.a(gate31inter0), .b(s_360), .O(gate31inter1));
  and2  gate3069(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate3070(.a(s_360), .O(gate31inter3));
  inv1  gate3071(.a(s_361), .O(gate31inter4));
  nand2 gate3072(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate3073(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate3074(.a(G4), .O(gate31inter7));
  inv1  gate3075(.a(G8), .O(gate31inter8));
  nand2 gate3076(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate3077(.a(s_361), .b(gate31inter3), .O(gate31inter10));
  nor2  gate3078(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate3079(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate3080(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate2409(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2410(.a(gate32inter0), .b(s_266), .O(gate32inter1));
  and2  gate2411(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2412(.a(s_266), .O(gate32inter3));
  inv1  gate2413(.a(s_267), .O(gate32inter4));
  nand2 gate2414(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2415(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2416(.a(G12), .O(gate32inter7));
  inv1  gate2417(.a(G16), .O(gate32inter8));
  nand2 gate2418(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2419(.a(s_267), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2420(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2421(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2422(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1233(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1234(.a(gate36inter0), .b(s_98), .O(gate36inter1));
  and2  gate1235(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1236(.a(s_98), .O(gate36inter3));
  inv1  gate1237(.a(s_99), .O(gate36inter4));
  nand2 gate1238(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1239(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1240(.a(G26), .O(gate36inter7));
  inv1  gate1241(.a(G30), .O(gate36inter8));
  nand2 gate1242(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1243(.a(s_99), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1244(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1245(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1246(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate2185(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2186(.a(gate37inter0), .b(s_234), .O(gate37inter1));
  and2  gate2187(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2188(.a(s_234), .O(gate37inter3));
  inv1  gate2189(.a(s_235), .O(gate37inter4));
  nand2 gate2190(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2191(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2192(.a(G19), .O(gate37inter7));
  inv1  gate2193(.a(G23), .O(gate37inter8));
  nand2 gate2194(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2195(.a(s_235), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2196(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2197(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2198(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1443(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1444(.a(gate39inter0), .b(s_128), .O(gate39inter1));
  and2  gate1445(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1446(.a(s_128), .O(gate39inter3));
  inv1  gate1447(.a(s_129), .O(gate39inter4));
  nand2 gate1448(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1449(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1450(.a(G20), .O(gate39inter7));
  inv1  gate1451(.a(G24), .O(gate39inter8));
  nand2 gate1452(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1453(.a(s_129), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1454(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1455(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1456(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate631(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate632(.a(gate40inter0), .b(s_12), .O(gate40inter1));
  and2  gate633(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate634(.a(s_12), .O(gate40inter3));
  inv1  gate635(.a(s_13), .O(gate40inter4));
  nand2 gate636(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate637(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate638(.a(G28), .O(gate40inter7));
  inv1  gate639(.a(G32), .O(gate40inter8));
  nand2 gate640(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate641(.a(s_13), .b(gate40inter3), .O(gate40inter10));
  nor2  gate642(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate643(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate644(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate547(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate548(.a(gate41inter0), .b(s_0), .O(gate41inter1));
  and2  gate549(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate550(.a(s_0), .O(gate41inter3));
  inv1  gate551(.a(s_1), .O(gate41inter4));
  nand2 gate552(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate553(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate554(.a(G1), .O(gate41inter7));
  inv1  gate555(.a(G266), .O(gate41inter8));
  nand2 gate556(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate557(.a(s_1), .b(gate41inter3), .O(gate41inter10));
  nor2  gate558(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate559(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate560(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1317(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1318(.a(gate43inter0), .b(s_110), .O(gate43inter1));
  and2  gate1319(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1320(.a(s_110), .O(gate43inter3));
  inv1  gate1321(.a(s_111), .O(gate43inter4));
  nand2 gate1322(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1323(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1324(.a(G3), .O(gate43inter7));
  inv1  gate1325(.a(G269), .O(gate43inter8));
  nand2 gate1326(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1327(.a(s_111), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1328(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1329(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1330(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2633(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2634(.a(gate44inter0), .b(s_298), .O(gate44inter1));
  and2  gate2635(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2636(.a(s_298), .O(gate44inter3));
  inv1  gate2637(.a(s_299), .O(gate44inter4));
  nand2 gate2638(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2639(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2640(.a(G4), .O(gate44inter7));
  inv1  gate2641(.a(G269), .O(gate44inter8));
  nand2 gate2642(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2643(.a(s_299), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2644(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2645(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2646(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2787(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2788(.a(gate46inter0), .b(s_320), .O(gate46inter1));
  and2  gate2789(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2790(.a(s_320), .O(gate46inter3));
  inv1  gate2791(.a(s_321), .O(gate46inter4));
  nand2 gate2792(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2793(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2794(.a(G6), .O(gate46inter7));
  inv1  gate2795(.a(G272), .O(gate46inter8));
  nand2 gate2796(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2797(.a(s_321), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2798(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2799(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2800(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1933(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1934(.a(gate47inter0), .b(s_198), .O(gate47inter1));
  and2  gate1935(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1936(.a(s_198), .O(gate47inter3));
  inv1  gate1937(.a(s_199), .O(gate47inter4));
  nand2 gate1938(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1939(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1940(.a(G7), .O(gate47inter7));
  inv1  gate1941(.a(G275), .O(gate47inter8));
  nand2 gate1942(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1943(.a(s_199), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1944(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1945(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1946(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2003(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2004(.a(gate48inter0), .b(s_208), .O(gate48inter1));
  and2  gate2005(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2006(.a(s_208), .O(gate48inter3));
  inv1  gate2007(.a(s_209), .O(gate48inter4));
  nand2 gate2008(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2009(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2010(.a(G8), .O(gate48inter7));
  inv1  gate2011(.a(G275), .O(gate48inter8));
  nand2 gate2012(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2013(.a(s_209), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2014(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2015(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2016(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1359(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1360(.a(gate51inter0), .b(s_116), .O(gate51inter1));
  and2  gate1361(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1362(.a(s_116), .O(gate51inter3));
  inv1  gate1363(.a(s_117), .O(gate51inter4));
  nand2 gate1364(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1365(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1366(.a(G11), .O(gate51inter7));
  inv1  gate1367(.a(G281), .O(gate51inter8));
  nand2 gate1368(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1369(.a(s_117), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1370(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1371(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1372(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1121(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1122(.a(gate52inter0), .b(s_82), .O(gate52inter1));
  and2  gate1123(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1124(.a(s_82), .O(gate52inter3));
  inv1  gate1125(.a(s_83), .O(gate52inter4));
  nand2 gate1126(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1127(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1128(.a(G12), .O(gate52inter7));
  inv1  gate1129(.a(G281), .O(gate52inter8));
  nand2 gate1130(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1131(.a(s_83), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1132(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1133(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1134(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1611(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1612(.a(gate53inter0), .b(s_152), .O(gate53inter1));
  and2  gate1613(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1614(.a(s_152), .O(gate53inter3));
  inv1  gate1615(.a(s_153), .O(gate53inter4));
  nand2 gate1616(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1617(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1618(.a(G13), .O(gate53inter7));
  inv1  gate1619(.a(G284), .O(gate53inter8));
  nand2 gate1620(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1621(.a(s_153), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1622(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1623(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1624(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1275(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1276(.a(gate55inter0), .b(s_104), .O(gate55inter1));
  and2  gate1277(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1278(.a(s_104), .O(gate55inter3));
  inv1  gate1279(.a(s_105), .O(gate55inter4));
  nand2 gate1280(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1281(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1282(.a(G15), .O(gate55inter7));
  inv1  gate1283(.a(G287), .O(gate55inter8));
  nand2 gate1284(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1285(.a(s_105), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1286(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1287(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1288(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2157(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2158(.a(gate56inter0), .b(s_230), .O(gate56inter1));
  and2  gate2159(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2160(.a(s_230), .O(gate56inter3));
  inv1  gate2161(.a(s_231), .O(gate56inter4));
  nand2 gate2162(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2163(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2164(.a(G16), .O(gate56inter7));
  inv1  gate2165(.a(G287), .O(gate56inter8));
  nand2 gate2166(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2167(.a(s_231), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2168(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2169(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2170(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2941(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2942(.a(gate59inter0), .b(s_342), .O(gate59inter1));
  and2  gate2943(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2944(.a(s_342), .O(gate59inter3));
  inv1  gate2945(.a(s_343), .O(gate59inter4));
  nand2 gate2946(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2947(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2948(.a(G19), .O(gate59inter7));
  inv1  gate2949(.a(G293), .O(gate59inter8));
  nand2 gate2950(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2951(.a(s_343), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2952(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2953(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2954(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1681(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1682(.a(gate62inter0), .b(s_162), .O(gate62inter1));
  and2  gate1683(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1684(.a(s_162), .O(gate62inter3));
  inv1  gate1685(.a(s_163), .O(gate62inter4));
  nand2 gate1686(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1687(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1688(.a(G22), .O(gate62inter7));
  inv1  gate1689(.a(G296), .O(gate62inter8));
  nand2 gate1690(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1691(.a(s_163), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1692(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1693(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1694(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1541(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1542(.a(gate63inter0), .b(s_142), .O(gate63inter1));
  and2  gate1543(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1544(.a(s_142), .O(gate63inter3));
  inv1  gate1545(.a(s_143), .O(gate63inter4));
  nand2 gate1546(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1547(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1548(.a(G23), .O(gate63inter7));
  inv1  gate1549(.a(G299), .O(gate63inter8));
  nand2 gate1550(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1551(.a(s_143), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1552(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1553(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1554(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2437(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2438(.a(gate66inter0), .b(s_270), .O(gate66inter1));
  and2  gate2439(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2440(.a(s_270), .O(gate66inter3));
  inv1  gate2441(.a(s_271), .O(gate66inter4));
  nand2 gate2442(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2443(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2444(.a(G26), .O(gate66inter7));
  inv1  gate2445(.a(G302), .O(gate66inter8));
  nand2 gate2446(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2447(.a(s_271), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2448(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2449(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2450(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate827(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate828(.a(gate67inter0), .b(s_40), .O(gate67inter1));
  and2  gate829(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate830(.a(s_40), .O(gate67inter3));
  inv1  gate831(.a(s_41), .O(gate67inter4));
  nand2 gate832(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate833(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate834(.a(G27), .O(gate67inter7));
  inv1  gate835(.a(G305), .O(gate67inter8));
  nand2 gate836(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate837(.a(s_41), .b(gate67inter3), .O(gate67inter10));
  nor2  gate838(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate839(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate840(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2395(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2396(.a(gate69inter0), .b(s_264), .O(gate69inter1));
  and2  gate2397(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2398(.a(s_264), .O(gate69inter3));
  inv1  gate2399(.a(s_265), .O(gate69inter4));
  nand2 gate2400(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2401(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2402(.a(G29), .O(gate69inter7));
  inv1  gate2403(.a(G308), .O(gate69inter8));
  nand2 gate2404(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2405(.a(s_265), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2406(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2407(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2408(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate617(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate618(.a(gate73inter0), .b(s_10), .O(gate73inter1));
  and2  gate619(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate620(.a(s_10), .O(gate73inter3));
  inv1  gate621(.a(s_11), .O(gate73inter4));
  nand2 gate622(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate623(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate624(.a(G1), .O(gate73inter7));
  inv1  gate625(.a(G314), .O(gate73inter8));
  nand2 gate626(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate627(.a(s_11), .b(gate73inter3), .O(gate73inter10));
  nor2  gate628(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate629(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate630(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2479(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2480(.a(gate77inter0), .b(s_276), .O(gate77inter1));
  and2  gate2481(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2482(.a(s_276), .O(gate77inter3));
  inv1  gate2483(.a(s_277), .O(gate77inter4));
  nand2 gate2484(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2485(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2486(.a(G2), .O(gate77inter7));
  inv1  gate2487(.a(G320), .O(gate77inter8));
  nand2 gate2488(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2489(.a(s_277), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2490(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2491(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2492(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate2115(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2116(.a(gate78inter0), .b(s_224), .O(gate78inter1));
  and2  gate2117(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2118(.a(s_224), .O(gate78inter3));
  inv1  gate2119(.a(s_225), .O(gate78inter4));
  nand2 gate2120(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2121(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2122(.a(G6), .O(gate78inter7));
  inv1  gate2123(.a(G320), .O(gate78inter8));
  nand2 gate2124(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2125(.a(s_225), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2126(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2127(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2128(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2885(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2886(.a(gate80inter0), .b(s_334), .O(gate80inter1));
  and2  gate2887(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2888(.a(s_334), .O(gate80inter3));
  inv1  gate2889(.a(s_335), .O(gate80inter4));
  nand2 gate2890(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2891(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2892(.a(G14), .O(gate80inter7));
  inv1  gate2893(.a(G323), .O(gate80inter8));
  nand2 gate2894(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2895(.a(s_335), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2896(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2897(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2898(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1247(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1248(.a(gate82inter0), .b(s_100), .O(gate82inter1));
  and2  gate1249(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1250(.a(s_100), .O(gate82inter3));
  inv1  gate1251(.a(s_101), .O(gate82inter4));
  nand2 gate1252(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1253(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1254(.a(G7), .O(gate82inter7));
  inv1  gate1255(.a(G326), .O(gate82inter8));
  nand2 gate1256(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1257(.a(s_101), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1258(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1259(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1260(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1555(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1556(.a(gate84inter0), .b(s_144), .O(gate84inter1));
  and2  gate1557(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1558(.a(s_144), .O(gate84inter3));
  inv1  gate1559(.a(s_145), .O(gate84inter4));
  nand2 gate1560(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1561(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1562(.a(G15), .O(gate84inter7));
  inv1  gate1563(.a(G329), .O(gate84inter8));
  nand2 gate1564(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1565(.a(s_145), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1566(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1567(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1568(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate3137(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate3138(.a(gate85inter0), .b(s_370), .O(gate85inter1));
  and2  gate3139(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate3140(.a(s_370), .O(gate85inter3));
  inv1  gate3141(.a(s_371), .O(gate85inter4));
  nand2 gate3142(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate3143(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate3144(.a(G4), .O(gate85inter7));
  inv1  gate3145(.a(G332), .O(gate85inter8));
  nand2 gate3146(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate3147(.a(s_371), .b(gate85inter3), .O(gate85inter10));
  nor2  gate3148(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate3149(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate3150(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1429(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1430(.a(gate86inter0), .b(s_126), .O(gate86inter1));
  and2  gate1431(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1432(.a(s_126), .O(gate86inter3));
  inv1  gate1433(.a(s_127), .O(gate86inter4));
  nand2 gate1434(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1435(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1436(.a(G8), .O(gate86inter7));
  inv1  gate1437(.a(G332), .O(gate86inter8));
  nand2 gate1438(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1439(.a(s_127), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1440(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1441(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1442(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2717(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2718(.a(gate88inter0), .b(s_310), .O(gate88inter1));
  and2  gate2719(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2720(.a(s_310), .O(gate88inter3));
  inv1  gate2721(.a(s_311), .O(gate88inter4));
  nand2 gate2722(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2723(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2724(.a(G16), .O(gate88inter7));
  inv1  gate2725(.a(G335), .O(gate88inter8));
  nand2 gate2726(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2727(.a(s_311), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2728(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2729(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2730(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1751(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1752(.a(gate89inter0), .b(s_172), .O(gate89inter1));
  and2  gate1753(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1754(.a(s_172), .O(gate89inter3));
  inv1  gate1755(.a(s_173), .O(gate89inter4));
  nand2 gate1756(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1757(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1758(.a(G17), .O(gate89inter7));
  inv1  gate1759(.a(G338), .O(gate89inter8));
  nand2 gate1760(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1761(.a(s_173), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1762(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1763(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1764(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2997(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2998(.a(gate92inter0), .b(s_350), .O(gate92inter1));
  and2  gate2999(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate3000(.a(s_350), .O(gate92inter3));
  inv1  gate3001(.a(s_351), .O(gate92inter4));
  nand2 gate3002(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate3003(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate3004(.a(G29), .O(gate92inter7));
  inv1  gate3005(.a(G341), .O(gate92inter8));
  nand2 gate3006(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate3007(.a(s_351), .b(gate92inter3), .O(gate92inter10));
  nor2  gate3008(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate3009(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate3010(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate2899(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2900(.a(gate93inter0), .b(s_336), .O(gate93inter1));
  and2  gate2901(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2902(.a(s_336), .O(gate93inter3));
  inv1  gate2903(.a(s_337), .O(gate93inter4));
  nand2 gate2904(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2905(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2906(.a(G18), .O(gate93inter7));
  inv1  gate2907(.a(G344), .O(gate93inter8));
  nand2 gate2908(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2909(.a(s_337), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2910(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2911(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2912(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1051(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1052(.a(gate95inter0), .b(s_72), .O(gate95inter1));
  and2  gate1053(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1054(.a(s_72), .O(gate95inter3));
  inv1  gate1055(.a(s_73), .O(gate95inter4));
  nand2 gate1056(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1057(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1058(.a(G26), .O(gate95inter7));
  inv1  gate1059(.a(G347), .O(gate95inter8));
  nand2 gate1060(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1061(.a(s_73), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1062(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1063(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1064(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate561(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate562(.a(gate96inter0), .b(s_2), .O(gate96inter1));
  and2  gate563(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate564(.a(s_2), .O(gate96inter3));
  inv1  gate565(.a(s_3), .O(gate96inter4));
  nand2 gate566(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate567(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate568(.a(G30), .O(gate96inter7));
  inv1  gate569(.a(G347), .O(gate96inter8));
  nand2 gate570(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate571(.a(s_3), .b(gate96inter3), .O(gate96inter10));
  nor2  gate572(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate573(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate574(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2577(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2578(.a(gate100inter0), .b(s_290), .O(gate100inter1));
  and2  gate2579(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2580(.a(s_290), .O(gate100inter3));
  inv1  gate2581(.a(s_291), .O(gate100inter4));
  nand2 gate2582(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2583(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2584(.a(G31), .O(gate100inter7));
  inv1  gate2585(.a(G353), .O(gate100inter8));
  nand2 gate2586(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2587(.a(s_291), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2588(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2589(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2590(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate673(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate674(.a(gate101inter0), .b(s_18), .O(gate101inter1));
  and2  gate675(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate676(.a(s_18), .O(gate101inter3));
  inv1  gate677(.a(s_19), .O(gate101inter4));
  nand2 gate678(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate679(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate680(.a(G20), .O(gate101inter7));
  inv1  gate681(.a(G356), .O(gate101inter8));
  nand2 gate682(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate683(.a(s_19), .b(gate101inter3), .O(gate101inter10));
  nor2  gate684(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate685(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate686(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2815(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2816(.a(gate105inter0), .b(s_324), .O(gate105inter1));
  and2  gate2817(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2818(.a(s_324), .O(gate105inter3));
  inv1  gate2819(.a(s_325), .O(gate105inter4));
  nand2 gate2820(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2821(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2822(.a(G362), .O(gate105inter7));
  inv1  gate2823(.a(G363), .O(gate105inter8));
  nand2 gate2824(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2825(.a(s_325), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2826(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2827(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2828(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1387(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1388(.a(gate106inter0), .b(s_120), .O(gate106inter1));
  and2  gate1389(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1390(.a(s_120), .O(gate106inter3));
  inv1  gate1391(.a(s_121), .O(gate106inter4));
  nand2 gate1392(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1393(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1394(.a(G364), .O(gate106inter7));
  inv1  gate1395(.a(G365), .O(gate106inter8));
  nand2 gate1396(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1397(.a(s_121), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1398(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1399(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1400(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1737(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1738(.a(gate108inter0), .b(s_170), .O(gate108inter1));
  and2  gate1739(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1740(.a(s_170), .O(gate108inter3));
  inv1  gate1741(.a(s_171), .O(gate108inter4));
  nand2 gate1742(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1743(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1744(.a(G368), .O(gate108inter7));
  inv1  gate1745(.a(G369), .O(gate108inter8));
  nand2 gate1746(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1747(.a(s_171), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1748(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1749(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1750(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate2269(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2270(.a(gate109inter0), .b(s_246), .O(gate109inter1));
  and2  gate2271(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2272(.a(s_246), .O(gate109inter3));
  inv1  gate2273(.a(s_247), .O(gate109inter4));
  nand2 gate2274(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2275(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2276(.a(G370), .O(gate109inter7));
  inv1  gate2277(.a(G371), .O(gate109inter8));
  nand2 gate2278(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2279(.a(s_247), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2280(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2281(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2282(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1975(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1976(.a(gate112inter0), .b(s_204), .O(gate112inter1));
  and2  gate1977(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1978(.a(s_204), .O(gate112inter3));
  inv1  gate1979(.a(s_205), .O(gate112inter4));
  nand2 gate1980(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1981(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1982(.a(G376), .O(gate112inter7));
  inv1  gate1983(.a(G377), .O(gate112inter8));
  nand2 gate1984(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1985(.a(s_205), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1986(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1987(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1988(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate967(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate968(.a(gate113inter0), .b(s_60), .O(gate113inter1));
  and2  gate969(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate970(.a(s_60), .O(gate113inter3));
  inv1  gate971(.a(s_61), .O(gate113inter4));
  nand2 gate972(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate973(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate974(.a(G378), .O(gate113inter7));
  inv1  gate975(.a(G379), .O(gate113inter8));
  nand2 gate976(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate977(.a(s_61), .b(gate113inter3), .O(gate113inter10));
  nor2  gate978(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate979(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate980(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1625(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1626(.a(gate118inter0), .b(s_154), .O(gate118inter1));
  and2  gate1627(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1628(.a(s_154), .O(gate118inter3));
  inv1  gate1629(.a(s_155), .O(gate118inter4));
  nand2 gate1630(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1631(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1632(.a(G388), .O(gate118inter7));
  inv1  gate1633(.a(G389), .O(gate118inter8));
  nand2 gate1634(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1635(.a(s_155), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1636(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1637(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1638(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2283(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2284(.a(gate119inter0), .b(s_248), .O(gate119inter1));
  and2  gate2285(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2286(.a(s_248), .O(gate119inter3));
  inv1  gate2287(.a(s_249), .O(gate119inter4));
  nand2 gate2288(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2289(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2290(.a(G390), .O(gate119inter7));
  inv1  gate2291(.a(G391), .O(gate119inter8));
  nand2 gate2292(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2293(.a(s_249), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2294(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2295(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2296(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate813(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate814(.a(gate121inter0), .b(s_38), .O(gate121inter1));
  and2  gate815(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate816(.a(s_38), .O(gate121inter3));
  inv1  gate817(.a(s_39), .O(gate121inter4));
  nand2 gate818(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate819(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate820(.a(G394), .O(gate121inter7));
  inv1  gate821(.a(G395), .O(gate121inter8));
  nand2 gate822(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate823(.a(s_39), .b(gate121inter3), .O(gate121inter10));
  nor2  gate824(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate825(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate826(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2171(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2172(.a(gate122inter0), .b(s_232), .O(gate122inter1));
  and2  gate2173(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2174(.a(s_232), .O(gate122inter3));
  inv1  gate2175(.a(s_233), .O(gate122inter4));
  nand2 gate2176(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2177(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2178(.a(G396), .O(gate122inter7));
  inv1  gate2179(.a(G397), .O(gate122inter8));
  nand2 gate2180(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2181(.a(s_233), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2182(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2183(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2184(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate2227(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2228(.a(gate123inter0), .b(s_240), .O(gate123inter1));
  and2  gate2229(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2230(.a(s_240), .O(gate123inter3));
  inv1  gate2231(.a(s_241), .O(gate123inter4));
  nand2 gate2232(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2233(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2234(.a(G398), .O(gate123inter7));
  inv1  gate2235(.a(G399), .O(gate123inter8));
  nand2 gate2236(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2237(.a(s_241), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2238(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2239(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2240(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate687(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate688(.a(gate124inter0), .b(s_20), .O(gate124inter1));
  and2  gate689(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate690(.a(s_20), .O(gate124inter3));
  inv1  gate691(.a(s_21), .O(gate124inter4));
  nand2 gate692(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate693(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate694(.a(G400), .O(gate124inter7));
  inv1  gate695(.a(G401), .O(gate124inter8));
  nand2 gate696(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate697(.a(s_21), .b(gate124inter3), .O(gate124inter10));
  nor2  gate698(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate699(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate700(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate785(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate786(.a(gate125inter0), .b(s_34), .O(gate125inter1));
  and2  gate787(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate788(.a(s_34), .O(gate125inter3));
  inv1  gate789(.a(s_35), .O(gate125inter4));
  nand2 gate790(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate791(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate792(.a(G402), .O(gate125inter7));
  inv1  gate793(.a(G403), .O(gate125inter8));
  nand2 gate794(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate795(.a(s_35), .b(gate125inter3), .O(gate125inter10));
  nor2  gate796(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate797(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate798(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2129(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2130(.a(gate131inter0), .b(s_226), .O(gate131inter1));
  and2  gate2131(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2132(.a(s_226), .O(gate131inter3));
  inv1  gate2133(.a(s_227), .O(gate131inter4));
  nand2 gate2134(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2135(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2136(.a(G414), .O(gate131inter7));
  inv1  gate2137(.a(G415), .O(gate131inter8));
  nand2 gate2138(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2139(.a(s_227), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2140(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2141(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2142(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1205(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1206(.a(gate132inter0), .b(s_94), .O(gate132inter1));
  and2  gate1207(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1208(.a(s_94), .O(gate132inter3));
  inv1  gate1209(.a(s_95), .O(gate132inter4));
  nand2 gate1210(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1211(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1212(.a(G416), .O(gate132inter7));
  inv1  gate1213(.a(G417), .O(gate132inter8));
  nand2 gate1214(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1215(.a(s_95), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1216(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1217(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1218(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate729(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate730(.a(gate142inter0), .b(s_26), .O(gate142inter1));
  and2  gate731(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate732(.a(s_26), .O(gate142inter3));
  inv1  gate733(.a(s_27), .O(gate142inter4));
  nand2 gate734(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate735(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate736(.a(G456), .O(gate142inter7));
  inv1  gate737(.a(G459), .O(gate142inter8));
  nand2 gate738(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate739(.a(s_27), .b(gate142inter3), .O(gate142inter10));
  nor2  gate740(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate741(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate742(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate3025(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate3026(.a(gate143inter0), .b(s_354), .O(gate143inter1));
  and2  gate3027(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate3028(.a(s_354), .O(gate143inter3));
  inv1  gate3029(.a(s_355), .O(gate143inter4));
  nand2 gate3030(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate3031(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate3032(.a(G462), .O(gate143inter7));
  inv1  gate3033(.a(G465), .O(gate143inter8));
  nand2 gate3034(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate3035(.a(s_355), .b(gate143inter3), .O(gate143inter10));
  nor2  gate3036(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate3037(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate3038(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1163(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1164(.a(gate144inter0), .b(s_88), .O(gate144inter1));
  and2  gate1165(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1166(.a(s_88), .O(gate144inter3));
  inv1  gate1167(.a(s_89), .O(gate144inter4));
  nand2 gate1168(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1169(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1170(.a(G468), .O(gate144inter7));
  inv1  gate1171(.a(G471), .O(gate144inter8));
  nand2 gate1172(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1173(.a(s_89), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1174(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1175(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1176(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate3109(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate3110(.a(gate145inter0), .b(s_366), .O(gate145inter1));
  and2  gate3111(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate3112(.a(s_366), .O(gate145inter3));
  inv1  gate3113(.a(s_367), .O(gate145inter4));
  nand2 gate3114(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate3115(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate3116(.a(G474), .O(gate145inter7));
  inv1  gate3117(.a(G477), .O(gate145inter8));
  nand2 gate3118(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate3119(.a(s_367), .b(gate145inter3), .O(gate145inter10));
  nor2  gate3120(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate3121(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate3122(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1891(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1892(.a(gate148inter0), .b(s_192), .O(gate148inter1));
  and2  gate1893(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1894(.a(s_192), .O(gate148inter3));
  inv1  gate1895(.a(s_193), .O(gate148inter4));
  nand2 gate1896(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1897(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1898(.a(G492), .O(gate148inter7));
  inv1  gate1899(.a(G495), .O(gate148inter8));
  nand2 gate1900(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1901(.a(s_193), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1902(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1903(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1904(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate3081(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate3082(.a(gate149inter0), .b(s_362), .O(gate149inter1));
  and2  gate3083(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate3084(.a(s_362), .O(gate149inter3));
  inv1  gate3085(.a(s_363), .O(gate149inter4));
  nand2 gate3086(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate3087(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate3088(.a(G498), .O(gate149inter7));
  inv1  gate3089(.a(G501), .O(gate149inter8));
  nand2 gate3090(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate3091(.a(s_363), .b(gate149inter3), .O(gate149inter10));
  nor2  gate3092(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate3093(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate3094(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1345(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1346(.a(gate152inter0), .b(s_114), .O(gate152inter1));
  and2  gate1347(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1348(.a(s_114), .O(gate152inter3));
  inv1  gate1349(.a(s_115), .O(gate152inter4));
  nand2 gate1350(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1351(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1352(.a(G516), .O(gate152inter7));
  inv1  gate1353(.a(G519), .O(gate152inter8));
  nand2 gate1354(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1355(.a(s_115), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1356(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1357(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1358(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1961(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1962(.a(gate155inter0), .b(s_202), .O(gate155inter1));
  and2  gate1963(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1964(.a(s_202), .O(gate155inter3));
  inv1  gate1965(.a(s_203), .O(gate155inter4));
  nand2 gate1966(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1967(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1968(.a(G432), .O(gate155inter7));
  inv1  gate1969(.a(G525), .O(gate155inter8));
  nand2 gate1970(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1971(.a(s_203), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1972(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1973(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1974(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2199(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2200(.a(gate157inter0), .b(s_236), .O(gate157inter1));
  and2  gate2201(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2202(.a(s_236), .O(gate157inter3));
  inv1  gate2203(.a(s_237), .O(gate157inter4));
  nand2 gate2204(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2205(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2206(.a(G438), .O(gate157inter7));
  inv1  gate2207(.a(G528), .O(gate157inter8));
  nand2 gate2208(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2209(.a(s_237), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2210(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2211(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2212(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1513(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1514(.a(gate158inter0), .b(s_138), .O(gate158inter1));
  and2  gate1515(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1516(.a(s_138), .O(gate158inter3));
  inv1  gate1517(.a(s_139), .O(gate158inter4));
  nand2 gate1518(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1519(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1520(.a(G441), .O(gate158inter7));
  inv1  gate1521(.a(G528), .O(gate158inter8));
  nand2 gate1522(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1523(.a(s_139), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1524(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1525(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1526(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2087(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2088(.a(gate159inter0), .b(s_220), .O(gate159inter1));
  and2  gate2089(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2090(.a(s_220), .O(gate159inter3));
  inv1  gate2091(.a(s_221), .O(gate159inter4));
  nand2 gate2092(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2093(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2094(.a(G444), .O(gate159inter7));
  inv1  gate2095(.a(G531), .O(gate159inter8));
  nand2 gate2096(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2097(.a(s_221), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2098(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2099(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2100(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate757(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate758(.a(gate160inter0), .b(s_30), .O(gate160inter1));
  and2  gate759(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate760(.a(s_30), .O(gate160inter3));
  inv1  gate761(.a(s_31), .O(gate160inter4));
  nand2 gate762(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate763(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate764(.a(G447), .O(gate160inter7));
  inv1  gate765(.a(G531), .O(gate160inter8));
  nand2 gate766(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate767(.a(s_31), .b(gate160inter3), .O(gate160inter10));
  nor2  gate768(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate769(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate770(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate2255(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2256(.a(gate161inter0), .b(s_244), .O(gate161inter1));
  and2  gate2257(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2258(.a(s_244), .O(gate161inter3));
  inv1  gate2259(.a(s_245), .O(gate161inter4));
  nand2 gate2260(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2261(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2262(.a(G450), .O(gate161inter7));
  inv1  gate2263(.a(G534), .O(gate161inter8));
  nand2 gate2264(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2265(.a(s_245), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2266(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2267(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2268(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate645(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate646(.a(gate162inter0), .b(s_14), .O(gate162inter1));
  and2  gate647(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate648(.a(s_14), .O(gate162inter3));
  inv1  gate649(.a(s_15), .O(gate162inter4));
  nand2 gate650(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate651(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate652(.a(G453), .O(gate162inter7));
  inv1  gate653(.a(G534), .O(gate162inter8));
  nand2 gate654(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate655(.a(s_15), .b(gate162inter3), .O(gate162inter10));
  nor2  gate656(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate657(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate658(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate869(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate870(.a(gate164inter0), .b(s_46), .O(gate164inter1));
  and2  gate871(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate872(.a(s_46), .O(gate164inter3));
  inv1  gate873(.a(s_47), .O(gate164inter4));
  nand2 gate874(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate875(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate876(.a(G459), .O(gate164inter7));
  inv1  gate877(.a(G537), .O(gate164inter8));
  nand2 gate878(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate879(.a(s_47), .b(gate164inter3), .O(gate164inter10));
  nor2  gate880(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate881(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate882(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate2073(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2074(.a(gate165inter0), .b(s_218), .O(gate165inter1));
  and2  gate2075(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2076(.a(s_218), .O(gate165inter3));
  inv1  gate2077(.a(s_219), .O(gate165inter4));
  nand2 gate2078(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2079(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2080(.a(G462), .O(gate165inter7));
  inv1  gate2081(.a(G540), .O(gate165inter8));
  nand2 gate2082(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2083(.a(s_219), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2084(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2085(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2086(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2605(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2606(.a(gate167inter0), .b(s_294), .O(gate167inter1));
  and2  gate2607(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2608(.a(s_294), .O(gate167inter3));
  inv1  gate2609(.a(s_295), .O(gate167inter4));
  nand2 gate2610(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2611(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2612(.a(G468), .O(gate167inter7));
  inv1  gate2613(.a(G543), .O(gate167inter8));
  nand2 gate2614(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2615(.a(s_295), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2616(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2617(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2618(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2521(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2522(.a(gate169inter0), .b(s_282), .O(gate169inter1));
  and2  gate2523(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2524(.a(s_282), .O(gate169inter3));
  inv1  gate2525(.a(s_283), .O(gate169inter4));
  nand2 gate2526(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2527(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2528(.a(G474), .O(gate169inter7));
  inv1  gate2529(.a(G546), .O(gate169inter8));
  nand2 gate2530(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2531(.a(s_283), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2532(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2533(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2534(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate715(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate716(.a(gate171inter0), .b(s_24), .O(gate171inter1));
  and2  gate717(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate718(.a(s_24), .O(gate171inter3));
  inv1  gate719(.a(s_25), .O(gate171inter4));
  nand2 gate720(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate721(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate722(.a(G480), .O(gate171inter7));
  inv1  gate723(.a(G549), .O(gate171inter8));
  nand2 gate724(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate725(.a(s_25), .b(gate171inter3), .O(gate171inter10));
  nor2  gate726(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate727(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate728(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2689(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2690(.a(gate173inter0), .b(s_306), .O(gate173inter1));
  and2  gate2691(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2692(.a(s_306), .O(gate173inter3));
  inv1  gate2693(.a(s_307), .O(gate173inter4));
  nand2 gate2694(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2695(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2696(.a(G486), .O(gate173inter7));
  inv1  gate2697(.a(G552), .O(gate173inter8));
  nand2 gate2698(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2699(.a(s_307), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2700(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2701(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2702(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate3011(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate3012(.a(gate175inter0), .b(s_352), .O(gate175inter1));
  and2  gate3013(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate3014(.a(s_352), .O(gate175inter3));
  inv1  gate3015(.a(s_353), .O(gate175inter4));
  nand2 gate3016(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate3017(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate3018(.a(G492), .O(gate175inter7));
  inv1  gate3019(.a(G555), .O(gate175inter8));
  nand2 gate3020(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate3021(.a(s_353), .b(gate175inter3), .O(gate175inter10));
  nor2  gate3022(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate3023(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate3024(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1149(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1150(.a(gate178inter0), .b(s_86), .O(gate178inter1));
  and2  gate1151(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1152(.a(s_86), .O(gate178inter3));
  inv1  gate1153(.a(s_87), .O(gate178inter4));
  nand2 gate1154(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1155(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1156(.a(G501), .O(gate178inter7));
  inv1  gate1157(.a(G558), .O(gate178inter8));
  nand2 gate1158(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1159(.a(s_87), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1160(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1161(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1162(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate1989(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1990(.a(gate179inter0), .b(s_206), .O(gate179inter1));
  and2  gate1991(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1992(.a(s_206), .O(gate179inter3));
  inv1  gate1993(.a(s_207), .O(gate179inter4));
  nand2 gate1994(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1995(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1996(.a(G504), .O(gate179inter7));
  inv1  gate1997(.a(G561), .O(gate179inter8));
  nand2 gate1998(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1999(.a(s_207), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2000(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2001(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2002(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1401(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1402(.a(gate180inter0), .b(s_122), .O(gate180inter1));
  and2  gate1403(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1404(.a(s_122), .O(gate180inter3));
  inv1  gate1405(.a(s_123), .O(gate180inter4));
  nand2 gate1406(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1407(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1408(.a(G507), .O(gate180inter7));
  inv1  gate1409(.a(G561), .O(gate180inter8));
  nand2 gate1410(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1411(.a(s_123), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1412(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1413(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1414(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1303(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1304(.a(gate181inter0), .b(s_108), .O(gate181inter1));
  and2  gate1305(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1306(.a(s_108), .O(gate181inter3));
  inv1  gate1307(.a(s_109), .O(gate181inter4));
  nand2 gate1308(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1309(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1310(.a(G510), .O(gate181inter7));
  inv1  gate1311(.a(G564), .O(gate181inter8));
  nand2 gate1312(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1313(.a(s_109), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1314(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1315(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1316(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1723(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1724(.a(gate182inter0), .b(s_168), .O(gate182inter1));
  and2  gate1725(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1726(.a(s_168), .O(gate182inter3));
  inv1  gate1727(.a(s_169), .O(gate182inter4));
  nand2 gate1728(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1729(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1730(.a(G513), .O(gate182inter7));
  inv1  gate1731(.a(G564), .O(gate182inter8));
  nand2 gate1732(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1733(.a(s_169), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1734(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1735(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1736(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2101(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2102(.a(gate185inter0), .b(s_222), .O(gate185inter1));
  and2  gate2103(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2104(.a(s_222), .O(gate185inter3));
  inv1  gate2105(.a(s_223), .O(gate185inter4));
  nand2 gate2106(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2107(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2108(.a(G570), .O(gate185inter7));
  inv1  gate2109(.a(G571), .O(gate185inter8));
  nand2 gate2110(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2111(.a(s_223), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2112(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2113(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2114(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1849(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1850(.a(gate187inter0), .b(s_186), .O(gate187inter1));
  and2  gate1851(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1852(.a(s_186), .O(gate187inter3));
  inv1  gate1853(.a(s_187), .O(gate187inter4));
  nand2 gate1854(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1855(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1856(.a(G574), .O(gate187inter7));
  inv1  gate1857(.a(G575), .O(gate187inter8));
  nand2 gate1858(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1859(.a(s_187), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1860(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1861(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1862(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate911(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate912(.a(gate192inter0), .b(s_52), .O(gate192inter1));
  and2  gate913(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate914(.a(s_52), .O(gate192inter3));
  inv1  gate915(.a(s_53), .O(gate192inter4));
  nand2 gate916(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate917(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate918(.a(G584), .O(gate192inter7));
  inv1  gate919(.a(G585), .O(gate192inter8));
  nand2 gate920(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate921(.a(s_53), .b(gate192inter3), .O(gate192inter10));
  nor2  gate922(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate923(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate924(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2549(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2550(.a(gate194inter0), .b(s_286), .O(gate194inter1));
  and2  gate2551(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2552(.a(s_286), .O(gate194inter3));
  inv1  gate2553(.a(s_287), .O(gate194inter4));
  nand2 gate2554(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2555(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2556(.a(G588), .O(gate194inter7));
  inv1  gate2557(.a(G589), .O(gate194inter8));
  nand2 gate2558(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2559(.a(s_287), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2560(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2561(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2562(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate2661(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2662(.a(gate196inter0), .b(s_302), .O(gate196inter1));
  and2  gate2663(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2664(.a(s_302), .O(gate196inter3));
  inv1  gate2665(.a(s_303), .O(gate196inter4));
  nand2 gate2666(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2667(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2668(.a(G592), .O(gate196inter7));
  inv1  gate2669(.a(G593), .O(gate196inter8));
  nand2 gate2670(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2671(.a(s_303), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2672(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2673(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2674(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1905(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1906(.a(gate197inter0), .b(s_194), .O(gate197inter1));
  and2  gate1907(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1908(.a(s_194), .O(gate197inter3));
  inv1  gate1909(.a(s_195), .O(gate197inter4));
  nand2 gate1910(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1911(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1912(.a(G594), .O(gate197inter7));
  inv1  gate1913(.a(G595), .O(gate197inter8));
  nand2 gate1914(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1915(.a(s_195), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1916(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1917(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1918(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2045(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2046(.a(gate207inter0), .b(s_214), .O(gate207inter1));
  and2  gate2047(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2048(.a(s_214), .O(gate207inter3));
  inv1  gate2049(.a(s_215), .O(gate207inter4));
  nand2 gate2050(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2051(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2052(.a(G622), .O(gate207inter7));
  inv1  gate2053(.a(G632), .O(gate207inter8));
  nand2 gate2054(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2055(.a(s_215), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2056(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2057(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2058(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1835(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1836(.a(gate209inter0), .b(s_184), .O(gate209inter1));
  and2  gate1837(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1838(.a(s_184), .O(gate209inter3));
  inv1  gate1839(.a(s_185), .O(gate209inter4));
  nand2 gate1840(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1841(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1842(.a(G602), .O(gate209inter7));
  inv1  gate1843(.a(G666), .O(gate209inter8));
  nand2 gate1844(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1845(.a(s_185), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1846(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1847(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1848(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate897(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate898(.a(gate215inter0), .b(s_50), .O(gate215inter1));
  and2  gate899(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate900(.a(s_50), .O(gate215inter3));
  inv1  gate901(.a(s_51), .O(gate215inter4));
  nand2 gate902(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate903(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate904(.a(G607), .O(gate215inter7));
  inv1  gate905(.a(G675), .O(gate215inter8));
  nand2 gate906(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate907(.a(s_51), .b(gate215inter3), .O(gate215inter10));
  nor2  gate908(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate909(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate910(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate2353(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2354(.a(gate216inter0), .b(s_258), .O(gate216inter1));
  and2  gate2355(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2356(.a(s_258), .O(gate216inter3));
  inv1  gate2357(.a(s_259), .O(gate216inter4));
  nand2 gate2358(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2359(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2360(.a(G617), .O(gate216inter7));
  inv1  gate2361(.a(G675), .O(gate216inter8));
  nand2 gate2362(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2363(.a(s_259), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2364(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2365(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2366(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2969(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2970(.a(gate217inter0), .b(s_346), .O(gate217inter1));
  and2  gate2971(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2972(.a(s_346), .O(gate217inter3));
  inv1  gate2973(.a(s_347), .O(gate217inter4));
  nand2 gate2974(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2975(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2976(.a(G622), .O(gate217inter7));
  inv1  gate2977(.a(G678), .O(gate217inter8));
  nand2 gate2978(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2979(.a(s_347), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2980(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2981(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2982(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1765(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1766(.a(gate218inter0), .b(s_174), .O(gate218inter1));
  and2  gate1767(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1768(.a(s_174), .O(gate218inter3));
  inv1  gate1769(.a(s_175), .O(gate218inter4));
  nand2 gate1770(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1771(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1772(.a(G627), .O(gate218inter7));
  inv1  gate1773(.a(G678), .O(gate218inter8));
  nand2 gate1774(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1775(.a(s_175), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1776(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1777(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1778(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate953(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate954(.a(gate220inter0), .b(s_58), .O(gate220inter1));
  and2  gate955(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate956(.a(s_58), .O(gate220inter3));
  inv1  gate957(.a(s_59), .O(gate220inter4));
  nand2 gate958(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate959(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate960(.a(G637), .O(gate220inter7));
  inv1  gate961(.a(G681), .O(gate220inter8));
  nand2 gate962(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate963(.a(s_59), .b(gate220inter3), .O(gate220inter10));
  nor2  gate964(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate965(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate966(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1667(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1668(.a(gate221inter0), .b(s_160), .O(gate221inter1));
  and2  gate1669(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1670(.a(s_160), .O(gate221inter3));
  inv1  gate1671(.a(s_161), .O(gate221inter4));
  nand2 gate1672(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1673(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1674(.a(G622), .O(gate221inter7));
  inv1  gate1675(.a(G684), .O(gate221inter8));
  nand2 gate1676(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1677(.a(s_161), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1678(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1679(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1680(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate3039(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate3040(.a(gate224inter0), .b(s_356), .O(gate224inter1));
  and2  gate3041(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate3042(.a(s_356), .O(gate224inter3));
  inv1  gate3043(.a(s_357), .O(gate224inter4));
  nand2 gate3044(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate3045(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate3046(.a(G637), .O(gate224inter7));
  inv1  gate3047(.a(G687), .O(gate224inter8));
  nand2 gate3048(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate3049(.a(s_357), .b(gate224inter3), .O(gate224inter10));
  nor2  gate3050(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate3051(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate3052(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate995(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate996(.a(gate225inter0), .b(s_64), .O(gate225inter1));
  and2  gate997(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate998(.a(s_64), .O(gate225inter3));
  inv1  gate999(.a(s_65), .O(gate225inter4));
  nand2 gate1000(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1001(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1002(.a(G690), .O(gate225inter7));
  inv1  gate1003(.a(G691), .O(gate225inter8));
  nand2 gate1004(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1005(.a(s_65), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1006(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1007(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1008(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1177(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1178(.a(gate227inter0), .b(s_90), .O(gate227inter1));
  and2  gate1179(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1180(.a(s_90), .O(gate227inter3));
  inv1  gate1181(.a(s_91), .O(gate227inter4));
  nand2 gate1182(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1183(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1184(.a(G694), .O(gate227inter7));
  inv1  gate1185(.a(G695), .O(gate227inter8));
  nand2 gate1186(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1187(.a(s_91), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1188(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1189(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1190(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate2983(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2984(.a(gate228inter0), .b(s_348), .O(gate228inter1));
  and2  gate2985(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2986(.a(s_348), .O(gate228inter3));
  inv1  gate2987(.a(s_349), .O(gate228inter4));
  nand2 gate2988(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2989(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2990(.a(G696), .O(gate228inter7));
  inv1  gate2991(.a(G697), .O(gate228inter8));
  nand2 gate2992(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2993(.a(s_349), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2994(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2995(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2996(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1457(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1458(.a(gate229inter0), .b(s_130), .O(gate229inter1));
  and2  gate1459(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1460(.a(s_130), .O(gate229inter3));
  inv1  gate1461(.a(s_131), .O(gate229inter4));
  nand2 gate1462(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1463(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1464(.a(G698), .O(gate229inter7));
  inv1  gate1465(.a(G699), .O(gate229inter8));
  nand2 gate1466(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1467(.a(s_131), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1468(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1469(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1470(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1639(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1640(.a(gate231inter0), .b(s_156), .O(gate231inter1));
  and2  gate1641(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1642(.a(s_156), .O(gate231inter3));
  inv1  gate1643(.a(s_157), .O(gate231inter4));
  nand2 gate1644(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1645(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1646(.a(G702), .O(gate231inter7));
  inv1  gate1647(.a(G703), .O(gate231inter8));
  nand2 gate1648(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1649(.a(s_157), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1650(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1651(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1652(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2591(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2592(.a(gate234inter0), .b(s_292), .O(gate234inter1));
  and2  gate2593(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2594(.a(s_292), .O(gate234inter3));
  inv1  gate2595(.a(s_293), .O(gate234inter4));
  nand2 gate2596(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2597(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2598(.a(G245), .O(gate234inter7));
  inv1  gate2599(.a(G721), .O(gate234inter8));
  nand2 gate2600(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2601(.a(s_293), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2602(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2603(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2604(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1583(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1584(.a(gate235inter0), .b(s_148), .O(gate235inter1));
  and2  gate1585(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1586(.a(s_148), .O(gate235inter3));
  inv1  gate1587(.a(s_149), .O(gate235inter4));
  nand2 gate1588(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1589(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1590(.a(G248), .O(gate235inter7));
  inv1  gate1591(.a(G724), .O(gate235inter8));
  nand2 gate1592(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1593(.a(s_149), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1594(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1595(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1596(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate925(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate926(.a(gate236inter0), .b(s_54), .O(gate236inter1));
  and2  gate927(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate928(.a(s_54), .O(gate236inter3));
  inv1  gate929(.a(s_55), .O(gate236inter4));
  nand2 gate930(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate931(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate932(.a(G251), .O(gate236inter7));
  inv1  gate933(.a(G727), .O(gate236inter8));
  nand2 gate934(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate935(.a(s_55), .b(gate236inter3), .O(gate236inter10));
  nor2  gate936(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate937(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate938(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2381(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2382(.a(gate238inter0), .b(s_262), .O(gate238inter1));
  and2  gate2383(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2384(.a(s_262), .O(gate238inter3));
  inv1  gate2385(.a(s_263), .O(gate238inter4));
  nand2 gate2386(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2387(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2388(.a(G257), .O(gate238inter7));
  inv1  gate2389(.a(G709), .O(gate238inter8));
  nand2 gate2390(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2391(.a(s_263), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2392(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2393(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2394(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2339(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2340(.a(gate241inter0), .b(s_256), .O(gate241inter1));
  and2  gate2341(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2342(.a(s_256), .O(gate241inter3));
  inv1  gate2343(.a(s_257), .O(gate241inter4));
  nand2 gate2344(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2345(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2346(.a(G242), .O(gate241inter7));
  inv1  gate2347(.a(G730), .O(gate241inter8));
  nand2 gate2348(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2349(.a(s_257), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2350(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2351(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2352(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1919(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1920(.a(gate242inter0), .b(s_196), .O(gate242inter1));
  and2  gate1921(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1922(.a(s_196), .O(gate242inter3));
  inv1  gate1923(.a(s_197), .O(gate242inter4));
  nand2 gate1924(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1925(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1926(.a(G718), .O(gate242inter7));
  inv1  gate1927(.a(G730), .O(gate242inter8));
  nand2 gate1928(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1929(.a(s_197), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1930(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1931(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1932(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2773(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2774(.a(gate246inter0), .b(s_318), .O(gate246inter1));
  and2  gate2775(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2776(.a(s_318), .O(gate246inter3));
  inv1  gate2777(.a(s_319), .O(gate246inter4));
  nand2 gate2778(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2779(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2780(.a(G724), .O(gate246inter7));
  inv1  gate2781(.a(G736), .O(gate246inter8));
  nand2 gate2782(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2783(.a(s_319), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2784(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2785(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2786(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1373(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1374(.a(gate258inter0), .b(s_118), .O(gate258inter1));
  and2  gate1375(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1376(.a(s_118), .O(gate258inter3));
  inv1  gate1377(.a(s_119), .O(gate258inter4));
  nand2 gate1378(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1379(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1380(.a(G756), .O(gate258inter7));
  inv1  gate1381(.a(G757), .O(gate258inter8));
  nand2 gate1382(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1383(.a(s_119), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1384(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1385(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1386(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1527(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1528(.a(gate260inter0), .b(s_140), .O(gate260inter1));
  and2  gate1529(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1530(.a(s_140), .O(gate260inter3));
  inv1  gate1531(.a(s_141), .O(gate260inter4));
  nand2 gate1532(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1533(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1534(.a(G760), .O(gate260inter7));
  inv1  gate1535(.a(G761), .O(gate260inter8));
  nand2 gate1536(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1537(.a(s_141), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1538(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1539(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1540(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2913(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2914(.a(gate262inter0), .b(s_338), .O(gate262inter1));
  and2  gate2915(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2916(.a(s_338), .O(gate262inter3));
  inv1  gate2917(.a(s_339), .O(gate262inter4));
  nand2 gate2918(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2919(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2920(.a(G764), .O(gate262inter7));
  inv1  gate2921(.a(G765), .O(gate262inter8));
  nand2 gate2922(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2923(.a(s_339), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2924(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2925(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2926(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1331(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1332(.a(gate263inter0), .b(s_112), .O(gate263inter1));
  and2  gate1333(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1334(.a(s_112), .O(gate263inter3));
  inv1  gate1335(.a(s_113), .O(gate263inter4));
  nand2 gate1336(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1337(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1338(.a(G766), .O(gate263inter7));
  inv1  gate1339(.a(G767), .O(gate263inter8));
  nand2 gate1340(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1341(.a(s_113), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1342(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1343(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1344(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1415(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1416(.a(gate265inter0), .b(s_124), .O(gate265inter1));
  and2  gate1417(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1418(.a(s_124), .O(gate265inter3));
  inv1  gate1419(.a(s_125), .O(gate265inter4));
  nand2 gate1420(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1421(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1422(.a(G642), .O(gate265inter7));
  inv1  gate1423(.a(G770), .O(gate265inter8));
  nand2 gate1424(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1425(.a(s_125), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1426(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1427(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1428(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate2143(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2144(.a(gate266inter0), .b(s_228), .O(gate266inter1));
  and2  gate2145(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2146(.a(s_228), .O(gate266inter3));
  inv1  gate2147(.a(s_229), .O(gate266inter4));
  nand2 gate2148(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2149(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2150(.a(G645), .O(gate266inter7));
  inv1  gate2151(.a(G773), .O(gate266inter8));
  nand2 gate2152(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2153(.a(s_229), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2154(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2155(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2156(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2535(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2536(.a(gate267inter0), .b(s_284), .O(gate267inter1));
  and2  gate2537(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2538(.a(s_284), .O(gate267inter3));
  inv1  gate2539(.a(s_285), .O(gate267inter4));
  nand2 gate2540(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2541(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2542(.a(G648), .O(gate267inter7));
  inv1  gate2543(.a(G776), .O(gate267inter8));
  nand2 gate2544(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2545(.a(s_285), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2546(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2547(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2548(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1009(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1010(.a(gate273inter0), .b(s_66), .O(gate273inter1));
  and2  gate1011(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1012(.a(s_66), .O(gate273inter3));
  inv1  gate1013(.a(s_67), .O(gate273inter4));
  nand2 gate1014(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1015(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1016(.a(G642), .O(gate273inter7));
  inv1  gate1017(.a(G794), .O(gate273inter8));
  nand2 gate1018(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1019(.a(s_67), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1020(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1021(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1022(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2311(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2312(.a(gate275inter0), .b(s_252), .O(gate275inter1));
  and2  gate2313(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2314(.a(s_252), .O(gate275inter3));
  inv1  gate2315(.a(s_253), .O(gate275inter4));
  nand2 gate2316(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2317(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2318(.a(G645), .O(gate275inter7));
  inv1  gate2319(.a(G797), .O(gate275inter8));
  nand2 gate2320(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2321(.a(s_253), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2322(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2323(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2324(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2843(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2844(.a(gate280inter0), .b(s_328), .O(gate280inter1));
  and2  gate2845(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2846(.a(s_328), .O(gate280inter3));
  inv1  gate2847(.a(s_329), .O(gate280inter4));
  nand2 gate2848(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2849(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2850(.a(G779), .O(gate280inter7));
  inv1  gate2851(.a(G803), .O(gate280inter8));
  nand2 gate2852(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2853(.a(s_329), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2854(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2855(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2856(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate2241(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2242(.a(gate281inter0), .b(s_242), .O(gate281inter1));
  and2  gate2243(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2244(.a(s_242), .O(gate281inter3));
  inv1  gate2245(.a(s_243), .O(gate281inter4));
  nand2 gate2246(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2247(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2248(.a(G654), .O(gate281inter7));
  inv1  gate2249(.a(G806), .O(gate281inter8));
  nand2 gate2250(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2251(.a(s_243), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2252(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2253(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2254(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate883(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate884(.a(gate282inter0), .b(s_48), .O(gate282inter1));
  and2  gate885(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate886(.a(s_48), .O(gate282inter3));
  inv1  gate887(.a(s_49), .O(gate282inter4));
  nand2 gate888(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate889(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate890(.a(G782), .O(gate282inter7));
  inv1  gate891(.a(G806), .O(gate282inter8));
  nand2 gate892(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate893(.a(s_49), .b(gate282inter3), .O(gate282inter10));
  nor2  gate894(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate895(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate896(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1135(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1136(.a(gate287inter0), .b(s_84), .O(gate287inter1));
  and2  gate1137(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1138(.a(s_84), .O(gate287inter3));
  inv1  gate1139(.a(s_85), .O(gate287inter4));
  nand2 gate1140(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1141(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1142(.a(G663), .O(gate287inter7));
  inv1  gate1143(.a(G815), .O(gate287inter8));
  nand2 gate1144(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1145(.a(s_85), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1146(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1147(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1148(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1709(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1710(.a(gate289inter0), .b(s_166), .O(gate289inter1));
  and2  gate1711(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1712(.a(s_166), .O(gate289inter3));
  inv1  gate1713(.a(s_167), .O(gate289inter4));
  nand2 gate1714(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1715(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1716(.a(G818), .O(gate289inter7));
  inv1  gate1717(.a(G819), .O(gate289inter8));
  nand2 gate1718(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1719(.a(s_167), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1720(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1721(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1722(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2619(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2620(.a(gate293inter0), .b(s_296), .O(gate293inter1));
  and2  gate2621(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2622(.a(s_296), .O(gate293inter3));
  inv1  gate2623(.a(s_297), .O(gate293inter4));
  nand2 gate2624(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2625(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2626(.a(G828), .O(gate293inter7));
  inv1  gate2627(.a(G829), .O(gate293inter8));
  nand2 gate2628(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2629(.a(s_297), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2630(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2631(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2632(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2675(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2676(.a(gate295inter0), .b(s_304), .O(gate295inter1));
  and2  gate2677(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2678(.a(s_304), .O(gate295inter3));
  inv1  gate2679(.a(s_305), .O(gate295inter4));
  nand2 gate2680(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2681(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2682(.a(G830), .O(gate295inter7));
  inv1  gate2683(.a(G831), .O(gate295inter8));
  nand2 gate2684(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2685(.a(s_305), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2686(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2687(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2688(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate659(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate660(.a(gate387inter0), .b(s_16), .O(gate387inter1));
  and2  gate661(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate662(.a(s_16), .O(gate387inter3));
  inv1  gate663(.a(s_17), .O(gate387inter4));
  nand2 gate664(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate665(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate666(.a(G1), .O(gate387inter7));
  inv1  gate667(.a(G1036), .O(gate387inter8));
  nand2 gate668(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate669(.a(s_17), .b(gate387inter3), .O(gate387inter10));
  nor2  gate670(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate671(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate672(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1947(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1948(.a(gate388inter0), .b(s_200), .O(gate388inter1));
  and2  gate1949(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1950(.a(s_200), .O(gate388inter3));
  inv1  gate1951(.a(s_201), .O(gate388inter4));
  nand2 gate1952(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1953(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1954(.a(G2), .O(gate388inter7));
  inv1  gate1955(.a(G1039), .O(gate388inter8));
  nand2 gate1956(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1957(.a(s_201), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1958(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1959(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1960(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate3053(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate3054(.a(gate393inter0), .b(s_358), .O(gate393inter1));
  and2  gate3055(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate3056(.a(s_358), .O(gate393inter3));
  inv1  gate3057(.a(s_359), .O(gate393inter4));
  nand2 gate3058(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate3059(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate3060(.a(G7), .O(gate393inter7));
  inv1  gate3061(.a(G1054), .O(gate393inter8));
  nand2 gate3062(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate3063(.a(s_359), .b(gate393inter3), .O(gate393inter10));
  nor2  gate3064(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate3065(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate3066(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2493(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2494(.a(gate394inter0), .b(s_278), .O(gate394inter1));
  and2  gate2495(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2496(.a(s_278), .O(gate394inter3));
  inv1  gate2497(.a(s_279), .O(gate394inter4));
  nand2 gate2498(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2499(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2500(.a(G8), .O(gate394inter7));
  inv1  gate2501(.a(G1057), .O(gate394inter8));
  nand2 gate2502(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2503(.a(s_279), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2504(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2505(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2506(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1597(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1598(.a(gate395inter0), .b(s_150), .O(gate395inter1));
  and2  gate1599(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1600(.a(s_150), .O(gate395inter3));
  inv1  gate1601(.a(s_151), .O(gate395inter4));
  nand2 gate1602(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1603(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1604(.a(G9), .O(gate395inter7));
  inv1  gate1605(.a(G1060), .O(gate395inter8));
  nand2 gate1606(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1607(.a(s_151), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1608(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1609(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1610(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2563(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2564(.a(gate397inter0), .b(s_288), .O(gate397inter1));
  and2  gate2565(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2566(.a(s_288), .O(gate397inter3));
  inv1  gate2567(.a(s_289), .O(gate397inter4));
  nand2 gate2568(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2569(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2570(.a(G11), .O(gate397inter7));
  inv1  gate2571(.a(G1066), .O(gate397inter8));
  nand2 gate2572(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2573(.a(s_289), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2574(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2575(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2576(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1569(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1570(.a(gate403inter0), .b(s_146), .O(gate403inter1));
  and2  gate1571(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1572(.a(s_146), .O(gate403inter3));
  inv1  gate1573(.a(s_147), .O(gate403inter4));
  nand2 gate1574(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1575(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1576(.a(G17), .O(gate403inter7));
  inv1  gate1577(.a(G1084), .O(gate403inter8));
  nand2 gate1578(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1579(.a(s_147), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1580(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1581(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1582(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate2213(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2214(.a(gate404inter0), .b(s_238), .O(gate404inter1));
  and2  gate2215(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2216(.a(s_238), .O(gate404inter3));
  inv1  gate2217(.a(s_239), .O(gate404inter4));
  nand2 gate2218(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2219(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2220(.a(G18), .O(gate404inter7));
  inv1  gate2221(.a(G1087), .O(gate404inter8));
  nand2 gate2222(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2223(.a(s_239), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2224(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2225(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2226(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate2423(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2424(.a(gate405inter0), .b(s_268), .O(gate405inter1));
  and2  gate2425(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2426(.a(s_268), .O(gate405inter3));
  inv1  gate2427(.a(s_269), .O(gate405inter4));
  nand2 gate2428(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2429(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2430(.a(G19), .O(gate405inter7));
  inv1  gate2431(.a(G1090), .O(gate405inter8));
  nand2 gate2432(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2433(.a(s_269), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2434(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2435(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2436(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate3123(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate3124(.a(gate408inter0), .b(s_368), .O(gate408inter1));
  and2  gate3125(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate3126(.a(s_368), .O(gate408inter3));
  inv1  gate3127(.a(s_369), .O(gate408inter4));
  nand2 gate3128(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate3129(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate3130(.a(G22), .O(gate408inter7));
  inv1  gate3131(.a(G1099), .O(gate408inter8));
  nand2 gate3132(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate3133(.a(s_369), .b(gate408inter3), .O(gate408inter10));
  nor2  gate3134(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate3135(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate3136(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate2759(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2760(.a(gate409inter0), .b(s_316), .O(gate409inter1));
  and2  gate2761(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2762(.a(s_316), .O(gate409inter3));
  inv1  gate2763(.a(s_317), .O(gate409inter4));
  nand2 gate2764(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2765(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2766(.a(G23), .O(gate409inter7));
  inv1  gate2767(.a(G1102), .O(gate409inter8));
  nand2 gate2768(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2769(.a(s_317), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2770(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2771(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2772(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate799(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate800(.a(gate410inter0), .b(s_36), .O(gate410inter1));
  and2  gate801(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate802(.a(s_36), .O(gate410inter3));
  inv1  gate803(.a(s_37), .O(gate410inter4));
  nand2 gate804(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate805(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate806(.a(G24), .O(gate410inter7));
  inv1  gate807(.a(G1105), .O(gate410inter8));
  nand2 gate808(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate809(.a(s_37), .b(gate410inter3), .O(gate410inter10));
  nor2  gate810(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate811(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate812(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate841(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate842(.a(gate411inter0), .b(s_42), .O(gate411inter1));
  and2  gate843(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate844(.a(s_42), .O(gate411inter3));
  inv1  gate845(.a(s_43), .O(gate411inter4));
  nand2 gate846(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate847(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate848(.a(G25), .O(gate411inter7));
  inv1  gate849(.a(G1108), .O(gate411inter8));
  nand2 gate850(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate851(.a(s_43), .b(gate411inter3), .O(gate411inter10));
  nor2  gate852(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate853(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate854(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1093(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1094(.a(gate415inter0), .b(s_78), .O(gate415inter1));
  and2  gate1095(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1096(.a(s_78), .O(gate415inter3));
  inv1  gate1097(.a(s_79), .O(gate415inter4));
  nand2 gate1098(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1099(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1100(.a(G29), .O(gate415inter7));
  inv1  gate1101(.a(G1120), .O(gate415inter8));
  nand2 gate1102(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1103(.a(s_79), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1104(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1105(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1106(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1107(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1108(.a(gate420inter0), .b(s_80), .O(gate420inter1));
  and2  gate1109(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1110(.a(s_80), .O(gate420inter3));
  inv1  gate1111(.a(s_81), .O(gate420inter4));
  nand2 gate1112(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1113(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1114(.a(G1036), .O(gate420inter7));
  inv1  gate1115(.a(G1132), .O(gate420inter8));
  nand2 gate1116(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1117(.a(s_81), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1118(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1119(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1120(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1499(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1500(.a(gate421inter0), .b(s_136), .O(gate421inter1));
  and2  gate1501(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1502(.a(s_136), .O(gate421inter3));
  inv1  gate1503(.a(s_137), .O(gate421inter4));
  nand2 gate1504(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1505(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1506(.a(G2), .O(gate421inter7));
  inv1  gate1507(.a(G1135), .O(gate421inter8));
  nand2 gate1508(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1509(.a(s_137), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1510(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1511(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1512(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1779(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1780(.a(gate422inter0), .b(s_176), .O(gate422inter1));
  and2  gate1781(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1782(.a(s_176), .O(gate422inter3));
  inv1  gate1783(.a(s_177), .O(gate422inter4));
  nand2 gate1784(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1785(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1786(.a(G1039), .O(gate422inter7));
  inv1  gate1787(.a(G1135), .O(gate422inter8));
  nand2 gate1788(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1789(.a(s_177), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1790(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1791(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1792(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2955(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2956(.a(gate428inter0), .b(s_344), .O(gate428inter1));
  and2  gate2957(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2958(.a(s_344), .O(gate428inter3));
  inv1  gate2959(.a(s_345), .O(gate428inter4));
  nand2 gate2960(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2961(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2962(.a(G1048), .O(gate428inter7));
  inv1  gate2963(.a(G1144), .O(gate428inter8));
  nand2 gate2964(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2965(.a(s_345), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2966(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2967(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2968(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1807(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1808(.a(gate437inter0), .b(s_180), .O(gate437inter1));
  and2  gate1809(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1810(.a(s_180), .O(gate437inter3));
  inv1  gate1811(.a(s_181), .O(gate437inter4));
  nand2 gate1812(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1813(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1814(.a(G10), .O(gate437inter7));
  inv1  gate1815(.a(G1159), .O(gate437inter8));
  nand2 gate1816(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1817(.a(s_181), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1818(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1819(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1820(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1877(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1878(.a(gate441inter0), .b(s_190), .O(gate441inter1));
  and2  gate1879(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1880(.a(s_190), .O(gate441inter3));
  inv1  gate1881(.a(s_191), .O(gate441inter4));
  nand2 gate1882(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1883(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1884(.a(G12), .O(gate441inter7));
  inv1  gate1885(.a(G1165), .O(gate441inter8));
  nand2 gate1886(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1887(.a(s_191), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1888(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1889(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1890(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1653(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1654(.a(gate445inter0), .b(s_158), .O(gate445inter1));
  and2  gate1655(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1656(.a(s_158), .O(gate445inter3));
  inv1  gate1657(.a(s_159), .O(gate445inter4));
  nand2 gate1658(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1659(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1660(.a(G14), .O(gate445inter7));
  inv1  gate1661(.a(G1171), .O(gate445inter8));
  nand2 gate1662(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1663(.a(s_159), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1664(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1665(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1666(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate2031(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2032(.a(gate446inter0), .b(s_212), .O(gate446inter1));
  and2  gate2033(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2034(.a(s_212), .O(gate446inter3));
  inv1  gate2035(.a(s_213), .O(gate446inter4));
  nand2 gate2036(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2037(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2038(.a(G1075), .O(gate446inter7));
  inv1  gate2039(.a(G1171), .O(gate446inter8));
  nand2 gate2040(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2041(.a(s_213), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2042(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2043(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2044(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1793(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1794(.a(gate448inter0), .b(s_178), .O(gate448inter1));
  and2  gate1795(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1796(.a(s_178), .O(gate448inter3));
  inv1  gate1797(.a(s_179), .O(gate448inter4));
  nand2 gate1798(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1799(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1800(.a(G1078), .O(gate448inter7));
  inv1  gate1801(.a(G1174), .O(gate448inter8));
  nand2 gate1802(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1803(.a(s_179), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1804(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1805(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1806(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1289(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1290(.a(gate449inter0), .b(s_106), .O(gate449inter1));
  and2  gate1291(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1292(.a(s_106), .O(gate449inter3));
  inv1  gate1293(.a(s_107), .O(gate449inter4));
  nand2 gate1294(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1295(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1296(.a(G16), .O(gate449inter7));
  inv1  gate1297(.a(G1177), .O(gate449inter8));
  nand2 gate1298(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1299(.a(s_107), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1300(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1301(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1302(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1471(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1472(.a(gate450inter0), .b(s_132), .O(gate450inter1));
  and2  gate1473(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1474(.a(s_132), .O(gate450inter3));
  inv1  gate1475(.a(s_133), .O(gate450inter4));
  nand2 gate1476(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1477(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1478(.a(G1081), .O(gate450inter7));
  inv1  gate1479(.a(G1177), .O(gate450inter8));
  nand2 gate1480(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1481(.a(s_133), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1482(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1483(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1484(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2325(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2326(.a(gate452inter0), .b(s_254), .O(gate452inter1));
  and2  gate2327(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2328(.a(s_254), .O(gate452inter3));
  inv1  gate2329(.a(s_255), .O(gate452inter4));
  nand2 gate2330(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2331(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2332(.a(G1084), .O(gate452inter7));
  inv1  gate2333(.a(G1180), .O(gate452inter8));
  nand2 gate2334(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2335(.a(s_255), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2336(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2337(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2338(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate575(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate576(.a(gate455inter0), .b(s_4), .O(gate455inter1));
  and2  gate577(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate578(.a(s_4), .O(gate455inter3));
  inv1  gate579(.a(s_5), .O(gate455inter4));
  nand2 gate580(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate581(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate582(.a(G19), .O(gate455inter7));
  inv1  gate583(.a(G1186), .O(gate455inter8));
  nand2 gate584(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate585(.a(s_5), .b(gate455inter3), .O(gate455inter10));
  nor2  gate586(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate587(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate588(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate589(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate590(.a(gate460inter0), .b(s_6), .O(gate460inter1));
  and2  gate591(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate592(.a(s_6), .O(gate460inter3));
  inv1  gate593(.a(s_7), .O(gate460inter4));
  nand2 gate594(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate595(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate596(.a(G1096), .O(gate460inter7));
  inv1  gate597(.a(G1192), .O(gate460inter8));
  nand2 gate598(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate599(.a(s_7), .b(gate460inter3), .O(gate460inter10));
  nor2  gate600(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate601(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate602(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2367(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2368(.a(gate466inter0), .b(s_260), .O(gate466inter1));
  and2  gate2369(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2370(.a(s_260), .O(gate466inter3));
  inv1  gate2371(.a(s_261), .O(gate466inter4));
  nand2 gate2372(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2373(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2374(.a(G1105), .O(gate466inter7));
  inv1  gate2375(.a(G1201), .O(gate466inter8));
  nand2 gate2376(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2377(.a(s_261), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2378(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2379(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2380(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate701(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate702(.a(gate467inter0), .b(s_22), .O(gate467inter1));
  and2  gate703(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate704(.a(s_22), .O(gate467inter3));
  inv1  gate705(.a(s_23), .O(gate467inter4));
  nand2 gate706(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate707(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate708(.a(G25), .O(gate467inter7));
  inv1  gate709(.a(G1204), .O(gate467inter8));
  nand2 gate710(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate711(.a(s_23), .b(gate467inter3), .O(gate467inter10));
  nor2  gate712(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate713(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate714(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2871(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2872(.a(gate471inter0), .b(s_332), .O(gate471inter1));
  and2  gate2873(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2874(.a(s_332), .O(gate471inter3));
  inv1  gate2875(.a(s_333), .O(gate471inter4));
  nand2 gate2876(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2877(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2878(.a(G27), .O(gate471inter7));
  inv1  gate2879(.a(G1210), .O(gate471inter8));
  nand2 gate2880(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2881(.a(s_333), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2882(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2883(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2884(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2829(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2830(.a(gate472inter0), .b(s_326), .O(gate472inter1));
  and2  gate2831(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2832(.a(s_326), .O(gate472inter3));
  inv1  gate2833(.a(s_327), .O(gate472inter4));
  nand2 gate2834(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2835(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2836(.a(G1114), .O(gate472inter7));
  inv1  gate2837(.a(G1210), .O(gate472inter8));
  nand2 gate2838(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2839(.a(s_327), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2840(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2841(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2842(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2927(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2928(.a(gate474inter0), .b(s_340), .O(gate474inter1));
  and2  gate2929(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2930(.a(s_340), .O(gate474inter3));
  inv1  gate2931(.a(s_341), .O(gate474inter4));
  nand2 gate2932(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2933(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2934(.a(G1117), .O(gate474inter7));
  inv1  gate2935(.a(G1213), .O(gate474inter8));
  nand2 gate2936(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2937(.a(s_341), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2938(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2939(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2940(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate2059(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2060(.a(gate475inter0), .b(s_216), .O(gate475inter1));
  and2  gate2061(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2062(.a(s_216), .O(gate475inter3));
  inv1  gate2063(.a(s_217), .O(gate475inter4));
  nand2 gate2064(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2065(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2066(.a(G29), .O(gate475inter7));
  inv1  gate2067(.a(G1216), .O(gate475inter8));
  nand2 gate2068(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2069(.a(s_217), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2070(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2071(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2072(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1191(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1192(.a(gate476inter0), .b(s_92), .O(gate476inter1));
  and2  gate1193(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1194(.a(s_92), .O(gate476inter3));
  inv1  gate1195(.a(s_93), .O(gate476inter4));
  nand2 gate1196(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1197(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1198(.a(G1120), .O(gate476inter7));
  inv1  gate1199(.a(G1216), .O(gate476inter8));
  nand2 gate1200(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1201(.a(s_93), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1202(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1203(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1204(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate2507(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2508(.a(gate477inter0), .b(s_280), .O(gate477inter1));
  and2  gate2509(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2510(.a(s_280), .O(gate477inter3));
  inv1  gate2511(.a(s_281), .O(gate477inter4));
  nand2 gate2512(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2513(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2514(.a(G30), .O(gate477inter7));
  inv1  gate2515(.a(G1219), .O(gate477inter8));
  nand2 gate2516(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2517(.a(s_281), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2518(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2519(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2520(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate2465(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2466(.a(gate481inter0), .b(s_274), .O(gate481inter1));
  and2  gate2467(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2468(.a(s_274), .O(gate481inter3));
  inv1  gate2469(.a(s_275), .O(gate481inter4));
  nand2 gate2470(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2471(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2472(.a(G32), .O(gate481inter7));
  inv1  gate2473(.a(G1225), .O(gate481inter8));
  nand2 gate2474(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2475(.a(s_275), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2476(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2477(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2478(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate2451(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2452(.a(gate482inter0), .b(s_272), .O(gate482inter1));
  and2  gate2453(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2454(.a(s_272), .O(gate482inter3));
  inv1  gate2455(.a(s_273), .O(gate482inter4));
  nand2 gate2456(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2457(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2458(.a(G1129), .O(gate482inter7));
  inv1  gate2459(.a(G1225), .O(gate482inter8));
  nand2 gate2460(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2461(.a(s_273), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2462(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2463(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2464(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1863(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1864(.a(gate483inter0), .b(s_188), .O(gate483inter1));
  and2  gate1865(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1866(.a(s_188), .O(gate483inter3));
  inv1  gate1867(.a(s_189), .O(gate483inter4));
  nand2 gate1868(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1869(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1870(.a(G1228), .O(gate483inter7));
  inv1  gate1871(.a(G1229), .O(gate483inter8));
  nand2 gate1872(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1873(.a(s_189), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1874(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1875(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1876(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate939(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate940(.a(gate485inter0), .b(s_56), .O(gate485inter1));
  and2  gate941(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate942(.a(s_56), .O(gate485inter3));
  inv1  gate943(.a(s_57), .O(gate485inter4));
  nand2 gate944(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate945(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate946(.a(G1232), .O(gate485inter7));
  inv1  gate947(.a(G1233), .O(gate485inter8));
  nand2 gate948(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate949(.a(s_57), .b(gate485inter3), .O(gate485inter10));
  nor2  gate950(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate951(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate952(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate2801(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2802(.a(gate487inter0), .b(s_322), .O(gate487inter1));
  and2  gate2803(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2804(.a(s_322), .O(gate487inter3));
  inv1  gate2805(.a(s_323), .O(gate487inter4));
  nand2 gate2806(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2807(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2808(.a(G1236), .O(gate487inter7));
  inv1  gate2809(.a(G1237), .O(gate487inter8));
  nand2 gate2810(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2811(.a(s_323), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2812(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2813(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2814(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2647(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2648(.a(gate490inter0), .b(s_300), .O(gate490inter1));
  and2  gate2649(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2650(.a(s_300), .O(gate490inter3));
  inv1  gate2651(.a(s_301), .O(gate490inter4));
  nand2 gate2652(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2653(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2654(.a(G1242), .O(gate490inter7));
  inv1  gate2655(.a(G1243), .O(gate490inter8));
  nand2 gate2656(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2657(.a(s_301), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2658(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2659(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2660(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1485(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1486(.a(gate497inter0), .b(s_134), .O(gate497inter1));
  and2  gate1487(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1488(.a(s_134), .O(gate497inter3));
  inv1  gate1489(.a(s_135), .O(gate497inter4));
  nand2 gate1490(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1491(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1492(.a(G1256), .O(gate497inter7));
  inv1  gate1493(.a(G1257), .O(gate497inter8));
  nand2 gate1494(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1495(.a(s_135), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1496(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1497(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1498(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate743(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate744(.a(gate499inter0), .b(s_28), .O(gate499inter1));
  and2  gate745(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate746(.a(s_28), .O(gate499inter3));
  inv1  gate747(.a(s_29), .O(gate499inter4));
  nand2 gate748(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate749(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate750(.a(G1260), .O(gate499inter7));
  inv1  gate751(.a(G1261), .O(gate499inter8));
  nand2 gate752(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate753(.a(s_29), .b(gate499inter3), .O(gate499inter10));
  nor2  gate754(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate755(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate756(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1037(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1038(.a(gate500inter0), .b(s_70), .O(gate500inter1));
  and2  gate1039(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1040(.a(s_70), .O(gate500inter3));
  inv1  gate1041(.a(s_71), .O(gate500inter4));
  nand2 gate1042(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1043(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1044(.a(G1262), .O(gate500inter7));
  inv1  gate1045(.a(G1263), .O(gate500inter8));
  nand2 gate1046(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1047(.a(s_71), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1048(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1049(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1050(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1023(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1024(.a(gate502inter0), .b(s_68), .O(gate502inter1));
  and2  gate1025(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1026(.a(s_68), .O(gate502inter3));
  inv1  gate1027(.a(s_69), .O(gate502inter4));
  nand2 gate1028(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1029(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1030(.a(G1266), .O(gate502inter7));
  inv1  gate1031(.a(G1267), .O(gate502inter8));
  nand2 gate1032(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1033(.a(s_69), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1034(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1035(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1036(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1065(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1066(.a(gate506inter0), .b(s_74), .O(gate506inter1));
  and2  gate1067(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1068(.a(s_74), .O(gate506inter3));
  inv1  gate1069(.a(s_75), .O(gate506inter4));
  nand2 gate1070(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1071(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1072(.a(G1274), .O(gate506inter7));
  inv1  gate1073(.a(G1275), .O(gate506inter8));
  nand2 gate1074(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1075(.a(s_75), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1076(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1077(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1078(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2297(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2298(.a(gate508inter0), .b(s_250), .O(gate508inter1));
  and2  gate2299(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2300(.a(s_250), .O(gate508inter3));
  inv1  gate2301(.a(s_251), .O(gate508inter4));
  nand2 gate2302(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2303(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2304(.a(G1278), .O(gate508inter7));
  inv1  gate2305(.a(G1279), .O(gate508inter8));
  nand2 gate2306(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2307(.a(s_251), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2308(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2309(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2310(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2745(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2746(.a(gate510inter0), .b(s_314), .O(gate510inter1));
  and2  gate2747(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2748(.a(s_314), .O(gate510inter3));
  inv1  gate2749(.a(s_315), .O(gate510inter4));
  nand2 gate2750(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2751(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2752(.a(G1282), .O(gate510inter7));
  inv1  gate2753(.a(G1283), .O(gate510inter8));
  nand2 gate2754(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2755(.a(s_315), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2756(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2757(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2758(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate2731(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2732(.a(gate511inter0), .b(s_312), .O(gate511inter1));
  and2  gate2733(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2734(.a(s_312), .O(gate511inter3));
  inv1  gate2735(.a(s_313), .O(gate511inter4));
  nand2 gate2736(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2737(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2738(.a(G1284), .O(gate511inter7));
  inv1  gate2739(.a(G1285), .O(gate511inter8));
  nand2 gate2740(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2741(.a(s_313), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2742(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2743(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2744(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate981(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate982(.a(gate512inter0), .b(s_62), .O(gate512inter1));
  and2  gate983(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate984(.a(s_62), .O(gate512inter3));
  inv1  gate985(.a(s_63), .O(gate512inter4));
  nand2 gate986(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate987(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate988(.a(G1286), .O(gate512inter7));
  inv1  gate989(.a(G1287), .O(gate512inter8));
  nand2 gate990(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate991(.a(s_63), .b(gate512inter3), .O(gate512inter10));
  nor2  gate992(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate993(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate994(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule