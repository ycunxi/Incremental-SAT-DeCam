module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1093(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1094(.a(gate15inter0), .b(s_78), .O(gate15inter1));
  and2  gate1095(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1096(.a(s_78), .O(gate15inter3));
  inv1  gate1097(.a(s_79), .O(gate15inter4));
  nand2 gate1098(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1099(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1100(.a(G13), .O(gate15inter7));
  inv1  gate1101(.a(G14), .O(gate15inter8));
  nand2 gate1102(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1103(.a(s_79), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1104(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1105(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1106(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1219(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1220(.a(gate21inter0), .b(s_96), .O(gate21inter1));
  and2  gate1221(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1222(.a(s_96), .O(gate21inter3));
  inv1  gate1223(.a(s_97), .O(gate21inter4));
  nand2 gate1224(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1225(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1226(.a(G25), .O(gate21inter7));
  inv1  gate1227(.a(G26), .O(gate21inter8));
  nand2 gate1228(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1229(.a(s_97), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1230(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1231(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1232(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1681(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1682(.a(gate27inter0), .b(s_162), .O(gate27inter1));
  and2  gate1683(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1684(.a(s_162), .O(gate27inter3));
  inv1  gate1685(.a(s_163), .O(gate27inter4));
  nand2 gate1686(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1687(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1688(.a(G2), .O(gate27inter7));
  inv1  gate1689(.a(G6), .O(gate27inter8));
  nand2 gate1690(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1691(.a(s_163), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1692(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1693(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1694(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1135(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1136(.a(gate35inter0), .b(s_84), .O(gate35inter1));
  and2  gate1137(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1138(.a(s_84), .O(gate35inter3));
  inv1  gate1139(.a(s_85), .O(gate35inter4));
  nand2 gate1140(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1141(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1142(.a(G18), .O(gate35inter7));
  inv1  gate1143(.a(G22), .O(gate35inter8));
  nand2 gate1144(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1145(.a(s_85), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1146(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1147(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1148(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1485(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1486(.a(gate37inter0), .b(s_134), .O(gate37inter1));
  and2  gate1487(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1488(.a(s_134), .O(gate37inter3));
  inv1  gate1489(.a(s_135), .O(gate37inter4));
  nand2 gate1490(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1491(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1492(.a(G19), .O(gate37inter7));
  inv1  gate1493(.a(G23), .O(gate37inter8));
  nand2 gate1494(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1495(.a(s_135), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1496(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1497(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1498(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1121(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1122(.a(gate40inter0), .b(s_82), .O(gate40inter1));
  and2  gate1123(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1124(.a(s_82), .O(gate40inter3));
  inv1  gate1125(.a(s_83), .O(gate40inter4));
  nand2 gate1126(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1127(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1128(.a(G28), .O(gate40inter7));
  inv1  gate1129(.a(G32), .O(gate40inter8));
  nand2 gate1130(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1131(.a(s_83), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1132(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1133(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1134(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1065(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1066(.a(gate43inter0), .b(s_74), .O(gate43inter1));
  and2  gate1067(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1068(.a(s_74), .O(gate43inter3));
  inv1  gate1069(.a(s_75), .O(gate43inter4));
  nand2 gate1070(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1071(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1072(.a(G3), .O(gate43inter7));
  inv1  gate1073(.a(G269), .O(gate43inter8));
  nand2 gate1074(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1075(.a(s_75), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1076(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1077(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1078(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate897(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate898(.a(gate45inter0), .b(s_50), .O(gate45inter1));
  and2  gate899(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate900(.a(s_50), .O(gate45inter3));
  inv1  gate901(.a(s_51), .O(gate45inter4));
  nand2 gate902(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate903(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate904(.a(G5), .O(gate45inter7));
  inv1  gate905(.a(G272), .O(gate45inter8));
  nand2 gate906(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate907(.a(s_51), .b(gate45inter3), .O(gate45inter10));
  nor2  gate908(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate909(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate910(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate743(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate744(.a(gate49inter0), .b(s_28), .O(gate49inter1));
  and2  gate745(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate746(.a(s_28), .O(gate49inter3));
  inv1  gate747(.a(s_29), .O(gate49inter4));
  nand2 gate748(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate749(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate750(.a(G9), .O(gate49inter7));
  inv1  gate751(.a(G278), .O(gate49inter8));
  nand2 gate752(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate753(.a(s_29), .b(gate49inter3), .O(gate49inter10));
  nor2  gate754(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate755(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate756(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1653(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1654(.a(gate50inter0), .b(s_158), .O(gate50inter1));
  and2  gate1655(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1656(.a(s_158), .O(gate50inter3));
  inv1  gate1657(.a(s_159), .O(gate50inter4));
  nand2 gate1658(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1659(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1660(.a(G10), .O(gate50inter7));
  inv1  gate1661(.a(G278), .O(gate50inter8));
  nand2 gate1662(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1663(.a(s_159), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1664(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1665(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1666(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1261(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1262(.a(gate51inter0), .b(s_102), .O(gate51inter1));
  and2  gate1263(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1264(.a(s_102), .O(gate51inter3));
  inv1  gate1265(.a(s_103), .O(gate51inter4));
  nand2 gate1266(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1267(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1268(.a(G11), .O(gate51inter7));
  inv1  gate1269(.a(G281), .O(gate51inter8));
  nand2 gate1270(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1271(.a(s_103), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1272(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1273(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1274(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1373(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1374(.a(gate57inter0), .b(s_118), .O(gate57inter1));
  and2  gate1375(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1376(.a(s_118), .O(gate57inter3));
  inv1  gate1377(.a(s_119), .O(gate57inter4));
  nand2 gate1378(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1379(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1380(.a(G17), .O(gate57inter7));
  inv1  gate1381(.a(G290), .O(gate57inter8));
  nand2 gate1382(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1383(.a(s_119), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1384(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1385(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1386(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1443(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1444(.a(gate68inter0), .b(s_128), .O(gate68inter1));
  and2  gate1445(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1446(.a(s_128), .O(gate68inter3));
  inv1  gate1447(.a(s_129), .O(gate68inter4));
  nand2 gate1448(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1449(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1450(.a(G28), .O(gate68inter7));
  inv1  gate1451(.a(G305), .O(gate68inter8));
  nand2 gate1452(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1453(.a(s_129), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1454(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1455(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1456(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1303(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1304(.a(gate74inter0), .b(s_108), .O(gate74inter1));
  and2  gate1305(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1306(.a(s_108), .O(gate74inter3));
  inv1  gate1307(.a(s_109), .O(gate74inter4));
  nand2 gate1308(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1309(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1310(.a(G5), .O(gate74inter7));
  inv1  gate1311(.a(G314), .O(gate74inter8));
  nand2 gate1312(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1313(.a(s_109), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1314(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1315(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1316(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1723(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1724(.a(gate80inter0), .b(s_168), .O(gate80inter1));
  and2  gate1725(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1726(.a(s_168), .O(gate80inter3));
  inv1  gate1727(.a(s_169), .O(gate80inter4));
  nand2 gate1728(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1729(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1730(.a(G14), .O(gate80inter7));
  inv1  gate1731(.a(G323), .O(gate80inter8));
  nand2 gate1732(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1733(.a(s_169), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1734(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1735(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1736(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1037(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1038(.a(gate85inter0), .b(s_70), .O(gate85inter1));
  and2  gate1039(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1040(.a(s_70), .O(gate85inter3));
  inv1  gate1041(.a(s_71), .O(gate85inter4));
  nand2 gate1042(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1043(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1044(.a(G4), .O(gate85inter7));
  inv1  gate1045(.a(G332), .O(gate85inter8));
  nand2 gate1046(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1047(.a(s_71), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1048(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1049(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1050(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate911(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate912(.a(gate86inter0), .b(s_52), .O(gate86inter1));
  and2  gate913(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate914(.a(s_52), .O(gate86inter3));
  inv1  gate915(.a(s_53), .O(gate86inter4));
  nand2 gate916(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate917(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate918(.a(G8), .O(gate86inter7));
  inv1  gate919(.a(G332), .O(gate86inter8));
  nand2 gate920(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate921(.a(s_53), .b(gate86inter3), .O(gate86inter10));
  nor2  gate922(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate923(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate924(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1695(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1696(.a(gate93inter0), .b(s_164), .O(gate93inter1));
  and2  gate1697(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1698(.a(s_164), .O(gate93inter3));
  inv1  gate1699(.a(s_165), .O(gate93inter4));
  nand2 gate1700(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1701(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1702(.a(G18), .O(gate93inter7));
  inv1  gate1703(.a(G344), .O(gate93inter8));
  nand2 gate1704(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1705(.a(s_165), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1706(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1707(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1708(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1177(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1178(.a(gate96inter0), .b(s_90), .O(gate96inter1));
  and2  gate1179(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1180(.a(s_90), .O(gate96inter3));
  inv1  gate1181(.a(s_91), .O(gate96inter4));
  nand2 gate1182(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1183(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1184(.a(G30), .O(gate96inter7));
  inv1  gate1185(.a(G347), .O(gate96inter8));
  nand2 gate1186(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1187(.a(s_91), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1188(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1189(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1190(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate967(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate968(.a(gate97inter0), .b(s_60), .O(gate97inter1));
  and2  gate969(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate970(.a(s_60), .O(gate97inter3));
  inv1  gate971(.a(s_61), .O(gate97inter4));
  nand2 gate972(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate973(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate974(.a(G19), .O(gate97inter7));
  inv1  gate975(.a(G350), .O(gate97inter8));
  nand2 gate976(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate977(.a(s_61), .b(gate97inter3), .O(gate97inter10));
  nor2  gate978(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate979(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate980(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate547(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate548(.a(gate98inter0), .b(s_0), .O(gate98inter1));
  and2  gate549(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate550(.a(s_0), .O(gate98inter3));
  inv1  gate551(.a(s_1), .O(gate98inter4));
  nand2 gate552(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate553(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate554(.a(G23), .O(gate98inter7));
  inv1  gate555(.a(G350), .O(gate98inter8));
  nand2 gate556(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate557(.a(s_1), .b(gate98inter3), .O(gate98inter10));
  nor2  gate558(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate559(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate560(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate701(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate702(.a(gate100inter0), .b(s_22), .O(gate100inter1));
  and2  gate703(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate704(.a(s_22), .O(gate100inter3));
  inv1  gate705(.a(s_23), .O(gate100inter4));
  nand2 gate706(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate707(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate708(.a(G31), .O(gate100inter7));
  inv1  gate709(.a(G353), .O(gate100inter8));
  nand2 gate710(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate711(.a(s_23), .b(gate100inter3), .O(gate100inter10));
  nor2  gate712(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate713(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate714(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate687(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate688(.a(gate104inter0), .b(s_20), .O(gate104inter1));
  and2  gate689(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate690(.a(s_20), .O(gate104inter3));
  inv1  gate691(.a(s_21), .O(gate104inter4));
  nand2 gate692(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate693(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate694(.a(G32), .O(gate104inter7));
  inv1  gate695(.a(G359), .O(gate104inter8));
  nand2 gate696(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate697(.a(s_21), .b(gate104inter3), .O(gate104inter10));
  nor2  gate698(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate699(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate700(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1499(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1500(.a(gate105inter0), .b(s_136), .O(gate105inter1));
  and2  gate1501(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1502(.a(s_136), .O(gate105inter3));
  inv1  gate1503(.a(s_137), .O(gate105inter4));
  nand2 gate1504(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1505(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1506(.a(G362), .O(gate105inter7));
  inv1  gate1507(.a(G363), .O(gate105inter8));
  nand2 gate1508(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1509(.a(s_137), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1510(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1511(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1512(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate729(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate730(.a(gate106inter0), .b(s_26), .O(gate106inter1));
  and2  gate731(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate732(.a(s_26), .O(gate106inter3));
  inv1  gate733(.a(s_27), .O(gate106inter4));
  nand2 gate734(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate735(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate736(.a(G364), .O(gate106inter7));
  inv1  gate737(.a(G365), .O(gate106inter8));
  nand2 gate738(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate739(.a(s_27), .b(gate106inter3), .O(gate106inter10));
  nor2  gate740(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate741(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate742(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1051(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1052(.a(gate107inter0), .b(s_72), .O(gate107inter1));
  and2  gate1053(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1054(.a(s_72), .O(gate107inter3));
  inv1  gate1055(.a(s_73), .O(gate107inter4));
  nand2 gate1056(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1057(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1058(.a(G366), .O(gate107inter7));
  inv1  gate1059(.a(G367), .O(gate107inter8));
  nand2 gate1060(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1061(.a(s_73), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1062(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1063(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1064(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate2045(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2046(.a(gate109inter0), .b(s_214), .O(gate109inter1));
  and2  gate2047(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2048(.a(s_214), .O(gate109inter3));
  inv1  gate2049(.a(s_215), .O(gate109inter4));
  nand2 gate2050(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2051(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2052(.a(G370), .O(gate109inter7));
  inv1  gate2053(.a(G371), .O(gate109inter8));
  nand2 gate2054(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2055(.a(s_215), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2056(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2057(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2058(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1961(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1962(.a(gate112inter0), .b(s_202), .O(gate112inter1));
  and2  gate1963(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1964(.a(s_202), .O(gate112inter3));
  inv1  gate1965(.a(s_203), .O(gate112inter4));
  nand2 gate1966(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1967(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1968(.a(G376), .O(gate112inter7));
  inv1  gate1969(.a(G377), .O(gate112inter8));
  nand2 gate1970(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1971(.a(s_203), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1972(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1973(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1974(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1023(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1024(.a(gate116inter0), .b(s_68), .O(gate116inter1));
  and2  gate1025(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1026(.a(s_68), .O(gate116inter3));
  inv1  gate1027(.a(s_69), .O(gate116inter4));
  nand2 gate1028(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1029(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1030(.a(G384), .O(gate116inter7));
  inv1  gate1031(.a(G385), .O(gate116inter8));
  nand2 gate1032(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1033(.a(s_69), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1034(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1035(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1036(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1919(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1920(.a(gate118inter0), .b(s_196), .O(gate118inter1));
  and2  gate1921(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1922(.a(s_196), .O(gate118inter3));
  inv1  gate1923(.a(s_197), .O(gate118inter4));
  nand2 gate1924(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1925(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1926(.a(G388), .O(gate118inter7));
  inv1  gate1927(.a(G389), .O(gate118inter8));
  nand2 gate1928(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1929(.a(s_197), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1930(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1931(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1932(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1009(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1010(.a(gate121inter0), .b(s_66), .O(gate121inter1));
  and2  gate1011(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1012(.a(s_66), .O(gate121inter3));
  inv1  gate1013(.a(s_67), .O(gate121inter4));
  nand2 gate1014(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1015(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1016(.a(G394), .O(gate121inter7));
  inv1  gate1017(.a(G395), .O(gate121inter8));
  nand2 gate1018(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1019(.a(s_67), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1020(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1021(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1022(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate813(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate814(.a(gate126inter0), .b(s_38), .O(gate126inter1));
  and2  gate815(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate816(.a(s_38), .O(gate126inter3));
  inv1  gate817(.a(s_39), .O(gate126inter4));
  nand2 gate818(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate819(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate820(.a(G404), .O(gate126inter7));
  inv1  gate821(.a(G405), .O(gate126inter8));
  nand2 gate822(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate823(.a(s_39), .b(gate126inter3), .O(gate126inter10));
  nor2  gate824(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate825(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate826(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate659(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate660(.a(gate134inter0), .b(s_16), .O(gate134inter1));
  and2  gate661(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate662(.a(s_16), .O(gate134inter3));
  inv1  gate663(.a(s_17), .O(gate134inter4));
  nand2 gate664(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate665(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate666(.a(G420), .O(gate134inter7));
  inv1  gate667(.a(G421), .O(gate134inter8));
  nand2 gate668(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate669(.a(s_17), .b(gate134inter3), .O(gate134inter10));
  nor2  gate670(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate671(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate672(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1149(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1150(.a(gate140inter0), .b(s_86), .O(gate140inter1));
  and2  gate1151(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1152(.a(s_86), .O(gate140inter3));
  inv1  gate1153(.a(s_87), .O(gate140inter4));
  nand2 gate1154(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1155(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1156(.a(G444), .O(gate140inter7));
  inv1  gate1157(.a(G447), .O(gate140inter8));
  nand2 gate1158(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1159(.a(s_87), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1160(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1161(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1162(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1947(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1948(.a(gate141inter0), .b(s_200), .O(gate141inter1));
  and2  gate1949(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1950(.a(s_200), .O(gate141inter3));
  inv1  gate1951(.a(s_201), .O(gate141inter4));
  nand2 gate1952(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1953(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1954(.a(G450), .O(gate141inter7));
  inv1  gate1955(.a(G453), .O(gate141inter8));
  nand2 gate1956(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1957(.a(s_201), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1958(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1959(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1960(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1597(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1598(.a(gate146inter0), .b(s_150), .O(gate146inter1));
  and2  gate1599(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1600(.a(s_150), .O(gate146inter3));
  inv1  gate1601(.a(s_151), .O(gate146inter4));
  nand2 gate1602(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1603(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1604(.a(G480), .O(gate146inter7));
  inv1  gate1605(.a(G483), .O(gate146inter8));
  nand2 gate1606(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1607(.a(s_151), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1608(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1609(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1610(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1807(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1808(.a(gate147inter0), .b(s_180), .O(gate147inter1));
  and2  gate1809(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1810(.a(s_180), .O(gate147inter3));
  inv1  gate1811(.a(s_181), .O(gate147inter4));
  nand2 gate1812(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1813(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1814(.a(G486), .O(gate147inter7));
  inv1  gate1815(.a(G489), .O(gate147inter8));
  nand2 gate1816(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1817(.a(s_181), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1818(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1819(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1820(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate883(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate884(.a(gate149inter0), .b(s_48), .O(gate149inter1));
  and2  gate885(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate886(.a(s_48), .O(gate149inter3));
  inv1  gate887(.a(s_49), .O(gate149inter4));
  nand2 gate888(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate889(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate890(.a(G498), .O(gate149inter7));
  inv1  gate891(.a(G501), .O(gate149inter8));
  nand2 gate892(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate893(.a(s_49), .b(gate149inter3), .O(gate149inter10));
  nor2  gate894(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate895(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate896(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate827(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate828(.a(gate153inter0), .b(s_40), .O(gate153inter1));
  and2  gate829(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate830(.a(s_40), .O(gate153inter3));
  inv1  gate831(.a(s_41), .O(gate153inter4));
  nand2 gate832(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate833(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate834(.a(G426), .O(gate153inter7));
  inv1  gate835(.a(G522), .O(gate153inter8));
  nand2 gate836(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate837(.a(s_41), .b(gate153inter3), .O(gate153inter10));
  nor2  gate838(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate839(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate840(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate575(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate576(.a(gate155inter0), .b(s_4), .O(gate155inter1));
  and2  gate577(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate578(.a(s_4), .O(gate155inter3));
  inv1  gate579(.a(s_5), .O(gate155inter4));
  nand2 gate580(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate581(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate582(.a(G432), .O(gate155inter7));
  inv1  gate583(.a(G525), .O(gate155inter8));
  nand2 gate584(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate585(.a(s_5), .b(gate155inter3), .O(gate155inter10));
  nor2  gate586(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate587(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate588(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1401(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1402(.a(gate158inter0), .b(s_122), .O(gate158inter1));
  and2  gate1403(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1404(.a(s_122), .O(gate158inter3));
  inv1  gate1405(.a(s_123), .O(gate158inter4));
  nand2 gate1406(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1407(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1408(.a(G441), .O(gate158inter7));
  inv1  gate1409(.a(G528), .O(gate158inter8));
  nand2 gate1410(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1411(.a(s_123), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1412(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1413(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1414(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1625(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1626(.a(gate159inter0), .b(s_154), .O(gate159inter1));
  and2  gate1627(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1628(.a(s_154), .O(gate159inter3));
  inv1  gate1629(.a(s_155), .O(gate159inter4));
  nand2 gate1630(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1631(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1632(.a(G444), .O(gate159inter7));
  inv1  gate1633(.a(G531), .O(gate159inter8));
  nand2 gate1634(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1635(.a(s_155), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1636(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1637(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1638(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate939(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate940(.a(gate165inter0), .b(s_56), .O(gate165inter1));
  and2  gate941(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate942(.a(s_56), .O(gate165inter3));
  inv1  gate943(.a(s_57), .O(gate165inter4));
  nand2 gate944(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate945(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate946(.a(G462), .O(gate165inter7));
  inv1  gate947(.a(G540), .O(gate165inter8));
  nand2 gate948(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate949(.a(s_57), .b(gate165inter3), .O(gate165inter10));
  nor2  gate950(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate951(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate952(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1863(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1864(.a(gate168inter0), .b(s_188), .O(gate168inter1));
  and2  gate1865(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1866(.a(s_188), .O(gate168inter3));
  inv1  gate1867(.a(s_189), .O(gate168inter4));
  nand2 gate1868(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1869(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1870(.a(G471), .O(gate168inter7));
  inv1  gate1871(.a(G543), .O(gate168inter8));
  nand2 gate1872(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1873(.a(s_189), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1874(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1875(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1876(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate869(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate870(.a(gate172inter0), .b(s_46), .O(gate172inter1));
  and2  gate871(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate872(.a(s_46), .O(gate172inter3));
  inv1  gate873(.a(s_47), .O(gate172inter4));
  nand2 gate874(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate875(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate876(.a(G483), .O(gate172inter7));
  inv1  gate877(.a(G549), .O(gate172inter8));
  nand2 gate878(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate879(.a(s_47), .b(gate172inter3), .O(gate172inter10));
  nor2  gate880(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate881(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate882(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate2087(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2088(.a(gate177inter0), .b(s_220), .O(gate177inter1));
  and2  gate2089(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2090(.a(s_220), .O(gate177inter3));
  inv1  gate2091(.a(s_221), .O(gate177inter4));
  nand2 gate2092(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2093(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2094(.a(G498), .O(gate177inter7));
  inv1  gate2095(.a(G558), .O(gate177inter8));
  nand2 gate2096(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2097(.a(s_221), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2098(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2099(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2100(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1541(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1542(.a(gate183inter0), .b(s_142), .O(gate183inter1));
  and2  gate1543(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1544(.a(s_142), .O(gate183inter3));
  inv1  gate1545(.a(s_143), .O(gate183inter4));
  nand2 gate1546(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1547(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1548(.a(G516), .O(gate183inter7));
  inv1  gate1549(.a(G567), .O(gate183inter8));
  nand2 gate1550(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1551(.a(s_143), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1552(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1553(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1554(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1737(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1738(.a(gate187inter0), .b(s_170), .O(gate187inter1));
  and2  gate1739(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1740(.a(s_170), .O(gate187inter3));
  inv1  gate1741(.a(s_171), .O(gate187inter4));
  nand2 gate1742(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1743(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1744(.a(G574), .O(gate187inter7));
  inv1  gate1745(.a(G575), .O(gate187inter8));
  nand2 gate1746(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1747(.a(s_171), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1748(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1749(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1750(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2059(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2060(.a(gate188inter0), .b(s_216), .O(gate188inter1));
  and2  gate2061(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2062(.a(s_216), .O(gate188inter3));
  inv1  gate2063(.a(s_217), .O(gate188inter4));
  nand2 gate2064(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2065(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2066(.a(G576), .O(gate188inter7));
  inv1  gate2067(.a(G577), .O(gate188inter8));
  nand2 gate2068(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2069(.a(s_217), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2070(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2071(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2072(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate995(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate996(.a(gate190inter0), .b(s_64), .O(gate190inter1));
  and2  gate997(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate998(.a(s_64), .O(gate190inter3));
  inv1  gate999(.a(s_65), .O(gate190inter4));
  nand2 gate1000(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1001(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1002(.a(G580), .O(gate190inter7));
  inv1  gate1003(.a(G581), .O(gate190inter8));
  nand2 gate1004(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1005(.a(s_65), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1006(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1007(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1008(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate841(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate842(.a(gate191inter0), .b(s_42), .O(gate191inter1));
  and2  gate843(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate844(.a(s_42), .O(gate191inter3));
  inv1  gate845(.a(s_43), .O(gate191inter4));
  nand2 gate846(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate847(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate848(.a(G582), .O(gate191inter7));
  inv1  gate849(.a(G583), .O(gate191inter8));
  nand2 gate850(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate851(.a(s_43), .b(gate191inter3), .O(gate191inter10));
  nor2  gate852(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate853(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate854(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate715(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate716(.a(gate194inter0), .b(s_24), .O(gate194inter1));
  and2  gate717(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate718(.a(s_24), .O(gate194inter3));
  inv1  gate719(.a(s_25), .O(gate194inter4));
  nand2 gate720(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate721(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate722(.a(G588), .O(gate194inter7));
  inv1  gate723(.a(G589), .O(gate194inter8));
  nand2 gate724(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate725(.a(s_25), .b(gate194inter3), .O(gate194inter10));
  nor2  gate726(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate727(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate728(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1527(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1528(.a(gate197inter0), .b(s_140), .O(gate197inter1));
  and2  gate1529(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1530(.a(s_140), .O(gate197inter3));
  inv1  gate1531(.a(s_141), .O(gate197inter4));
  nand2 gate1532(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1533(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1534(.a(G594), .O(gate197inter7));
  inv1  gate1535(.a(G595), .O(gate197inter8));
  nand2 gate1536(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1537(.a(s_141), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1538(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1539(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1540(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1345(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1346(.a(gate199inter0), .b(s_114), .O(gate199inter1));
  and2  gate1347(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1348(.a(s_114), .O(gate199inter3));
  inv1  gate1349(.a(s_115), .O(gate199inter4));
  nand2 gate1350(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1351(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1352(.a(G598), .O(gate199inter7));
  inv1  gate1353(.a(G599), .O(gate199inter8));
  nand2 gate1354(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1355(.a(s_115), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1356(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1357(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1358(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1933(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1934(.a(gate202inter0), .b(s_198), .O(gate202inter1));
  and2  gate1935(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1936(.a(s_198), .O(gate202inter3));
  inv1  gate1937(.a(s_199), .O(gate202inter4));
  nand2 gate1938(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1939(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1940(.a(G612), .O(gate202inter7));
  inv1  gate1941(.a(G617), .O(gate202inter8));
  nand2 gate1942(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1943(.a(s_199), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1944(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1945(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1946(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate757(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate758(.a(gate205inter0), .b(s_30), .O(gate205inter1));
  and2  gate759(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate760(.a(s_30), .O(gate205inter3));
  inv1  gate761(.a(s_31), .O(gate205inter4));
  nand2 gate762(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate763(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate764(.a(G622), .O(gate205inter7));
  inv1  gate765(.a(G627), .O(gate205inter8));
  nand2 gate766(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate767(.a(s_31), .b(gate205inter3), .O(gate205inter10));
  nor2  gate768(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate769(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate770(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1471(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1472(.a(gate209inter0), .b(s_132), .O(gate209inter1));
  and2  gate1473(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1474(.a(s_132), .O(gate209inter3));
  inv1  gate1475(.a(s_133), .O(gate209inter4));
  nand2 gate1476(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1477(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1478(.a(G602), .O(gate209inter7));
  inv1  gate1479(.a(G666), .O(gate209inter8));
  nand2 gate1480(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1481(.a(s_133), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1482(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1483(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1484(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1163(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1164(.a(gate211inter0), .b(s_88), .O(gate211inter1));
  and2  gate1165(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1166(.a(s_88), .O(gate211inter3));
  inv1  gate1167(.a(s_89), .O(gate211inter4));
  nand2 gate1168(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1169(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1170(.a(G612), .O(gate211inter7));
  inv1  gate1171(.a(G669), .O(gate211inter8));
  nand2 gate1172(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1173(.a(s_89), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1174(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1175(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1176(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2031(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2032(.a(gate212inter0), .b(s_212), .O(gate212inter1));
  and2  gate2033(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2034(.a(s_212), .O(gate212inter3));
  inv1  gate2035(.a(s_213), .O(gate212inter4));
  nand2 gate2036(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2037(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2038(.a(G617), .O(gate212inter7));
  inv1  gate2039(.a(G669), .O(gate212inter8));
  nand2 gate2040(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2041(.a(s_213), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2042(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2043(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2044(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1849(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1850(.a(gate214inter0), .b(s_186), .O(gate214inter1));
  and2  gate1851(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1852(.a(s_186), .O(gate214inter3));
  inv1  gate1853(.a(s_187), .O(gate214inter4));
  nand2 gate1854(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1855(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1856(.a(G612), .O(gate214inter7));
  inv1  gate1857(.a(G672), .O(gate214inter8));
  nand2 gate1858(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1859(.a(s_187), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1860(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1861(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1862(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1331(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1332(.a(gate219inter0), .b(s_112), .O(gate219inter1));
  and2  gate1333(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1334(.a(s_112), .O(gate219inter3));
  inv1  gate1335(.a(s_113), .O(gate219inter4));
  nand2 gate1336(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1337(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1338(.a(G632), .O(gate219inter7));
  inv1  gate1339(.a(G681), .O(gate219inter8));
  nand2 gate1340(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1341(.a(s_113), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1342(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1343(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1344(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1205(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1206(.a(gate221inter0), .b(s_94), .O(gate221inter1));
  and2  gate1207(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1208(.a(s_94), .O(gate221inter3));
  inv1  gate1209(.a(s_95), .O(gate221inter4));
  nand2 gate1210(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1211(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1212(.a(G622), .O(gate221inter7));
  inv1  gate1213(.a(G684), .O(gate221inter8));
  nand2 gate1214(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1215(.a(s_95), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1216(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1217(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1218(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1275(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1276(.a(gate222inter0), .b(s_104), .O(gate222inter1));
  and2  gate1277(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1278(.a(s_104), .O(gate222inter3));
  inv1  gate1279(.a(s_105), .O(gate222inter4));
  nand2 gate1280(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1281(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1282(.a(G632), .O(gate222inter7));
  inv1  gate1283(.a(G684), .O(gate222inter8));
  nand2 gate1284(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1285(.a(s_105), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1286(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1287(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1288(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate673(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate674(.a(gate224inter0), .b(s_18), .O(gate224inter1));
  and2  gate675(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate676(.a(s_18), .O(gate224inter3));
  inv1  gate677(.a(s_19), .O(gate224inter4));
  nand2 gate678(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate679(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate680(.a(G637), .O(gate224inter7));
  inv1  gate681(.a(G687), .O(gate224inter8));
  nand2 gate682(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate683(.a(s_19), .b(gate224inter3), .O(gate224inter10));
  nor2  gate684(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate685(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate686(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1289(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1290(.a(gate233inter0), .b(s_106), .O(gate233inter1));
  and2  gate1291(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1292(.a(s_106), .O(gate233inter3));
  inv1  gate1293(.a(s_107), .O(gate233inter4));
  nand2 gate1294(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1295(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1296(.a(G242), .O(gate233inter7));
  inv1  gate1297(.a(G718), .O(gate233inter8));
  nand2 gate1298(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1299(.a(s_107), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1300(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1301(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1302(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1555(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1556(.a(gate236inter0), .b(s_144), .O(gate236inter1));
  and2  gate1557(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1558(.a(s_144), .O(gate236inter3));
  inv1  gate1559(.a(s_145), .O(gate236inter4));
  nand2 gate1560(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1561(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1562(.a(G251), .O(gate236inter7));
  inv1  gate1563(.a(G727), .O(gate236inter8));
  nand2 gate1564(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1565(.a(s_145), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1566(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1567(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1568(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate771(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate772(.a(gate237inter0), .b(s_32), .O(gate237inter1));
  and2  gate773(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate774(.a(s_32), .O(gate237inter3));
  inv1  gate775(.a(s_33), .O(gate237inter4));
  nand2 gate776(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate777(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate778(.a(G254), .O(gate237inter7));
  inv1  gate779(.a(G706), .O(gate237inter8));
  nand2 gate780(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate781(.a(s_33), .b(gate237inter3), .O(gate237inter10));
  nor2  gate782(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate783(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate784(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate785(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate786(.a(gate245inter0), .b(s_34), .O(gate245inter1));
  and2  gate787(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate788(.a(s_34), .O(gate245inter3));
  inv1  gate789(.a(s_35), .O(gate245inter4));
  nand2 gate790(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate791(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate792(.a(G248), .O(gate245inter7));
  inv1  gate793(.a(G736), .O(gate245inter8));
  nand2 gate794(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate795(.a(s_35), .b(gate245inter3), .O(gate245inter10));
  nor2  gate796(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate797(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate798(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1107(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1108(.a(gate247inter0), .b(s_80), .O(gate247inter1));
  and2  gate1109(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1110(.a(s_80), .O(gate247inter3));
  inv1  gate1111(.a(s_81), .O(gate247inter4));
  nand2 gate1112(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1113(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1114(.a(G251), .O(gate247inter7));
  inv1  gate1115(.a(G739), .O(gate247inter8));
  nand2 gate1116(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1117(.a(s_81), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1118(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1119(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1120(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1639(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1640(.a(gate249inter0), .b(s_156), .O(gate249inter1));
  and2  gate1641(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1642(.a(s_156), .O(gate249inter3));
  inv1  gate1643(.a(s_157), .O(gate249inter4));
  nand2 gate1644(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1645(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1646(.a(G254), .O(gate249inter7));
  inv1  gate1647(.a(G742), .O(gate249inter8));
  nand2 gate1648(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1649(.a(s_157), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1650(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1651(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1652(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1779(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1780(.a(gate253inter0), .b(s_176), .O(gate253inter1));
  and2  gate1781(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1782(.a(s_176), .O(gate253inter3));
  inv1  gate1783(.a(s_177), .O(gate253inter4));
  nand2 gate1784(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1785(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1786(.a(G260), .O(gate253inter7));
  inv1  gate1787(.a(G748), .O(gate253inter8));
  nand2 gate1788(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1789(.a(s_177), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1790(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1791(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1792(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate645(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate646(.a(gate256inter0), .b(s_14), .O(gate256inter1));
  and2  gate647(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate648(.a(s_14), .O(gate256inter3));
  inv1  gate649(.a(s_15), .O(gate256inter4));
  nand2 gate650(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate651(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate652(.a(G715), .O(gate256inter7));
  inv1  gate653(.a(G751), .O(gate256inter8));
  nand2 gate654(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate655(.a(s_15), .b(gate256inter3), .O(gate256inter10));
  nor2  gate656(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate657(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate658(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1317(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1318(.a(gate262inter0), .b(s_110), .O(gate262inter1));
  and2  gate1319(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1320(.a(s_110), .O(gate262inter3));
  inv1  gate1321(.a(s_111), .O(gate262inter4));
  nand2 gate1322(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1323(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1324(.a(G764), .O(gate262inter7));
  inv1  gate1325(.a(G765), .O(gate262inter8));
  nand2 gate1326(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1327(.a(s_111), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1328(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1329(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1330(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate2003(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2004(.a(gate266inter0), .b(s_208), .O(gate266inter1));
  and2  gate2005(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2006(.a(s_208), .O(gate266inter3));
  inv1  gate2007(.a(s_209), .O(gate266inter4));
  nand2 gate2008(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2009(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2010(.a(G645), .O(gate266inter7));
  inv1  gate2011(.a(G773), .O(gate266inter8));
  nand2 gate2012(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2013(.a(s_209), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2014(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2015(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2016(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate981(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate982(.a(gate277inter0), .b(s_62), .O(gate277inter1));
  and2  gate983(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate984(.a(s_62), .O(gate277inter3));
  inv1  gate985(.a(s_63), .O(gate277inter4));
  nand2 gate986(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate987(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate988(.a(G648), .O(gate277inter7));
  inv1  gate989(.a(G800), .O(gate277inter8));
  nand2 gate990(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate991(.a(s_63), .b(gate277inter3), .O(gate277inter10));
  nor2  gate992(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate993(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate994(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1569(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1570(.a(gate290inter0), .b(s_146), .O(gate290inter1));
  and2  gate1571(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1572(.a(s_146), .O(gate290inter3));
  inv1  gate1573(.a(s_147), .O(gate290inter4));
  nand2 gate1574(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1575(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1576(.a(G820), .O(gate290inter7));
  inv1  gate1577(.a(G821), .O(gate290inter8));
  nand2 gate1578(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1579(.a(s_147), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1580(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1581(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1582(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1765(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1766(.a(gate294inter0), .b(s_174), .O(gate294inter1));
  and2  gate1767(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1768(.a(s_174), .O(gate294inter3));
  inv1  gate1769(.a(s_175), .O(gate294inter4));
  nand2 gate1770(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1771(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1772(.a(G832), .O(gate294inter7));
  inv1  gate1773(.a(G833), .O(gate294inter8));
  nand2 gate1774(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1775(.a(s_175), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1776(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1777(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1778(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2073(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2074(.a(gate393inter0), .b(s_218), .O(gate393inter1));
  and2  gate2075(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2076(.a(s_218), .O(gate393inter3));
  inv1  gate2077(.a(s_219), .O(gate393inter4));
  nand2 gate2078(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2079(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2080(.a(G7), .O(gate393inter7));
  inv1  gate2081(.a(G1054), .O(gate393inter8));
  nand2 gate2082(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2083(.a(s_219), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2084(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2085(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2086(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1191(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1192(.a(gate396inter0), .b(s_92), .O(gate396inter1));
  and2  gate1193(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1194(.a(s_92), .O(gate396inter3));
  inv1  gate1195(.a(s_93), .O(gate396inter4));
  nand2 gate1196(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1197(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1198(.a(G10), .O(gate396inter7));
  inv1  gate1199(.a(G1063), .O(gate396inter8));
  nand2 gate1200(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1201(.a(s_93), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1202(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1203(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1204(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1835(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1836(.a(gate397inter0), .b(s_184), .O(gate397inter1));
  and2  gate1837(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1838(.a(s_184), .O(gate397inter3));
  inv1  gate1839(.a(s_185), .O(gate397inter4));
  nand2 gate1840(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1841(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1842(.a(G11), .O(gate397inter7));
  inv1  gate1843(.a(G1066), .O(gate397inter8));
  nand2 gate1844(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1845(.a(s_185), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1846(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1847(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1848(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1387(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1388(.a(gate399inter0), .b(s_120), .O(gate399inter1));
  and2  gate1389(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1390(.a(s_120), .O(gate399inter3));
  inv1  gate1391(.a(s_121), .O(gate399inter4));
  nand2 gate1392(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1393(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1394(.a(G13), .O(gate399inter7));
  inv1  gate1395(.a(G1072), .O(gate399inter8));
  nand2 gate1396(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1397(.a(s_121), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1398(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1399(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1400(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate617(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate618(.a(gate400inter0), .b(s_10), .O(gate400inter1));
  and2  gate619(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate620(.a(s_10), .O(gate400inter3));
  inv1  gate621(.a(s_11), .O(gate400inter4));
  nand2 gate622(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate623(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate624(.a(G14), .O(gate400inter7));
  inv1  gate625(.a(G1075), .O(gate400inter8));
  nand2 gate626(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate627(.a(s_11), .b(gate400inter3), .O(gate400inter10));
  nor2  gate628(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate629(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate630(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1457(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1458(.a(gate401inter0), .b(s_130), .O(gate401inter1));
  and2  gate1459(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1460(.a(s_130), .O(gate401inter3));
  inv1  gate1461(.a(s_131), .O(gate401inter4));
  nand2 gate1462(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1463(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1464(.a(G15), .O(gate401inter7));
  inv1  gate1465(.a(G1078), .O(gate401inter8));
  nand2 gate1466(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1467(.a(s_131), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1468(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1469(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1470(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1667(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1668(.a(gate403inter0), .b(s_160), .O(gate403inter1));
  and2  gate1669(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1670(.a(s_160), .O(gate403inter3));
  inv1  gate1671(.a(s_161), .O(gate403inter4));
  nand2 gate1672(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1673(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1674(.a(G17), .O(gate403inter7));
  inv1  gate1675(.a(G1084), .O(gate403inter8));
  nand2 gate1676(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1677(.a(s_161), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1678(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1679(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1680(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1793(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1794(.a(gate407inter0), .b(s_178), .O(gate407inter1));
  and2  gate1795(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1796(.a(s_178), .O(gate407inter3));
  inv1  gate1797(.a(s_179), .O(gate407inter4));
  nand2 gate1798(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1799(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1800(.a(G21), .O(gate407inter7));
  inv1  gate1801(.a(G1096), .O(gate407inter8));
  nand2 gate1802(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1803(.a(s_179), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1804(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1805(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1806(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1247(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1248(.a(gate409inter0), .b(s_100), .O(gate409inter1));
  and2  gate1249(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1250(.a(s_100), .O(gate409inter3));
  inv1  gate1251(.a(s_101), .O(gate409inter4));
  nand2 gate1252(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1253(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1254(.a(G23), .O(gate409inter7));
  inv1  gate1255(.a(G1102), .O(gate409inter8));
  nand2 gate1256(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1257(.a(s_101), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1258(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1259(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1260(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1975(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1976(.a(gate411inter0), .b(s_204), .O(gate411inter1));
  and2  gate1977(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1978(.a(s_204), .O(gate411inter3));
  inv1  gate1979(.a(s_205), .O(gate411inter4));
  nand2 gate1980(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1981(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1982(.a(G25), .O(gate411inter7));
  inv1  gate1983(.a(G1108), .O(gate411inter8));
  nand2 gate1984(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1985(.a(s_205), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1986(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1987(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1988(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1359(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1360(.a(gate413inter0), .b(s_116), .O(gate413inter1));
  and2  gate1361(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1362(.a(s_116), .O(gate413inter3));
  inv1  gate1363(.a(s_117), .O(gate413inter4));
  nand2 gate1364(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1365(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1366(.a(G27), .O(gate413inter7));
  inv1  gate1367(.a(G1114), .O(gate413inter8));
  nand2 gate1368(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1369(.a(s_117), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1370(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1371(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1372(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate603(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate604(.a(gate417inter0), .b(s_8), .O(gate417inter1));
  and2  gate605(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate606(.a(s_8), .O(gate417inter3));
  inv1  gate607(.a(s_9), .O(gate417inter4));
  nand2 gate608(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate609(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate610(.a(G31), .O(gate417inter7));
  inv1  gate611(.a(G1126), .O(gate417inter8));
  nand2 gate612(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate613(.a(s_9), .b(gate417inter3), .O(gate417inter10));
  nor2  gate614(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate615(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate616(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1821(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1822(.a(gate422inter0), .b(s_182), .O(gate422inter1));
  and2  gate1823(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1824(.a(s_182), .O(gate422inter3));
  inv1  gate1825(.a(s_183), .O(gate422inter4));
  nand2 gate1826(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1827(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1828(.a(G1039), .O(gate422inter7));
  inv1  gate1829(.a(G1135), .O(gate422inter8));
  nand2 gate1830(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1831(.a(s_183), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1832(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1833(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1834(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1891(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1892(.a(gate424inter0), .b(s_192), .O(gate424inter1));
  and2  gate1893(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1894(.a(s_192), .O(gate424inter3));
  inv1  gate1895(.a(s_193), .O(gate424inter4));
  nand2 gate1896(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1897(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1898(.a(G1042), .O(gate424inter7));
  inv1  gate1899(.a(G1138), .O(gate424inter8));
  nand2 gate1900(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1901(.a(s_193), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1902(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1903(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1904(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1079(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1080(.a(gate425inter0), .b(s_76), .O(gate425inter1));
  and2  gate1081(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1082(.a(s_76), .O(gate425inter3));
  inv1  gate1083(.a(s_77), .O(gate425inter4));
  nand2 gate1084(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1085(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1086(.a(G4), .O(gate425inter7));
  inv1  gate1087(.a(G1141), .O(gate425inter8));
  nand2 gate1088(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1089(.a(s_77), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1090(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1091(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1092(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1513(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1514(.a(gate429inter0), .b(s_138), .O(gate429inter1));
  and2  gate1515(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1516(.a(s_138), .O(gate429inter3));
  inv1  gate1517(.a(s_139), .O(gate429inter4));
  nand2 gate1518(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1519(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1520(.a(G6), .O(gate429inter7));
  inv1  gate1521(.a(G1147), .O(gate429inter8));
  nand2 gate1522(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1523(.a(s_139), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1524(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1525(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1526(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate631(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate632(.a(gate431inter0), .b(s_12), .O(gate431inter1));
  and2  gate633(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate634(.a(s_12), .O(gate431inter3));
  inv1  gate635(.a(s_13), .O(gate431inter4));
  nand2 gate636(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate637(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate638(.a(G7), .O(gate431inter7));
  inv1  gate639(.a(G1150), .O(gate431inter8));
  nand2 gate640(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate641(.a(s_13), .b(gate431inter3), .O(gate431inter10));
  nor2  gate642(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate643(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate644(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1905(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1906(.a(gate437inter0), .b(s_194), .O(gate437inter1));
  and2  gate1907(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1908(.a(s_194), .O(gate437inter3));
  inv1  gate1909(.a(s_195), .O(gate437inter4));
  nand2 gate1910(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1911(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1912(.a(G10), .O(gate437inter7));
  inv1  gate1913(.a(G1159), .O(gate437inter8));
  nand2 gate1914(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1915(.a(s_195), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1916(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1917(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1918(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1415(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1416(.a(gate446inter0), .b(s_124), .O(gate446inter1));
  and2  gate1417(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1418(.a(s_124), .O(gate446inter3));
  inv1  gate1419(.a(s_125), .O(gate446inter4));
  nand2 gate1420(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1421(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1422(.a(G1075), .O(gate446inter7));
  inv1  gate1423(.a(G1171), .O(gate446inter8));
  nand2 gate1424(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1425(.a(s_125), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1426(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1427(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1428(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate799(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate800(.a(gate456inter0), .b(s_36), .O(gate456inter1));
  and2  gate801(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate802(.a(s_36), .O(gate456inter3));
  inv1  gate803(.a(s_37), .O(gate456inter4));
  nand2 gate804(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate805(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate806(.a(G1090), .O(gate456inter7));
  inv1  gate807(.a(G1186), .O(gate456inter8));
  nand2 gate808(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate809(.a(s_37), .b(gate456inter3), .O(gate456inter10));
  nor2  gate810(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate811(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate812(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1751(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1752(.a(gate458inter0), .b(s_172), .O(gate458inter1));
  and2  gate1753(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1754(.a(s_172), .O(gate458inter3));
  inv1  gate1755(.a(s_173), .O(gate458inter4));
  nand2 gate1756(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1757(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1758(.a(G1093), .O(gate458inter7));
  inv1  gate1759(.a(G1189), .O(gate458inter8));
  nand2 gate1760(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1761(.a(s_173), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1762(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1763(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1764(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1583(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1584(.a(gate459inter0), .b(s_148), .O(gate459inter1));
  and2  gate1585(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1586(.a(s_148), .O(gate459inter3));
  inv1  gate1587(.a(s_149), .O(gate459inter4));
  nand2 gate1588(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1589(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1590(.a(G21), .O(gate459inter7));
  inv1  gate1591(.a(G1192), .O(gate459inter8));
  nand2 gate1592(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1593(.a(s_149), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1594(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1595(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1596(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1709(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1710(.a(gate466inter0), .b(s_166), .O(gate466inter1));
  and2  gate1711(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1712(.a(s_166), .O(gate466inter3));
  inv1  gate1713(.a(s_167), .O(gate466inter4));
  nand2 gate1714(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1715(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1716(.a(G1105), .O(gate466inter7));
  inv1  gate1717(.a(G1201), .O(gate466inter8));
  nand2 gate1718(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1719(.a(s_167), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1720(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1721(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1722(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1611(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1612(.a(gate470inter0), .b(s_152), .O(gate470inter1));
  and2  gate1613(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1614(.a(s_152), .O(gate470inter3));
  inv1  gate1615(.a(s_153), .O(gate470inter4));
  nand2 gate1616(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1617(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1618(.a(G1111), .O(gate470inter7));
  inv1  gate1619(.a(G1207), .O(gate470inter8));
  nand2 gate1620(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1621(.a(s_153), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1622(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1623(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1624(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate925(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate926(.a(gate474inter0), .b(s_54), .O(gate474inter1));
  and2  gate927(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate928(.a(s_54), .O(gate474inter3));
  inv1  gate929(.a(s_55), .O(gate474inter4));
  nand2 gate930(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate931(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate932(.a(G1117), .O(gate474inter7));
  inv1  gate933(.a(G1213), .O(gate474inter8));
  nand2 gate934(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate935(.a(s_55), .b(gate474inter3), .O(gate474inter10));
  nor2  gate936(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate937(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate938(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate953(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate954(.a(gate475inter0), .b(s_58), .O(gate475inter1));
  and2  gate955(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate956(.a(s_58), .O(gate475inter3));
  inv1  gate957(.a(s_59), .O(gate475inter4));
  nand2 gate958(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate959(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate960(.a(G29), .O(gate475inter7));
  inv1  gate961(.a(G1216), .O(gate475inter8));
  nand2 gate962(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate963(.a(s_59), .b(gate475inter3), .O(gate475inter10));
  nor2  gate964(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate965(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate966(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1233(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1234(.a(gate477inter0), .b(s_98), .O(gate477inter1));
  and2  gate1235(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1236(.a(s_98), .O(gate477inter3));
  inv1  gate1237(.a(s_99), .O(gate477inter4));
  nand2 gate1238(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1239(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1240(.a(G30), .O(gate477inter7));
  inv1  gate1241(.a(G1219), .O(gate477inter8));
  nand2 gate1242(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1243(.a(s_99), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1244(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1245(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1246(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1429(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1430(.a(gate479inter0), .b(s_126), .O(gate479inter1));
  and2  gate1431(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1432(.a(s_126), .O(gate479inter3));
  inv1  gate1433(.a(s_127), .O(gate479inter4));
  nand2 gate1434(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1435(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1436(.a(G31), .O(gate479inter7));
  inv1  gate1437(.a(G1222), .O(gate479inter8));
  nand2 gate1438(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1439(.a(s_127), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1440(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1441(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1442(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate589(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate590(.a(gate480inter0), .b(s_6), .O(gate480inter1));
  and2  gate591(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate592(.a(s_6), .O(gate480inter3));
  inv1  gate593(.a(s_7), .O(gate480inter4));
  nand2 gate594(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate595(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate596(.a(G1126), .O(gate480inter7));
  inv1  gate597(.a(G1222), .O(gate480inter8));
  nand2 gate598(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate599(.a(s_7), .b(gate480inter3), .O(gate480inter10));
  nor2  gate600(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate601(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate602(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate855(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate856(.a(gate488inter0), .b(s_44), .O(gate488inter1));
  and2  gate857(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate858(.a(s_44), .O(gate488inter3));
  inv1  gate859(.a(s_45), .O(gate488inter4));
  nand2 gate860(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate861(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate862(.a(G1238), .O(gate488inter7));
  inv1  gate863(.a(G1239), .O(gate488inter8));
  nand2 gate864(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate865(.a(s_45), .b(gate488inter3), .O(gate488inter10));
  nor2  gate866(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate867(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate868(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate2017(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2018(.a(gate489inter0), .b(s_210), .O(gate489inter1));
  and2  gate2019(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2020(.a(s_210), .O(gate489inter3));
  inv1  gate2021(.a(s_211), .O(gate489inter4));
  nand2 gate2022(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2023(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2024(.a(G1240), .O(gate489inter7));
  inv1  gate2025(.a(G1241), .O(gate489inter8));
  nand2 gate2026(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2027(.a(s_211), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2028(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2029(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2030(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1989(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1990(.a(gate492inter0), .b(s_206), .O(gate492inter1));
  and2  gate1991(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1992(.a(s_206), .O(gate492inter3));
  inv1  gate1993(.a(s_207), .O(gate492inter4));
  nand2 gate1994(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1995(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1996(.a(G1246), .O(gate492inter7));
  inv1  gate1997(.a(G1247), .O(gate492inter8));
  nand2 gate1998(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1999(.a(s_207), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2000(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2001(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2002(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1877(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1878(.a(gate495inter0), .b(s_190), .O(gate495inter1));
  and2  gate1879(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1880(.a(s_190), .O(gate495inter3));
  inv1  gate1881(.a(s_191), .O(gate495inter4));
  nand2 gate1882(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1883(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1884(.a(G1252), .O(gate495inter7));
  inv1  gate1885(.a(G1253), .O(gate495inter8));
  nand2 gate1886(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1887(.a(s_191), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1888(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1889(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1890(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate561(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate562(.a(gate506inter0), .b(s_2), .O(gate506inter1));
  and2  gate563(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate564(.a(s_2), .O(gate506inter3));
  inv1  gate565(.a(s_3), .O(gate506inter4));
  nand2 gate566(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate567(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate568(.a(G1274), .O(gate506inter7));
  inv1  gate569(.a(G1275), .O(gate506inter8));
  nand2 gate570(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate571(.a(s_3), .b(gate506inter3), .O(gate506inter10));
  nor2  gate572(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate573(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate574(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule