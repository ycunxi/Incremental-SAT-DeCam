module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1051(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1052(.a(gate12inter0), .b(s_72), .O(gate12inter1));
  and2  gate1053(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1054(.a(s_72), .O(gate12inter3));
  inv1  gate1055(.a(s_73), .O(gate12inter4));
  nand2 gate1056(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1057(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1058(.a(G7), .O(gate12inter7));
  inv1  gate1059(.a(G8), .O(gate12inter8));
  nand2 gate1060(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1061(.a(s_73), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1062(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1063(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1064(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate925(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate926(.a(gate13inter0), .b(s_54), .O(gate13inter1));
  and2  gate927(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate928(.a(s_54), .O(gate13inter3));
  inv1  gate929(.a(s_55), .O(gate13inter4));
  nand2 gate930(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate931(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate932(.a(G9), .O(gate13inter7));
  inv1  gate933(.a(G10), .O(gate13inter8));
  nand2 gate934(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate935(.a(s_55), .b(gate13inter3), .O(gate13inter10));
  nor2  gate936(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate937(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate938(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1401(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1402(.a(gate14inter0), .b(s_122), .O(gate14inter1));
  and2  gate1403(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1404(.a(s_122), .O(gate14inter3));
  inv1  gate1405(.a(s_123), .O(gate14inter4));
  nand2 gate1406(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1407(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1408(.a(G11), .O(gate14inter7));
  inv1  gate1409(.a(G12), .O(gate14inter8));
  nand2 gate1410(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1411(.a(s_123), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1412(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1413(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1414(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate729(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate730(.a(gate16inter0), .b(s_26), .O(gate16inter1));
  and2  gate731(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate732(.a(s_26), .O(gate16inter3));
  inv1  gate733(.a(s_27), .O(gate16inter4));
  nand2 gate734(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate735(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate736(.a(G15), .O(gate16inter7));
  inv1  gate737(.a(G16), .O(gate16inter8));
  nand2 gate738(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate739(.a(s_27), .b(gate16inter3), .O(gate16inter10));
  nor2  gate740(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate741(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate742(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate981(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate982(.a(gate24inter0), .b(s_62), .O(gate24inter1));
  and2  gate983(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate984(.a(s_62), .O(gate24inter3));
  inv1  gate985(.a(s_63), .O(gate24inter4));
  nand2 gate986(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate987(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate988(.a(G31), .O(gate24inter7));
  inv1  gate989(.a(G32), .O(gate24inter8));
  nand2 gate990(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate991(.a(s_63), .b(gate24inter3), .O(gate24inter10));
  nor2  gate992(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate993(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate994(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1023(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1024(.a(gate26inter0), .b(s_68), .O(gate26inter1));
  and2  gate1025(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1026(.a(s_68), .O(gate26inter3));
  inv1  gate1027(.a(s_69), .O(gate26inter4));
  nand2 gate1028(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1029(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1030(.a(G9), .O(gate26inter7));
  inv1  gate1031(.a(G13), .O(gate26inter8));
  nand2 gate1032(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1033(.a(s_69), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1034(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1035(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1036(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1457(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1458(.a(gate31inter0), .b(s_130), .O(gate31inter1));
  and2  gate1459(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1460(.a(s_130), .O(gate31inter3));
  inv1  gate1461(.a(s_131), .O(gate31inter4));
  nand2 gate1462(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1463(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1464(.a(G4), .O(gate31inter7));
  inv1  gate1465(.a(G8), .O(gate31inter8));
  nand2 gate1466(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1467(.a(s_131), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1468(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1469(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1470(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate855(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate856(.a(gate34inter0), .b(s_44), .O(gate34inter1));
  and2  gate857(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate858(.a(s_44), .O(gate34inter3));
  inv1  gate859(.a(s_45), .O(gate34inter4));
  nand2 gate860(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate861(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate862(.a(G25), .O(gate34inter7));
  inv1  gate863(.a(G29), .O(gate34inter8));
  nand2 gate864(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate865(.a(s_45), .b(gate34inter3), .O(gate34inter10));
  nor2  gate866(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate867(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate868(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1583(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1584(.a(gate40inter0), .b(s_148), .O(gate40inter1));
  and2  gate1585(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1586(.a(s_148), .O(gate40inter3));
  inv1  gate1587(.a(s_149), .O(gate40inter4));
  nand2 gate1588(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1589(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1590(.a(G28), .O(gate40inter7));
  inv1  gate1591(.a(G32), .O(gate40inter8));
  nand2 gate1592(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1593(.a(s_149), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1594(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1595(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1596(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1933(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1934(.a(gate60inter0), .b(s_198), .O(gate60inter1));
  and2  gate1935(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1936(.a(s_198), .O(gate60inter3));
  inv1  gate1937(.a(s_199), .O(gate60inter4));
  nand2 gate1938(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1939(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1940(.a(G20), .O(gate60inter7));
  inv1  gate1941(.a(G293), .O(gate60inter8));
  nand2 gate1942(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1943(.a(s_199), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1944(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1945(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1946(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate715(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate716(.a(gate62inter0), .b(s_24), .O(gate62inter1));
  and2  gate717(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate718(.a(s_24), .O(gate62inter3));
  inv1  gate719(.a(s_25), .O(gate62inter4));
  nand2 gate720(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate721(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate722(.a(G22), .O(gate62inter7));
  inv1  gate723(.a(G296), .O(gate62inter8));
  nand2 gate724(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate725(.a(s_25), .b(gate62inter3), .O(gate62inter10));
  nor2  gate726(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate727(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate728(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1205(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1206(.a(gate65inter0), .b(s_94), .O(gate65inter1));
  and2  gate1207(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1208(.a(s_94), .O(gate65inter3));
  inv1  gate1209(.a(s_95), .O(gate65inter4));
  nand2 gate1210(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1211(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1212(.a(G25), .O(gate65inter7));
  inv1  gate1213(.a(G302), .O(gate65inter8));
  nand2 gate1214(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1215(.a(s_95), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1216(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1217(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1218(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1219(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1220(.a(gate66inter0), .b(s_96), .O(gate66inter1));
  and2  gate1221(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1222(.a(s_96), .O(gate66inter3));
  inv1  gate1223(.a(s_97), .O(gate66inter4));
  nand2 gate1224(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1225(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1226(.a(G26), .O(gate66inter7));
  inv1  gate1227(.a(G302), .O(gate66inter8));
  nand2 gate1228(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1229(.a(s_97), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1230(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1231(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1232(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1079(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1080(.a(gate69inter0), .b(s_76), .O(gate69inter1));
  and2  gate1081(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1082(.a(s_76), .O(gate69inter3));
  inv1  gate1083(.a(s_77), .O(gate69inter4));
  nand2 gate1084(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1085(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1086(.a(G29), .O(gate69inter7));
  inv1  gate1087(.a(G308), .O(gate69inter8));
  nand2 gate1088(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1089(.a(s_77), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1090(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1091(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1092(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1387(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1388(.a(gate75inter0), .b(s_120), .O(gate75inter1));
  and2  gate1389(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1390(.a(s_120), .O(gate75inter3));
  inv1  gate1391(.a(s_121), .O(gate75inter4));
  nand2 gate1392(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1393(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1394(.a(G9), .O(gate75inter7));
  inv1  gate1395(.a(G317), .O(gate75inter8));
  nand2 gate1396(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1397(.a(s_121), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1398(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1399(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1400(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate687(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate688(.a(gate78inter0), .b(s_20), .O(gate78inter1));
  and2  gate689(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate690(.a(s_20), .O(gate78inter3));
  inv1  gate691(.a(s_21), .O(gate78inter4));
  nand2 gate692(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate693(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate694(.a(G6), .O(gate78inter7));
  inv1  gate695(.a(G320), .O(gate78inter8));
  nand2 gate696(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate697(.a(s_21), .b(gate78inter3), .O(gate78inter10));
  nor2  gate698(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate699(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate700(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1569(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1570(.a(gate80inter0), .b(s_146), .O(gate80inter1));
  and2  gate1571(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1572(.a(s_146), .O(gate80inter3));
  inv1  gate1573(.a(s_147), .O(gate80inter4));
  nand2 gate1574(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1575(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1576(.a(G14), .O(gate80inter7));
  inv1  gate1577(.a(G323), .O(gate80inter8));
  nand2 gate1578(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1579(.a(s_147), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1580(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1581(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1582(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1233(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1234(.a(gate83inter0), .b(s_98), .O(gate83inter1));
  and2  gate1235(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1236(.a(s_98), .O(gate83inter3));
  inv1  gate1237(.a(s_99), .O(gate83inter4));
  nand2 gate1238(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1239(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1240(.a(G11), .O(gate83inter7));
  inv1  gate1241(.a(G329), .O(gate83inter8));
  nand2 gate1242(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1243(.a(s_99), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1244(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1245(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1246(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate757(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate758(.a(gate87inter0), .b(s_30), .O(gate87inter1));
  and2  gate759(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate760(.a(s_30), .O(gate87inter3));
  inv1  gate761(.a(s_31), .O(gate87inter4));
  nand2 gate762(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate763(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate764(.a(G12), .O(gate87inter7));
  inv1  gate765(.a(G335), .O(gate87inter8));
  nand2 gate766(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate767(.a(s_31), .b(gate87inter3), .O(gate87inter10));
  nor2  gate768(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate769(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate770(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate589(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate590(.a(gate89inter0), .b(s_6), .O(gate89inter1));
  and2  gate591(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate592(.a(s_6), .O(gate89inter3));
  inv1  gate593(.a(s_7), .O(gate89inter4));
  nand2 gate594(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate595(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate596(.a(G17), .O(gate89inter7));
  inv1  gate597(.a(G338), .O(gate89inter8));
  nand2 gate598(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate599(.a(s_7), .b(gate89inter3), .O(gate89inter10));
  nor2  gate600(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate601(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate602(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate911(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate912(.a(gate92inter0), .b(s_52), .O(gate92inter1));
  and2  gate913(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate914(.a(s_52), .O(gate92inter3));
  inv1  gate915(.a(s_53), .O(gate92inter4));
  nand2 gate916(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate917(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate918(.a(G29), .O(gate92inter7));
  inv1  gate919(.a(G341), .O(gate92inter8));
  nand2 gate920(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate921(.a(s_53), .b(gate92inter3), .O(gate92inter10));
  nor2  gate922(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate923(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate924(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1373(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1374(.a(gate94inter0), .b(s_118), .O(gate94inter1));
  and2  gate1375(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1376(.a(s_118), .O(gate94inter3));
  inv1  gate1377(.a(s_119), .O(gate94inter4));
  nand2 gate1378(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1379(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1380(.a(G22), .O(gate94inter7));
  inv1  gate1381(.a(G344), .O(gate94inter8));
  nand2 gate1382(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1383(.a(s_119), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1384(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1385(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1386(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1009(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1010(.a(gate99inter0), .b(s_66), .O(gate99inter1));
  and2  gate1011(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1012(.a(s_66), .O(gate99inter3));
  inv1  gate1013(.a(s_67), .O(gate99inter4));
  nand2 gate1014(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1015(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1016(.a(G27), .O(gate99inter7));
  inv1  gate1017(.a(G353), .O(gate99inter8));
  nand2 gate1018(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1019(.a(s_67), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1020(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1021(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1022(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1485(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1486(.a(gate108inter0), .b(s_134), .O(gate108inter1));
  and2  gate1487(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1488(.a(s_134), .O(gate108inter3));
  inv1  gate1489(.a(s_135), .O(gate108inter4));
  nand2 gate1490(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1491(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1492(.a(G368), .O(gate108inter7));
  inv1  gate1493(.a(G369), .O(gate108inter8));
  nand2 gate1494(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1495(.a(s_135), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1496(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1497(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1498(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1331(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1332(.a(gate113inter0), .b(s_112), .O(gate113inter1));
  and2  gate1333(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1334(.a(s_112), .O(gate113inter3));
  inv1  gate1335(.a(s_113), .O(gate113inter4));
  nand2 gate1336(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1337(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1338(.a(G378), .O(gate113inter7));
  inv1  gate1339(.a(G379), .O(gate113inter8));
  nand2 gate1340(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1341(.a(s_113), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1342(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1343(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1344(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1471(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1472(.a(gate115inter0), .b(s_132), .O(gate115inter1));
  and2  gate1473(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1474(.a(s_132), .O(gate115inter3));
  inv1  gate1475(.a(s_133), .O(gate115inter4));
  nand2 gate1476(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1477(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1478(.a(G382), .O(gate115inter7));
  inv1  gate1479(.a(G383), .O(gate115inter8));
  nand2 gate1480(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1481(.a(s_133), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1482(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1483(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1484(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1415(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1416(.a(gate120inter0), .b(s_124), .O(gate120inter1));
  and2  gate1417(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1418(.a(s_124), .O(gate120inter3));
  inv1  gate1419(.a(s_125), .O(gate120inter4));
  nand2 gate1420(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1421(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1422(.a(G392), .O(gate120inter7));
  inv1  gate1423(.a(G393), .O(gate120inter8));
  nand2 gate1424(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1425(.a(s_125), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1426(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1427(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1428(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1513(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1514(.a(gate123inter0), .b(s_138), .O(gate123inter1));
  and2  gate1515(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1516(.a(s_138), .O(gate123inter3));
  inv1  gate1517(.a(s_139), .O(gate123inter4));
  nand2 gate1518(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1519(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1520(.a(G398), .O(gate123inter7));
  inv1  gate1521(.a(G399), .O(gate123inter8));
  nand2 gate1522(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1523(.a(s_139), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1524(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1525(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1526(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1597(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1598(.a(gate126inter0), .b(s_150), .O(gate126inter1));
  and2  gate1599(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1600(.a(s_150), .O(gate126inter3));
  inv1  gate1601(.a(s_151), .O(gate126inter4));
  nand2 gate1602(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1603(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1604(.a(G404), .O(gate126inter7));
  inv1  gate1605(.a(G405), .O(gate126inter8));
  nand2 gate1606(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1607(.a(s_151), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1608(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1609(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1610(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1695(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1696(.a(gate128inter0), .b(s_164), .O(gate128inter1));
  and2  gate1697(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1698(.a(s_164), .O(gate128inter3));
  inv1  gate1699(.a(s_165), .O(gate128inter4));
  nand2 gate1700(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1701(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1702(.a(G408), .O(gate128inter7));
  inv1  gate1703(.a(G409), .O(gate128inter8));
  nand2 gate1704(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1705(.a(s_165), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1706(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1707(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1708(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate897(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate898(.a(gate129inter0), .b(s_50), .O(gate129inter1));
  and2  gate899(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate900(.a(s_50), .O(gate129inter3));
  inv1  gate901(.a(s_51), .O(gate129inter4));
  nand2 gate902(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate903(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate904(.a(G410), .O(gate129inter7));
  inv1  gate905(.a(G411), .O(gate129inter8));
  nand2 gate906(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate907(.a(s_51), .b(gate129inter3), .O(gate129inter10));
  nor2  gate908(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate909(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate910(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate813(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate814(.a(gate130inter0), .b(s_38), .O(gate130inter1));
  and2  gate815(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate816(.a(s_38), .O(gate130inter3));
  inv1  gate817(.a(s_39), .O(gate130inter4));
  nand2 gate818(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate819(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate820(.a(G412), .O(gate130inter7));
  inv1  gate821(.a(G413), .O(gate130inter8));
  nand2 gate822(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate823(.a(s_39), .b(gate130inter3), .O(gate130inter10));
  nor2  gate824(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate825(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate826(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate673(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate674(.a(gate131inter0), .b(s_18), .O(gate131inter1));
  and2  gate675(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate676(.a(s_18), .O(gate131inter3));
  inv1  gate677(.a(s_19), .O(gate131inter4));
  nand2 gate678(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate679(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate680(.a(G414), .O(gate131inter7));
  inv1  gate681(.a(G415), .O(gate131inter8));
  nand2 gate682(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate683(.a(s_19), .b(gate131inter3), .O(gate131inter10));
  nor2  gate684(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate685(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate686(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1821(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1822(.a(gate134inter0), .b(s_182), .O(gate134inter1));
  and2  gate1823(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1824(.a(s_182), .O(gate134inter3));
  inv1  gate1825(.a(s_183), .O(gate134inter4));
  nand2 gate1826(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1827(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1828(.a(G420), .O(gate134inter7));
  inv1  gate1829(.a(G421), .O(gate134inter8));
  nand2 gate1830(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1831(.a(s_183), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1832(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1833(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1834(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate1247(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1248(.a(gate135inter0), .b(s_100), .O(gate135inter1));
  and2  gate1249(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1250(.a(s_100), .O(gate135inter3));
  inv1  gate1251(.a(s_101), .O(gate135inter4));
  nand2 gate1252(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1253(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1254(.a(G422), .O(gate135inter7));
  inv1  gate1255(.a(G423), .O(gate135inter8));
  nand2 gate1256(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1257(.a(s_101), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1258(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1259(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1260(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate827(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate828(.a(gate136inter0), .b(s_40), .O(gate136inter1));
  and2  gate829(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate830(.a(s_40), .O(gate136inter3));
  inv1  gate831(.a(s_41), .O(gate136inter4));
  nand2 gate832(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate833(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate834(.a(G424), .O(gate136inter7));
  inv1  gate835(.a(G425), .O(gate136inter8));
  nand2 gate836(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate837(.a(s_41), .b(gate136inter3), .O(gate136inter10));
  nor2  gate838(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate839(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate840(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate603(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate604(.a(gate139inter0), .b(s_8), .O(gate139inter1));
  and2  gate605(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate606(.a(s_8), .O(gate139inter3));
  inv1  gate607(.a(s_9), .O(gate139inter4));
  nand2 gate608(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate609(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate610(.a(G438), .O(gate139inter7));
  inv1  gate611(.a(G441), .O(gate139inter8));
  nand2 gate612(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate613(.a(s_9), .b(gate139inter3), .O(gate139inter10));
  nor2  gate614(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate615(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate616(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1625(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1626(.a(gate140inter0), .b(s_154), .O(gate140inter1));
  and2  gate1627(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1628(.a(s_154), .O(gate140inter3));
  inv1  gate1629(.a(s_155), .O(gate140inter4));
  nand2 gate1630(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1631(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1632(.a(G444), .O(gate140inter7));
  inv1  gate1633(.a(G447), .O(gate140inter8));
  nand2 gate1634(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1635(.a(s_155), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1636(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1637(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1638(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate799(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate800(.a(gate141inter0), .b(s_36), .O(gate141inter1));
  and2  gate801(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate802(.a(s_36), .O(gate141inter3));
  inv1  gate803(.a(s_37), .O(gate141inter4));
  nand2 gate804(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate805(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate806(.a(G450), .O(gate141inter7));
  inv1  gate807(.a(G453), .O(gate141inter8));
  nand2 gate808(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate809(.a(s_37), .b(gate141inter3), .O(gate141inter10));
  nor2  gate810(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate811(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate812(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate659(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate660(.a(gate143inter0), .b(s_16), .O(gate143inter1));
  and2  gate661(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate662(.a(s_16), .O(gate143inter3));
  inv1  gate663(.a(s_17), .O(gate143inter4));
  nand2 gate664(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate665(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate666(.a(G462), .O(gate143inter7));
  inv1  gate667(.a(G465), .O(gate143inter8));
  nand2 gate668(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate669(.a(s_17), .b(gate143inter3), .O(gate143inter10));
  nor2  gate670(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate671(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate672(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1037(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1038(.a(gate144inter0), .b(s_70), .O(gate144inter1));
  and2  gate1039(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1040(.a(s_70), .O(gate144inter3));
  inv1  gate1041(.a(s_71), .O(gate144inter4));
  nand2 gate1042(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1043(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1044(.a(G468), .O(gate144inter7));
  inv1  gate1045(.a(G471), .O(gate144inter8));
  nand2 gate1046(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1047(.a(s_71), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1048(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1049(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1050(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1443(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1444(.a(gate145inter0), .b(s_128), .O(gate145inter1));
  and2  gate1445(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1446(.a(s_128), .O(gate145inter3));
  inv1  gate1447(.a(s_129), .O(gate145inter4));
  nand2 gate1448(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1449(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1450(.a(G474), .O(gate145inter7));
  inv1  gate1451(.a(G477), .O(gate145inter8));
  nand2 gate1452(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1453(.a(s_129), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1454(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1455(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1456(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1541(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1542(.a(gate152inter0), .b(s_142), .O(gate152inter1));
  and2  gate1543(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1544(.a(s_142), .O(gate152inter3));
  inv1  gate1545(.a(s_143), .O(gate152inter4));
  nand2 gate1546(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1547(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1548(.a(G516), .O(gate152inter7));
  inv1  gate1549(.a(G519), .O(gate152inter8));
  nand2 gate1550(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1551(.a(s_143), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1552(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1553(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1554(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate785(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate786(.a(gate156inter0), .b(s_34), .O(gate156inter1));
  and2  gate787(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate788(.a(s_34), .O(gate156inter3));
  inv1  gate789(.a(s_35), .O(gate156inter4));
  nand2 gate790(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate791(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate792(.a(G435), .O(gate156inter7));
  inv1  gate793(.a(G525), .O(gate156inter8));
  nand2 gate794(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate795(.a(s_35), .b(gate156inter3), .O(gate156inter10));
  nor2  gate796(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate797(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate798(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1093(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1094(.a(gate159inter0), .b(s_78), .O(gate159inter1));
  and2  gate1095(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1096(.a(s_78), .O(gate159inter3));
  inv1  gate1097(.a(s_79), .O(gate159inter4));
  nand2 gate1098(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1099(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1100(.a(G444), .O(gate159inter7));
  inv1  gate1101(.a(G531), .O(gate159inter8));
  nand2 gate1102(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1103(.a(s_79), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1104(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1105(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1106(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate953(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate954(.a(gate170inter0), .b(s_58), .O(gate170inter1));
  and2  gate955(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate956(.a(s_58), .O(gate170inter3));
  inv1  gate957(.a(s_59), .O(gate170inter4));
  nand2 gate958(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate959(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate960(.a(G477), .O(gate170inter7));
  inv1  gate961(.a(G546), .O(gate170inter8));
  nand2 gate962(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate963(.a(s_59), .b(gate170inter3), .O(gate170inter10));
  nor2  gate964(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate965(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate966(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1779(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1780(.a(gate172inter0), .b(s_176), .O(gate172inter1));
  and2  gate1781(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1782(.a(s_176), .O(gate172inter3));
  inv1  gate1783(.a(s_177), .O(gate172inter4));
  nand2 gate1784(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1785(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1786(.a(G483), .O(gate172inter7));
  inv1  gate1787(.a(G549), .O(gate172inter8));
  nand2 gate1788(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1789(.a(s_177), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1790(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1791(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1792(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1345(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1346(.a(gate175inter0), .b(s_114), .O(gate175inter1));
  and2  gate1347(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1348(.a(s_114), .O(gate175inter3));
  inv1  gate1349(.a(s_115), .O(gate175inter4));
  nand2 gate1350(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1351(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1352(.a(G492), .O(gate175inter7));
  inv1  gate1353(.a(G555), .O(gate175inter8));
  nand2 gate1354(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1355(.a(s_115), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1356(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1357(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1358(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1275(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1276(.a(gate181inter0), .b(s_104), .O(gate181inter1));
  and2  gate1277(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1278(.a(s_104), .O(gate181inter3));
  inv1  gate1279(.a(s_105), .O(gate181inter4));
  nand2 gate1280(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1281(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1282(.a(G510), .O(gate181inter7));
  inv1  gate1283(.a(G564), .O(gate181inter8));
  nand2 gate1284(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1285(.a(s_105), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1286(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1287(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1288(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1429(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1430(.a(gate185inter0), .b(s_126), .O(gate185inter1));
  and2  gate1431(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1432(.a(s_126), .O(gate185inter3));
  inv1  gate1433(.a(s_127), .O(gate185inter4));
  nand2 gate1434(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1435(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1436(.a(G570), .O(gate185inter7));
  inv1  gate1437(.a(G571), .O(gate185inter8));
  nand2 gate1438(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1439(.a(s_127), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1440(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1441(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1442(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1919(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1920(.a(gate186inter0), .b(s_196), .O(gate186inter1));
  and2  gate1921(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1922(.a(s_196), .O(gate186inter3));
  inv1  gate1923(.a(s_197), .O(gate186inter4));
  nand2 gate1924(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1925(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1926(.a(G572), .O(gate186inter7));
  inv1  gate1927(.a(G573), .O(gate186inter8));
  nand2 gate1928(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1929(.a(s_197), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1930(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1931(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1932(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1667(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1668(.a(gate197inter0), .b(s_160), .O(gate197inter1));
  and2  gate1669(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1670(.a(s_160), .O(gate197inter3));
  inv1  gate1671(.a(s_161), .O(gate197inter4));
  nand2 gate1672(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1673(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1674(.a(G594), .O(gate197inter7));
  inv1  gate1675(.a(G595), .O(gate197inter8));
  nand2 gate1676(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1677(.a(s_161), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1678(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1679(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1680(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate701(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate702(.a(gate199inter0), .b(s_22), .O(gate199inter1));
  and2  gate703(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate704(.a(s_22), .O(gate199inter3));
  inv1  gate705(.a(s_23), .O(gate199inter4));
  nand2 gate706(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate707(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate708(.a(G598), .O(gate199inter7));
  inv1  gate709(.a(G599), .O(gate199inter8));
  nand2 gate710(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate711(.a(s_23), .b(gate199inter3), .O(gate199inter10));
  nor2  gate712(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate713(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate714(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1149(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1150(.a(gate200inter0), .b(s_86), .O(gate200inter1));
  and2  gate1151(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1152(.a(s_86), .O(gate200inter3));
  inv1  gate1153(.a(s_87), .O(gate200inter4));
  nand2 gate1154(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1155(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1156(.a(G600), .O(gate200inter7));
  inv1  gate1157(.a(G601), .O(gate200inter8));
  nand2 gate1158(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1159(.a(s_87), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1160(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1161(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1162(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1191(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1192(.a(gate201inter0), .b(s_92), .O(gate201inter1));
  and2  gate1193(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1194(.a(s_92), .O(gate201inter3));
  inv1  gate1195(.a(s_93), .O(gate201inter4));
  nand2 gate1196(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1197(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1198(.a(G602), .O(gate201inter7));
  inv1  gate1199(.a(G607), .O(gate201inter8));
  nand2 gate1200(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1201(.a(s_93), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1202(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1203(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1204(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1681(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1682(.a(gate202inter0), .b(s_162), .O(gate202inter1));
  and2  gate1683(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1684(.a(s_162), .O(gate202inter3));
  inv1  gate1685(.a(s_163), .O(gate202inter4));
  nand2 gate1686(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1687(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1688(.a(G612), .O(gate202inter7));
  inv1  gate1689(.a(G617), .O(gate202inter8));
  nand2 gate1690(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1691(.a(s_163), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1692(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1693(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1694(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1289(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1290(.a(gate203inter0), .b(s_106), .O(gate203inter1));
  and2  gate1291(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1292(.a(s_106), .O(gate203inter3));
  inv1  gate1293(.a(s_107), .O(gate203inter4));
  nand2 gate1294(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1295(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1296(.a(G602), .O(gate203inter7));
  inv1  gate1297(.a(G612), .O(gate203inter8));
  nand2 gate1298(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1299(.a(s_107), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1300(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1301(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1302(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate645(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate646(.a(gate208inter0), .b(s_14), .O(gate208inter1));
  and2  gate647(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate648(.a(s_14), .O(gate208inter3));
  inv1  gate649(.a(s_15), .O(gate208inter4));
  nand2 gate650(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate651(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate652(.a(G627), .O(gate208inter7));
  inv1  gate653(.a(G637), .O(gate208inter8));
  nand2 gate654(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate655(.a(s_15), .b(gate208inter3), .O(gate208inter10));
  nor2  gate656(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate657(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate658(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1555(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1556(.a(gate209inter0), .b(s_144), .O(gate209inter1));
  and2  gate1557(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1558(.a(s_144), .O(gate209inter3));
  inv1  gate1559(.a(s_145), .O(gate209inter4));
  nand2 gate1560(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1561(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1562(.a(G602), .O(gate209inter7));
  inv1  gate1563(.a(G666), .O(gate209inter8));
  nand2 gate1564(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1565(.a(s_145), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1566(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1567(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1568(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1835(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1836(.a(gate212inter0), .b(s_184), .O(gate212inter1));
  and2  gate1837(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1838(.a(s_184), .O(gate212inter3));
  inv1  gate1839(.a(s_185), .O(gate212inter4));
  nand2 gate1840(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1841(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1842(.a(G617), .O(gate212inter7));
  inv1  gate1843(.a(G669), .O(gate212inter8));
  nand2 gate1844(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1845(.a(s_185), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1846(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1847(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1848(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1849(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1850(.a(gate216inter0), .b(s_186), .O(gate216inter1));
  and2  gate1851(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1852(.a(s_186), .O(gate216inter3));
  inv1  gate1853(.a(s_187), .O(gate216inter4));
  nand2 gate1854(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1855(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1856(.a(G617), .O(gate216inter7));
  inv1  gate1857(.a(G675), .O(gate216inter8));
  nand2 gate1858(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1859(.a(s_187), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1860(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1861(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1862(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate995(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate996(.a(gate220inter0), .b(s_64), .O(gate220inter1));
  and2  gate997(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate998(.a(s_64), .O(gate220inter3));
  inv1  gate999(.a(s_65), .O(gate220inter4));
  nand2 gate1000(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1001(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1002(.a(G637), .O(gate220inter7));
  inv1  gate1003(.a(G681), .O(gate220inter8));
  nand2 gate1004(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1005(.a(s_65), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1006(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1007(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1008(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate883(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate884(.a(gate223inter0), .b(s_48), .O(gate223inter1));
  and2  gate885(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate886(.a(s_48), .O(gate223inter3));
  inv1  gate887(.a(s_49), .O(gate223inter4));
  nand2 gate888(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate889(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate890(.a(G627), .O(gate223inter7));
  inv1  gate891(.a(G687), .O(gate223inter8));
  nand2 gate892(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate893(.a(s_49), .b(gate223inter3), .O(gate223inter10));
  nor2  gate894(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate895(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate896(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate939(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate940(.a(gate229inter0), .b(s_56), .O(gate229inter1));
  and2  gate941(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate942(.a(s_56), .O(gate229inter3));
  inv1  gate943(.a(s_57), .O(gate229inter4));
  nand2 gate944(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate945(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate946(.a(G698), .O(gate229inter7));
  inv1  gate947(.a(G699), .O(gate229inter8));
  nand2 gate948(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate949(.a(s_57), .b(gate229inter3), .O(gate229inter10));
  nor2  gate950(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate951(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate952(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1121(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1122(.a(gate231inter0), .b(s_82), .O(gate231inter1));
  and2  gate1123(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1124(.a(s_82), .O(gate231inter3));
  inv1  gate1125(.a(s_83), .O(gate231inter4));
  nand2 gate1126(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1127(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1128(.a(G702), .O(gate231inter7));
  inv1  gate1129(.a(G703), .O(gate231inter8));
  nand2 gate1130(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1131(.a(s_83), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1132(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1133(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1134(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate841(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate842(.a(gate235inter0), .b(s_42), .O(gate235inter1));
  and2  gate843(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate844(.a(s_42), .O(gate235inter3));
  inv1  gate845(.a(s_43), .O(gate235inter4));
  nand2 gate846(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate847(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate848(.a(G248), .O(gate235inter7));
  inv1  gate849(.a(G724), .O(gate235inter8));
  nand2 gate850(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate851(.a(s_43), .b(gate235inter3), .O(gate235inter10));
  nor2  gate852(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate853(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate854(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1723(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1724(.a(gate237inter0), .b(s_168), .O(gate237inter1));
  and2  gate1725(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1726(.a(s_168), .O(gate237inter3));
  inv1  gate1727(.a(s_169), .O(gate237inter4));
  nand2 gate1728(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1729(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1730(.a(G254), .O(gate237inter7));
  inv1  gate1731(.a(G706), .O(gate237inter8));
  nand2 gate1732(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1733(.a(s_169), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1734(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1735(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1736(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate771(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate772(.a(gate257inter0), .b(s_32), .O(gate257inter1));
  and2  gate773(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate774(.a(s_32), .O(gate257inter3));
  inv1  gate775(.a(s_33), .O(gate257inter4));
  nand2 gate776(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate777(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate778(.a(G754), .O(gate257inter7));
  inv1  gate779(.a(G755), .O(gate257inter8));
  nand2 gate780(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate781(.a(s_33), .b(gate257inter3), .O(gate257inter10));
  nor2  gate782(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate783(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate784(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate869(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate870(.a(gate263inter0), .b(s_46), .O(gate263inter1));
  and2  gate871(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate872(.a(s_46), .O(gate263inter3));
  inv1  gate873(.a(s_47), .O(gate263inter4));
  nand2 gate874(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate875(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate876(.a(G766), .O(gate263inter7));
  inv1  gate877(.a(G767), .O(gate263inter8));
  nand2 gate878(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate879(.a(s_47), .b(gate263inter3), .O(gate263inter10));
  nor2  gate880(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate881(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate882(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1765(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1766(.a(gate278inter0), .b(s_174), .O(gate278inter1));
  and2  gate1767(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1768(.a(s_174), .O(gate278inter3));
  inv1  gate1769(.a(s_175), .O(gate278inter4));
  nand2 gate1770(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1771(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1772(.a(G776), .O(gate278inter7));
  inv1  gate1773(.a(G800), .O(gate278inter8));
  nand2 gate1774(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1775(.a(s_175), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1776(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1777(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1778(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1163(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1164(.a(gate286inter0), .b(s_88), .O(gate286inter1));
  and2  gate1165(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1166(.a(s_88), .O(gate286inter3));
  inv1  gate1167(.a(s_89), .O(gate286inter4));
  nand2 gate1168(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1169(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1170(.a(G788), .O(gate286inter7));
  inv1  gate1171(.a(G812), .O(gate286inter8));
  nand2 gate1172(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1173(.a(s_89), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1174(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1175(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1176(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1737(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1738(.a(gate289inter0), .b(s_170), .O(gate289inter1));
  and2  gate1739(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1740(.a(s_170), .O(gate289inter3));
  inv1  gate1741(.a(s_171), .O(gate289inter4));
  nand2 gate1742(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1743(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1744(.a(G818), .O(gate289inter7));
  inv1  gate1745(.a(G819), .O(gate289inter8));
  nand2 gate1746(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1747(.a(s_171), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1748(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1749(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1750(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1065(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1066(.a(gate292inter0), .b(s_74), .O(gate292inter1));
  and2  gate1067(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1068(.a(s_74), .O(gate292inter3));
  inv1  gate1069(.a(s_75), .O(gate292inter4));
  nand2 gate1070(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1071(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1072(.a(G824), .O(gate292inter7));
  inv1  gate1073(.a(G825), .O(gate292inter8));
  nand2 gate1074(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1075(.a(s_75), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1076(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1077(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1078(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate575(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate576(.a(gate296inter0), .b(s_4), .O(gate296inter1));
  and2  gate577(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate578(.a(s_4), .O(gate296inter3));
  inv1  gate579(.a(s_5), .O(gate296inter4));
  nand2 gate580(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate581(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate582(.a(G826), .O(gate296inter7));
  inv1  gate583(.a(G827), .O(gate296inter8));
  nand2 gate584(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate585(.a(s_5), .b(gate296inter3), .O(gate296inter10));
  nor2  gate586(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate587(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate588(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1863(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1864(.a(gate392inter0), .b(s_188), .O(gate392inter1));
  and2  gate1865(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1866(.a(s_188), .O(gate392inter3));
  inv1  gate1867(.a(s_189), .O(gate392inter4));
  nand2 gate1868(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1869(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1870(.a(G6), .O(gate392inter7));
  inv1  gate1871(.a(G1051), .O(gate392inter8));
  nand2 gate1872(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1873(.a(s_189), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1874(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1875(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1876(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1905(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1906(.a(gate396inter0), .b(s_194), .O(gate396inter1));
  and2  gate1907(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1908(.a(s_194), .O(gate396inter3));
  inv1  gate1909(.a(s_195), .O(gate396inter4));
  nand2 gate1910(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1911(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1912(.a(G10), .O(gate396inter7));
  inv1  gate1913(.a(G1063), .O(gate396inter8));
  nand2 gate1914(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1915(.a(s_195), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1916(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1917(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1918(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1751(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1752(.a(gate398inter0), .b(s_172), .O(gate398inter1));
  and2  gate1753(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1754(.a(s_172), .O(gate398inter3));
  inv1  gate1755(.a(s_173), .O(gate398inter4));
  nand2 gate1756(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1757(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1758(.a(G12), .O(gate398inter7));
  inv1  gate1759(.a(G1069), .O(gate398inter8));
  nand2 gate1760(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1761(.a(s_173), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1762(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1763(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1764(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1499(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1500(.a(gate399inter0), .b(s_136), .O(gate399inter1));
  and2  gate1501(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1502(.a(s_136), .O(gate399inter3));
  inv1  gate1503(.a(s_137), .O(gate399inter4));
  nand2 gate1504(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1505(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1506(.a(G13), .O(gate399inter7));
  inv1  gate1507(.a(G1072), .O(gate399inter8));
  nand2 gate1508(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1509(.a(s_137), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1510(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1511(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1512(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1877(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1878(.a(gate405inter0), .b(s_190), .O(gate405inter1));
  and2  gate1879(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1880(.a(s_190), .O(gate405inter3));
  inv1  gate1881(.a(s_191), .O(gate405inter4));
  nand2 gate1882(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1883(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1884(.a(G19), .O(gate405inter7));
  inv1  gate1885(.a(G1090), .O(gate405inter8));
  nand2 gate1886(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1887(.a(s_191), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1888(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1889(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1890(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1653(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1654(.a(gate407inter0), .b(s_158), .O(gate407inter1));
  and2  gate1655(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1656(.a(s_158), .O(gate407inter3));
  inv1  gate1657(.a(s_159), .O(gate407inter4));
  nand2 gate1658(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1659(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1660(.a(G21), .O(gate407inter7));
  inv1  gate1661(.a(G1096), .O(gate407inter8));
  nand2 gate1662(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1663(.a(s_159), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1664(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1665(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1666(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1107(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1108(.a(gate413inter0), .b(s_80), .O(gate413inter1));
  and2  gate1109(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1110(.a(s_80), .O(gate413inter3));
  inv1  gate1111(.a(s_81), .O(gate413inter4));
  nand2 gate1112(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1113(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1114(.a(G27), .O(gate413inter7));
  inv1  gate1115(.a(G1114), .O(gate413inter8));
  nand2 gate1116(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1117(.a(s_81), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1118(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1119(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1120(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1807(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1808(.a(gate416inter0), .b(s_180), .O(gate416inter1));
  and2  gate1809(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1810(.a(s_180), .O(gate416inter3));
  inv1  gate1811(.a(s_181), .O(gate416inter4));
  nand2 gate1812(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1813(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1814(.a(G30), .O(gate416inter7));
  inv1  gate1815(.a(G1123), .O(gate416inter8));
  nand2 gate1816(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1817(.a(s_181), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1818(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1819(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1820(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1793(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1794(.a(gate426inter0), .b(s_178), .O(gate426inter1));
  and2  gate1795(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1796(.a(s_178), .O(gate426inter3));
  inv1  gate1797(.a(s_179), .O(gate426inter4));
  nand2 gate1798(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1799(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1800(.a(G1045), .O(gate426inter7));
  inv1  gate1801(.a(G1141), .O(gate426inter8));
  nand2 gate1802(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1803(.a(s_179), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1804(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1805(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1806(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate967(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate968(.a(gate430inter0), .b(s_60), .O(gate430inter1));
  and2  gate969(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate970(.a(s_60), .O(gate430inter3));
  inv1  gate971(.a(s_61), .O(gate430inter4));
  nand2 gate972(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate973(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate974(.a(G1051), .O(gate430inter7));
  inv1  gate975(.a(G1147), .O(gate430inter8));
  nand2 gate976(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate977(.a(s_61), .b(gate430inter3), .O(gate430inter10));
  nor2  gate978(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate979(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate980(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1639(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1640(.a(gate435inter0), .b(s_156), .O(gate435inter1));
  and2  gate1641(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1642(.a(s_156), .O(gate435inter3));
  inv1  gate1643(.a(s_157), .O(gate435inter4));
  nand2 gate1644(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1645(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1646(.a(G9), .O(gate435inter7));
  inv1  gate1647(.a(G1156), .O(gate435inter8));
  nand2 gate1648(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1649(.a(s_157), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1650(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1651(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1652(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1303(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1304(.a(gate441inter0), .b(s_108), .O(gate441inter1));
  and2  gate1305(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1306(.a(s_108), .O(gate441inter3));
  inv1  gate1307(.a(s_109), .O(gate441inter4));
  nand2 gate1308(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1309(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1310(.a(G12), .O(gate441inter7));
  inv1  gate1311(.a(G1165), .O(gate441inter8));
  nand2 gate1312(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1313(.a(s_109), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1314(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1315(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1316(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1261(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1262(.a(gate447inter0), .b(s_102), .O(gate447inter1));
  and2  gate1263(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1264(.a(s_102), .O(gate447inter3));
  inv1  gate1265(.a(s_103), .O(gate447inter4));
  nand2 gate1266(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1267(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1268(.a(G15), .O(gate447inter7));
  inv1  gate1269(.a(G1174), .O(gate447inter8));
  nand2 gate1270(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1271(.a(s_103), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1272(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1273(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1274(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1317(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1318(.a(gate460inter0), .b(s_110), .O(gate460inter1));
  and2  gate1319(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1320(.a(s_110), .O(gate460inter3));
  inv1  gate1321(.a(s_111), .O(gate460inter4));
  nand2 gate1322(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1323(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1324(.a(G1096), .O(gate460inter7));
  inv1  gate1325(.a(G1192), .O(gate460inter8));
  nand2 gate1326(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1327(.a(s_111), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1328(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1329(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1330(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate561(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate562(.a(gate465inter0), .b(s_2), .O(gate465inter1));
  and2  gate563(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate564(.a(s_2), .O(gate465inter3));
  inv1  gate565(.a(s_3), .O(gate465inter4));
  nand2 gate566(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate567(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate568(.a(G24), .O(gate465inter7));
  inv1  gate569(.a(G1201), .O(gate465inter8));
  nand2 gate570(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate571(.a(s_3), .b(gate465inter3), .O(gate465inter10));
  nor2  gate572(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate573(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate574(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate617(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate618(.a(gate472inter0), .b(s_10), .O(gate472inter1));
  and2  gate619(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate620(.a(s_10), .O(gate472inter3));
  inv1  gate621(.a(s_11), .O(gate472inter4));
  nand2 gate622(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate623(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate624(.a(G1114), .O(gate472inter7));
  inv1  gate625(.a(G1210), .O(gate472inter8));
  nand2 gate626(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate627(.a(s_11), .b(gate472inter3), .O(gate472inter10));
  nor2  gate628(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate629(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate630(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1177(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1178(.a(gate474inter0), .b(s_90), .O(gate474inter1));
  and2  gate1179(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1180(.a(s_90), .O(gate474inter3));
  inv1  gate1181(.a(s_91), .O(gate474inter4));
  nand2 gate1182(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1183(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1184(.a(G1117), .O(gate474inter7));
  inv1  gate1185(.a(G1213), .O(gate474inter8));
  nand2 gate1186(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1187(.a(s_91), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1188(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1189(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1190(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1709(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1710(.a(gate480inter0), .b(s_166), .O(gate480inter1));
  and2  gate1711(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1712(.a(s_166), .O(gate480inter3));
  inv1  gate1713(.a(s_167), .O(gate480inter4));
  nand2 gate1714(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1715(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1716(.a(G1126), .O(gate480inter7));
  inv1  gate1717(.a(G1222), .O(gate480inter8));
  nand2 gate1718(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1719(.a(s_167), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1720(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1721(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1722(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1135(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1136(.a(gate485inter0), .b(s_84), .O(gate485inter1));
  and2  gate1137(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1138(.a(s_84), .O(gate485inter3));
  inv1  gate1139(.a(s_85), .O(gate485inter4));
  nand2 gate1140(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1141(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1142(.a(G1232), .O(gate485inter7));
  inv1  gate1143(.a(G1233), .O(gate485inter8));
  nand2 gate1144(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1145(.a(s_85), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1146(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1147(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1148(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate547(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate548(.a(gate491inter0), .b(s_0), .O(gate491inter1));
  and2  gate549(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate550(.a(s_0), .O(gate491inter3));
  inv1  gate551(.a(s_1), .O(gate491inter4));
  nand2 gate552(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate553(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate554(.a(G1244), .O(gate491inter7));
  inv1  gate555(.a(G1245), .O(gate491inter8));
  nand2 gate556(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate557(.a(s_1), .b(gate491inter3), .O(gate491inter10));
  nor2  gate558(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate559(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate560(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1359(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1360(.a(gate501inter0), .b(s_116), .O(gate501inter1));
  and2  gate1361(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1362(.a(s_116), .O(gate501inter3));
  inv1  gate1363(.a(s_117), .O(gate501inter4));
  nand2 gate1364(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1365(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1366(.a(G1264), .O(gate501inter7));
  inv1  gate1367(.a(G1265), .O(gate501inter8));
  nand2 gate1368(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1369(.a(s_117), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1370(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1371(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1372(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1611(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1612(.a(gate503inter0), .b(s_152), .O(gate503inter1));
  and2  gate1613(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1614(.a(s_152), .O(gate503inter3));
  inv1  gate1615(.a(s_153), .O(gate503inter4));
  nand2 gate1616(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1617(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1618(.a(G1268), .O(gate503inter7));
  inv1  gate1619(.a(G1269), .O(gate503inter8));
  nand2 gate1620(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1621(.a(s_153), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1622(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1623(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1624(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1947(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1948(.a(gate505inter0), .b(s_200), .O(gate505inter1));
  and2  gate1949(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1950(.a(s_200), .O(gate505inter3));
  inv1  gate1951(.a(s_201), .O(gate505inter4));
  nand2 gate1952(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1953(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1954(.a(G1272), .O(gate505inter7));
  inv1  gate1955(.a(G1273), .O(gate505inter8));
  nand2 gate1956(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1957(.a(s_201), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1958(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1959(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1960(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate631(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate632(.a(gate506inter0), .b(s_12), .O(gate506inter1));
  and2  gate633(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate634(.a(s_12), .O(gate506inter3));
  inv1  gate635(.a(s_13), .O(gate506inter4));
  nand2 gate636(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate637(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate638(.a(G1274), .O(gate506inter7));
  inv1  gate639(.a(G1275), .O(gate506inter8));
  nand2 gate640(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate641(.a(s_13), .b(gate506inter3), .O(gate506inter10));
  nor2  gate642(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate643(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate644(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1891(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1892(.a(gate508inter0), .b(s_192), .O(gate508inter1));
  and2  gate1893(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1894(.a(s_192), .O(gate508inter3));
  inv1  gate1895(.a(s_193), .O(gate508inter4));
  nand2 gate1896(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1897(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1898(.a(G1278), .O(gate508inter7));
  inv1  gate1899(.a(G1279), .O(gate508inter8));
  nand2 gate1900(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1901(.a(s_193), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1902(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1903(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1904(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate743(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate744(.a(gate511inter0), .b(s_28), .O(gate511inter1));
  and2  gate745(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate746(.a(s_28), .O(gate511inter3));
  inv1  gate747(.a(s_29), .O(gate511inter4));
  nand2 gate748(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate749(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate750(.a(G1284), .O(gate511inter7));
  inv1  gate751(.a(G1285), .O(gate511inter8));
  nand2 gate752(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate753(.a(s_29), .b(gate511inter3), .O(gate511inter10));
  nor2  gate754(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate755(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate756(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1527(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1528(.a(gate512inter0), .b(s_140), .O(gate512inter1));
  and2  gate1529(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1530(.a(s_140), .O(gate512inter3));
  inv1  gate1531(.a(s_141), .O(gate512inter4));
  nand2 gate1532(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1533(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1534(.a(G1286), .O(gate512inter7));
  inv1  gate1535(.a(G1287), .O(gate512inter8));
  nand2 gate1536(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1537(.a(s_141), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1538(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1539(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1540(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule