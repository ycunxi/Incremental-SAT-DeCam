module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate858inter0, gate858inter1, gate858inter2, gate858inter3, gate858inter4, gate858inter5, gate858inter6, gate858inter7, gate858inter8, gate858inter9, gate858inter10, gate858inter11, gate858inter12, gate875inter0, gate875inter1, gate875inter2, gate875inter3, gate875inter4, gate875inter5, gate875inter6, gate875inter7, gate875inter8, gate875inter9, gate875inter10, gate875inter11, gate875inter12, gate819inter0, gate819inter1, gate819inter2, gate819inter3, gate819inter4, gate819inter5, gate819inter6, gate819inter7, gate819inter8, gate819inter9, gate819inter10, gate819inter11, gate819inter12, gate636inter0, gate636inter1, gate636inter2, gate636inter3, gate636inter4, gate636inter5, gate636inter6, gate636inter7, gate636inter8, gate636inter9, gate636inter10, gate636inter11, gate636inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate803inter0, gate803inter1, gate803inter2, gate803inter3, gate803inter4, gate803inter5, gate803inter6, gate803inter7, gate803inter8, gate803inter9, gate803inter10, gate803inter11, gate803inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate539inter0, gate539inter1, gate539inter2, gate539inter3, gate539inter4, gate539inter5, gate539inter6, gate539inter7, gate539inter8, gate539inter9, gate539inter10, gate539inter11, gate539inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate526inter0, gate526inter1, gate526inter2, gate526inter3, gate526inter4, gate526inter5, gate526inter6, gate526inter7, gate526inter8, gate526inter9, gate526inter10, gate526inter11, gate526inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate789inter0, gate789inter1, gate789inter2, gate789inter3, gate789inter4, gate789inter5, gate789inter6, gate789inter7, gate789inter8, gate789inter9, gate789inter10, gate789inter11, gate789inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate828inter0, gate828inter1, gate828inter2, gate828inter3, gate828inter4, gate828inter5, gate828inter6, gate828inter7, gate828inter8, gate828inter9, gate828inter10, gate828inter11, gate828inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate550inter0, gate550inter1, gate550inter2, gate550inter3, gate550inter4, gate550inter5, gate550inter6, gate550inter7, gate550inter8, gate550inter9, gate550inter10, gate550inter11, gate550inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate876inter0, gate876inter1, gate876inter2, gate876inter3, gate876inter4, gate876inter5, gate876inter6, gate876inter7, gate876inter8, gate876inter9, gate876inter10, gate876inter11, gate876inter12, gate758inter0, gate758inter1, gate758inter2, gate758inter3, gate758inter4, gate758inter5, gate758inter6, gate758inter7, gate758inter8, gate758inter9, gate758inter10, gate758inter11, gate758inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate320inter0, gate320inter1, gate320inter2, gate320inter3, gate320inter4, gate320inter5, gate320inter6, gate320inter7, gate320inter8, gate320inter9, gate320inter10, gate320inter11, gate320inter12, gate854inter0, gate854inter1, gate854inter2, gate854inter3, gate854inter4, gate854inter5, gate854inter6, gate854inter7, gate854inter8, gate854inter9, gate854inter10, gate854inter11, gate854inter12, gate561inter0, gate561inter1, gate561inter2, gate561inter3, gate561inter4, gate561inter5, gate561inter6, gate561inter7, gate561inter8, gate561inter9, gate561inter10, gate561inter11, gate561inter12, gate820inter0, gate820inter1, gate820inter2, gate820inter3, gate820inter4, gate820inter5, gate820inter6, gate820inter7, gate820inter8, gate820inter9, gate820inter10, gate820inter11, gate820inter12, gate605inter0, gate605inter1, gate605inter2, gate605inter3, gate605inter4, gate605inter5, gate605inter6, gate605inter7, gate605inter8, gate605inter9, gate605inter10, gate605inter11, gate605inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate631inter0, gate631inter1, gate631inter2, gate631inter3, gate631inter4, gate631inter5, gate631inter6, gate631inter7, gate631inter8, gate631inter9, gate631inter10, gate631inter11, gate631inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate809inter0, gate809inter1, gate809inter2, gate809inter3, gate809inter4, gate809inter5, gate809inter6, gate809inter7, gate809inter8, gate809inter9, gate809inter10, gate809inter11, gate809inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate750inter0, gate750inter1, gate750inter2, gate750inter3, gate750inter4, gate750inter5, gate750inter6, gate750inter7, gate750inter8, gate750inter9, gate750inter10, gate750inter11, gate750inter12, gate867inter0, gate867inter1, gate867inter2, gate867inter3, gate867inter4, gate867inter5, gate867inter6, gate867inter7, gate867inter8, gate867inter9, gate867inter10, gate867inter11, gate867inter12, gate527inter0, gate527inter1, gate527inter2, gate527inter3, gate527inter4, gate527inter5, gate527inter6, gate527inter7, gate527inter8, gate527inter9, gate527inter10, gate527inter11, gate527inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate345inter0, gate345inter1, gate345inter2, gate345inter3, gate345inter4, gate345inter5, gate345inter6, gate345inter7, gate345inter8, gate345inter9, gate345inter10, gate345inter11, gate345inter12, gate542inter0, gate542inter1, gate542inter2, gate542inter3, gate542inter4, gate542inter5, gate542inter6, gate542inter7, gate542inter8, gate542inter9, gate542inter10, gate542inter11, gate542inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate775inter0, gate775inter1, gate775inter2, gate775inter3, gate775inter4, gate775inter5, gate775inter6, gate775inter7, gate775inter8, gate775inter9, gate775inter10, gate775inter11, gate775inter12, gate519inter0, gate519inter1, gate519inter2, gate519inter3, gate519inter4, gate519inter5, gate519inter6, gate519inter7, gate519inter8, gate519inter9, gate519inter10, gate519inter11, gate519inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate850inter0, gate850inter1, gate850inter2, gate850inter3, gate850inter4, gate850inter5, gate850inter6, gate850inter7, gate850inter8, gate850inter9, gate850inter10, gate850inter11, gate850inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate572inter0, gate572inter1, gate572inter2, gate572inter3, gate572inter4, gate572inter5, gate572inter6, gate572inter7, gate572inter8, gate572inter9, gate572inter10, gate572inter11, gate572inter12, gate802inter0, gate802inter1, gate802inter2, gate802inter3, gate802inter4, gate802inter5, gate802inter6, gate802inter7, gate802inter8, gate802inter9, gate802inter10, gate802inter11, gate802inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate632inter0, gate632inter1, gate632inter2, gate632inter3, gate632inter4, gate632inter5, gate632inter6, gate632inter7, gate632inter8, gate632inter9, gate632inter10, gate632inter11, gate632inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate318inter0, gate318inter1, gate318inter2, gate318inter3, gate318inter4, gate318inter5, gate318inter6, gate318inter7, gate318inter8, gate318inter9, gate318inter10, gate318inter11, gate318inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );

  xor2  gate1945(.a(N331), .b(N306), .O(gate75inter0));
  nand2 gate1946(.a(gate75inter0), .b(s_152), .O(gate75inter1));
  and2  gate1947(.a(N331), .b(N306), .O(gate75inter2));
  inv1  gate1948(.a(s_152), .O(gate75inter3));
  inv1  gate1949(.a(s_153), .O(gate75inter4));
  nand2 gate1950(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1951(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1952(.a(N306), .O(gate75inter7));
  inv1  gate1953(.a(N331), .O(gate75inter8));
  nand2 gate1954(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1955(.a(s_153), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1956(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1957(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1958(.a(gate75inter12), .b(gate75inter1), .O(N550));
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate1973(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate1974(.a(gate96inter0), .b(s_156), .O(gate96inter1));
  and2  gate1975(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate1976(.a(s_156), .O(gate96inter3));
  inv1  gate1977(.a(s_157), .O(gate96inter4));
  nand2 gate1978(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1979(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1980(.a(N326), .O(gate96inter7));
  inv1  gate1981(.a(N277), .O(gate96inter8));
  nand2 gate1982(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1983(.a(s_157), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1984(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1985(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1986(.a(gate96inter12), .b(gate96inter1), .O(N601));
nand2 gate97( .a(N326), .b(N280), .O(N602) );

  xor2  gate1749(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate1750(.a(gate98inter0), .b(s_124), .O(gate98inter1));
  and2  gate1751(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate1752(.a(s_124), .O(gate98inter3));
  inv1  gate1753(.a(s_125), .O(gate98inter4));
  nand2 gate1754(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1755(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1756(.a(N260), .O(gate98inter7));
  inv1  gate1757(.a(N72), .O(gate98inter8));
  nand2 gate1758(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1759(.a(s_125), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1760(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1761(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1762(.a(gate98inter12), .b(gate98inter1), .O(N603));
nand2 gate99( .a(N260), .b(N300), .O(N608) );

  xor2  gate1147(.a(N300), .b(N256), .O(gate100inter0));
  nand2 gate1148(.a(gate100inter0), .b(s_38), .O(gate100inter1));
  and2  gate1149(.a(N300), .b(N256), .O(gate100inter2));
  inv1  gate1150(.a(s_38), .O(gate100inter3));
  inv1  gate1151(.a(s_39), .O(gate100inter4));
  nand2 gate1152(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1153(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1154(.a(N256), .O(gate100inter7));
  inv1  gate1155(.a(N300), .O(gate100inter8));
  nand2 gate1156(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1157(.a(s_39), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1158(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1159(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1160(.a(gate100inter12), .b(gate100inter1), .O(N612));
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );

  xor2  gate965(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate966(.a(gate236inter0), .b(s_12), .O(gate236inter1));
  and2  gate967(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate968(.a(s_12), .O(gate236inter3));
  inv1  gate969(.a(s_13), .O(gate236inter4));
  nand2 gate970(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate971(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate972(.a(N622), .O(gate236inter7));
  inv1  gate973(.a(N891), .O(gate236inter8));
  nand2 gate974(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate975(.a(s_13), .b(gate236inter3), .O(gate236inter10));
  nor2  gate976(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate977(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate978(.a(gate236inter12), .b(gate236inter1), .O(N1064));

  xor2  gate1217(.a(N895), .b(N655), .O(gate237inter0));
  nand2 gate1218(.a(gate237inter0), .b(s_48), .O(gate237inter1));
  and2  gate1219(.a(N895), .b(N655), .O(gate237inter2));
  inv1  gate1220(.a(s_48), .O(gate237inter3));
  inv1  gate1221(.a(s_49), .O(gate237inter4));
  nand2 gate1222(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1223(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1224(.a(N655), .O(gate237inter7));
  inv1  gate1225(.a(N895), .O(gate237inter8));
  nand2 gate1226(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1227(.a(s_49), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1228(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1229(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1230(.a(gate237inter12), .b(gate237inter1), .O(N1067));

  xor2  gate1581(.a(N896), .b(N652), .O(gate238inter0));
  nand2 gate1582(.a(gate238inter0), .b(s_100), .O(gate238inter1));
  and2  gate1583(.a(N896), .b(N652), .O(gate238inter2));
  inv1  gate1584(.a(s_100), .O(gate238inter3));
  inv1  gate1585(.a(s_101), .O(gate238inter4));
  nand2 gate1586(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1587(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1588(.a(N652), .O(gate238inter7));
  inv1  gate1589(.a(N896), .O(gate238inter8));
  nand2 gate1590(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1591(.a(s_101), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1592(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1593(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1594(.a(gate238inter12), .b(gate238inter1), .O(N1068));
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );

  xor2  gate1063(.a(N991), .b(N727), .O(gate241inter0));
  nand2 gate1064(.a(gate241inter0), .b(s_26), .O(gate241inter1));
  and2  gate1065(.a(N991), .b(N727), .O(gate241inter2));
  inv1  gate1066(.a(s_26), .O(gate241inter3));
  inv1  gate1067(.a(s_27), .O(gate241inter4));
  nand2 gate1068(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1069(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1070(.a(N727), .O(gate241inter7));
  inv1  gate1071(.a(N991), .O(gate241inter8));
  nand2 gate1072(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1073(.a(s_27), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1074(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1075(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1076(.a(gate241inter12), .b(gate241inter1), .O(N1121));
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );

  xor2  gate1161(.a(N1009), .b(N748), .O(gate248inter0));
  nand2 gate1162(.a(gate248inter0), .b(s_40), .O(gate248inter1));
  and2  gate1163(.a(N1009), .b(N748), .O(gate248inter2));
  inv1  gate1164(.a(s_40), .O(gate248inter3));
  inv1  gate1165(.a(s_41), .O(gate248inter4));
  nand2 gate1166(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1167(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1168(.a(N748), .O(gate248inter7));
  inv1  gate1169(.a(N1009), .O(gate248inter8));
  nand2 gate1170(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1171(.a(s_41), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1172(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1173(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1174(.a(gate248inter12), .b(gate248inter1), .O(N1133));
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );

  xor2  gate1231(.a(N1064), .b(N1063), .O(gate259inter0));
  nand2 gate1232(.a(gate259inter0), .b(s_50), .O(gate259inter1));
  and2  gate1233(.a(N1064), .b(N1063), .O(gate259inter2));
  inv1  gate1234(.a(s_50), .O(gate259inter3));
  inv1  gate1235(.a(s_51), .O(gate259inter4));
  nand2 gate1236(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1237(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1238(.a(N1063), .O(gate259inter7));
  inv1  gate1239(.a(N1064), .O(gate259inter8));
  nand2 gate1240(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1241(.a(s_51), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1242(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1243(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1244(.a(gate259inter12), .b(gate259inter1), .O(N1158));
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );

  xor2  gate1959(.a(N938), .b(N1010), .O(gate271inter0));
  nand2 gate1960(.a(gate271inter0), .b(s_154), .O(gate271inter1));
  and2  gate1961(.a(N938), .b(N1010), .O(gate271inter2));
  inv1  gate1962(.a(s_154), .O(gate271inter3));
  inv1  gate1963(.a(s_155), .O(gate271inter4));
  nand2 gate1964(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1965(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1966(.a(N1010), .O(gate271inter7));
  inv1  gate1967(.a(N938), .O(gate271inter8));
  nand2 gate1968(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1969(.a(s_155), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1970(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1971(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1972(.a(gate271inter12), .b(gate271inter1), .O(N1206));
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate1413(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate1414(.a(gate273inter0), .b(s_76), .O(gate273inter1));
  and2  gate1415(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate1416(.a(s_76), .O(gate273inter3));
  inv1  gate1417(.a(s_77), .O(gate273inter4));
  nand2 gate1418(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1419(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1420(.a(N1013), .O(gate273inter7));
  inv1  gate1421(.a(N942), .O(gate273inter8));
  nand2 gate1422(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1423(.a(s_77), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1424(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1425(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1426(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate1777(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate1778(.a(gate275inter0), .b(s_128), .O(gate275inter1));
  and2  gate1779(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate1780(.a(s_128), .O(gate275inter3));
  inv1  gate1781(.a(s_129), .O(gate275inter4));
  nand2 gate1782(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1783(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1784(.a(N1016), .O(gate275inter7));
  inv1  gate1785(.a(N946), .O(gate275inter8));
  nand2 gate1786(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1787(.a(s_129), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1788(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1789(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1790(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate993(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate994(.a(gate277inter0), .b(s_16), .O(gate277inter1));
  and2  gate995(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate996(.a(s_16), .O(gate277inter3));
  inv1  gate997(.a(s_17), .O(gate277inter4));
  nand2 gate998(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate999(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1000(.a(N1019), .O(gate277inter7));
  inv1  gate1001(.a(N950), .O(gate277inter8));
  nand2 gate1002(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1003(.a(s_17), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1004(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1005(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1006(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );

  xor2  gate1399(.a(N954), .b(N1022), .O(gate279inter0));
  nand2 gate1400(.a(gate279inter0), .b(s_74), .O(gate279inter1));
  and2  gate1401(.a(N954), .b(N1022), .O(gate279inter2));
  inv1  gate1402(.a(s_74), .O(gate279inter3));
  inv1  gate1403(.a(s_75), .O(gate279inter4));
  nand2 gate1404(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1405(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1406(.a(N1022), .O(gate279inter7));
  inv1  gate1407(.a(N954), .O(gate279inter8));
  nand2 gate1408(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1409(.a(s_75), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1410(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1411(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1412(.a(gate279inter12), .b(gate279inter1), .O(N1214));
inv1 gate280( .a(N1025), .O(N1215) );

  xor2  gate1679(.a(N958), .b(N1025), .O(gate281inter0));
  nand2 gate1680(.a(gate281inter0), .b(s_114), .O(gate281inter1));
  and2  gate1681(.a(N958), .b(N1025), .O(gate281inter2));
  inv1  gate1682(.a(s_114), .O(gate281inter3));
  inv1  gate1683(.a(s_115), .O(gate281inter4));
  nand2 gate1684(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1685(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1686(.a(N1025), .O(gate281inter7));
  inv1  gate1687(.a(N958), .O(gate281inter8));
  nand2 gate1688(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1689(.a(s_115), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1690(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1691(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1692(.a(gate281inter12), .b(gate281inter1), .O(N1216));
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate1833(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate1834(.a(gate312inter0), .b(s_136), .O(gate312inter1));
  and2  gate1835(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate1836(.a(s_136), .O(gate312inter3));
  inv1  gate1837(.a(s_137), .O(gate312inter4));
  nand2 gate1838(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate1839(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate1840(.a(N631), .O(gate312inter7));
  inv1  gate1841(.a(N1159), .O(gate312inter8));
  nand2 gate1842(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate1843(.a(s_137), .b(gate312inter3), .O(gate312inter10));
  nor2  gate1844(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate1845(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate1846(.a(gate312inter12), .b(gate312inter1), .O(N1267));
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );

  xor2  gate1805(.a(N1207), .b(N691), .O(gate314inter0));
  nand2 gate1806(.a(gate314inter0), .b(s_132), .O(gate314inter1));
  and2  gate1807(.a(N1207), .b(N691), .O(gate314inter2));
  inv1  gate1808(.a(s_132), .O(gate314inter3));
  inv1  gate1809(.a(s_133), .O(gate314inter4));
  nand2 gate1810(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate1811(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate1812(.a(N691), .O(gate314inter7));
  inv1  gate1813(.a(N1207), .O(gate314inter8));
  nand2 gate1814(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate1815(.a(s_133), .b(gate314inter3), .O(gate314inter10));
  nor2  gate1816(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate1817(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate1818(.a(gate314inter12), .b(gate314inter1), .O(N1310));
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );

  xor2  gate2001(.a(N1215), .b(N703), .O(gate318inter0));
  nand2 gate2002(.a(gate318inter0), .b(s_160), .O(gate318inter1));
  and2  gate2003(.a(N1215), .b(N703), .O(gate318inter2));
  inv1  gate2004(.a(s_160), .O(gate318inter3));
  inv1  gate2005(.a(s_161), .O(gate318inter4));
  nand2 gate2006(.a(gate318inter4), .b(gate318inter3), .O(gate318inter5));
  nor2  gate2007(.a(gate318inter5), .b(gate318inter2), .O(gate318inter6));
  inv1  gate2008(.a(N703), .O(gate318inter7));
  inv1  gate2009(.a(N1215), .O(gate318inter8));
  nand2 gate2010(.a(gate318inter8), .b(gate318inter7), .O(gate318inter9));
  nand2 gate2011(.a(s_161), .b(gate318inter3), .O(gate318inter10));
  nor2  gate2012(.a(gate318inter10), .b(gate318inter9), .O(gate318inter11));
  nor2  gate2013(.a(gate318inter11), .b(gate318inter6), .O(gate318inter12));
  nand2 gate2014(.a(gate318inter12), .b(gate318inter1), .O(N1314));
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );

  xor2  gate1301(.a(N1223), .b(N709), .O(gate320inter0));
  nand2 gate1302(.a(gate320inter0), .b(s_60), .O(gate320inter1));
  and2  gate1303(.a(N1223), .b(N709), .O(gate320inter2));
  inv1  gate1304(.a(s_60), .O(gate320inter3));
  inv1  gate1305(.a(s_61), .O(gate320inter4));
  nand2 gate1306(.a(gate320inter4), .b(gate320inter3), .O(gate320inter5));
  nor2  gate1307(.a(gate320inter5), .b(gate320inter2), .O(gate320inter6));
  inv1  gate1308(.a(N709), .O(gate320inter7));
  inv1  gate1309(.a(N1223), .O(gate320inter8));
  nand2 gate1310(.a(gate320inter8), .b(gate320inter7), .O(gate320inter9));
  nand2 gate1311(.a(s_61), .b(gate320inter3), .O(gate320inter10));
  nor2  gate1312(.a(gate320inter10), .b(gate320inter9), .O(gate320inter11));
  nor2  gate1313(.a(gate320inter11), .b(gate320inter6), .O(gate320inter12));
  nand2 gate1314(.a(gate320inter12), .b(gate320inter1), .O(N1316));
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );

  xor2  gate1021(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate1022(.a(gate326inter0), .b(s_20), .O(gate326inter1));
  and2  gate1023(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate1024(.a(s_20), .O(gate326inter3));
  inv1  gate1025(.a(s_21), .O(gate326inter4));
  nand2 gate1026(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate1027(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate1028(.a(N733), .O(gate326inter7));
  inv1  gate1029(.a(N1241), .O(gate326inter8));
  nand2 gate1030(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate1031(.a(s_21), .b(gate326inter3), .O(gate326inter10));
  nor2  gate1032(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate1033(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate1034(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );

  xor2  gate1049(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate1050(.a(gate342inter0), .b(s_24), .O(gate342inter1));
  and2  gate1051(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate1052(.a(s_24), .O(gate342inter3));
  inv1  gate1053(.a(s_25), .O(gate342inter4));
  nand2 gate1054(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate1055(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate1056(.a(N1316), .O(gate342inter7));
  inv1  gate1057(.a(N1224), .O(gate342inter8));
  nand2 gate1058(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate1059(.a(s_25), .b(gate342inter3), .O(gate342inter10));
  nor2  gate1060(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate1061(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate1062(.a(gate342inter12), .b(gate342inter1), .O(N1373));
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );

  xor2  gate1539(.a(N1231), .b(N1322), .O(gate345inter0));
  nand2 gate1540(.a(gate345inter0), .b(s_94), .O(gate345inter1));
  and2  gate1541(.a(N1231), .b(N1322), .O(gate345inter2));
  inv1  gate1542(.a(s_94), .O(gate345inter3));
  inv1  gate1543(.a(s_95), .O(gate345inter4));
  nand2 gate1544(.a(gate345inter4), .b(gate345inter3), .O(gate345inter5));
  nor2  gate1545(.a(gate345inter5), .b(gate345inter2), .O(gate345inter6));
  inv1  gate1546(.a(N1322), .O(gate345inter7));
  inv1  gate1547(.a(N1231), .O(gate345inter8));
  nand2 gate1548(.a(gate345inter8), .b(gate345inter7), .O(gate345inter9));
  nand2 gate1549(.a(s_95), .b(gate345inter3), .O(gate345inter10));
  nor2  gate1550(.a(gate345inter10), .b(gate345inter9), .O(gate345inter11));
  nor2  gate1551(.a(gate345inter11), .b(gate345inter6), .O(gate345inter12));
  nand2 gate1552(.a(gate345inter12), .b(gate345inter1), .O(N1383));
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate937(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate938(.a(gate376inter0), .b(s_8), .O(gate376inter1));
  and2  gate939(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate940(.a(s_8), .O(gate376inter3));
  inv1  gate941(.a(s_9), .O(gate376inter4));
  nand2 gate942(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate943(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate944(.a(N1364), .O(gate376inter7));
  inv1  gate945(.a(N1154), .O(gate376inter8));
  nand2 gate946(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate947(.a(s_9), .b(gate376inter3), .O(gate376inter10));
  nor2  gate948(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate949(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate950(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );

  xor2  gate1987(.a(N1222), .b(N1370), .O(gate387inter0));
  nand2 gate1988(.a(gate387inter0), .b(s_158), .O(gate387inter1));
  and2  gate1989(.a(N1222), .b(N1370), .O(gate387inter2));
  inv1  gate1990(.a(s_158), .O(gate387inter3));
  inv1  gate1991(.a(s_159), .O(gate387inter4));
  nand2 gate1992(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1993(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1994(.a(N1370), .O(gate387inter7));
  inv1  gate1995(.a(N1222), .O(gate387inter8));
  nand2 gate1996(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1997(.a(s_159), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1998(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1999(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2000(.a(gate387inter12), .b(gate387inter1), .O(N1469));
inv1 gate388( .a(N1376), .O(N1470) );

  xor2  gate1889(.a(N1227), .b(N1376), .O(gate389inter0));
  nand2 gate1890(.a(gate389inter0), .b(s_144), .O(gate389inter1));
  and2  gate1891(.a(N1227), .b(N1376), .O(gate389inter2));
  inv1  gate1892(.a(s_144), .O(gate389inter3));
  inv1  gate1893(.a(s_145), .O(gate389inter4));
  nand2 gate1894(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1895(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1896(.a(N1376), .O(gate389inter7));
  inv1  gate1897(.a(N1227), .O(gate389inter8));
  nand2 gate1898(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1899(.a(s_145), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1900(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1901(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1902(.a(gate389inter12), .b(gate389inter1), .O(N1471));

  xor2  gate1595(.a(N1433), .b(N1387), .O(gate390inter0));
  nand2 gate1596(.a(gate390inter0), .b(s_102), .O(gate390inter1));
  and2  gate1597(.a(N1433), .b(N1387), .O(gate390inter2));
  inv1  gate1598(.a(s_102), .O(gate390inter3));
  inv1  gate1599(.a(s_103), .O(gate390inter4));
  nand2 gate1600(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1601(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1602(.a(N1387), .O(gate390inter7));
  inv1  gate1603(.a(N1433), .O(gate390inter8));
  nand2 gate1604(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1605(.a(s_103), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1606(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1607(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1608(.a(gate390inter12), .b(gate390inter1), .O(N1472));
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );

  xor2  gate1903(.a(N1448), .b(N943), .O(gate398inter0));
  nand2 gate1904(.a(gate398inter0), .b(s_146), .O(gate398inter1));
  and2  gate1905(.a(N1448), .b(N943), .O(gate398inter2));
  inv1  gate1906(.a(s_146), .O(gate398inter3));
  inv1  gate1907(.a(s_147), .O(gate398inter4));
  nand2 gate1908(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1909(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1910(.a(N943), .O(gate398inter7));
  inv1  gate1911(.a(N1448), .O(gate398inter8));
  nand2 gate1912(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1913(.a(s_147), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1914(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1915(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1916(.a(gate398inter12), .b(gate398inter1), .O(N1489));
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );

  xor2  gate1427(.a(N1452), .b(N947), .O(gate401inter0));
  nand2 gate1428(.a(gate401inter0), .b(s_78), .O(gate401inter1));
  and2  gate1429(.a(N1452), .b(N947), .O(gate401inter2));
  inv1  gate1430(.a(s_78), .O(gate401inter3));
  inv1  gate1431(.a(s_79), .O(gate401inter4));
  nand2 gate1432(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1433(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1434(.a(N947), .O(gate401inter7));
  inv1  gate1435(.a(N1452), .O(gate401inter8));
  nand2 gate1436(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1437(.a(s_79), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1438(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1439(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1440(.a(gate401inter12), .b(gate401inter1), .O(N1492));
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );

  xor2  gate1819(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate1820(.a(gate406inter0), .b(s_134), .O(gate406inter1));
  and2  gate1821(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate1822(.a(s_134), .O(gate406inter3));
  inv1  gate1823(.a(s_135), .O(gate406inter4));
  nand2 gate1824(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1825(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1826(.a(N998), .O(gate406inter7));
  inv1  gate1827(.a(N1463), .O(gate406inter8));
  nand2 gate1828(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1829(.a(s_135), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1830(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1831(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1832(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );

  xor2  gate1287(.a(N1470), .b(N973), .O(gate409inter0));
  nand2 gate1288(.a(gate409inter0), .b(s_58), .O(gate409inter1));
  and2  gate1289(.a(N1470), .b(N973), .O(gate409inter2));
  inv1  gate1290(.a(s_58), .O(gate409inter3));
  inv1  gate1291(.a(s_59), .O(gate409inter4));
  nand2 gate1292(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1293(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1294(.a(N973), .O(gate409inter7));
  inv1  gate1295(.a(N1470), .O(gate409inter8));
  nand2 gate1296(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1297(.a(s_59), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1298(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1299(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1300(.a(gate409inter12), .b(gate409inter1), .O(N1501));
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );

  xor2  gate1847(.a(N1489), .b(N1447), .O(gate414inter0));
  nand2 gate1848(.a(gate414inter0), .b(s_138), .O(gate414inter1));
  and2  gate1849(.a(N1489), .b(N1447), .O(gate414inter2));
  inv1  gate1850(.a(s_138), .O(gate414inter3));
  inv1  gate1851(.a(s_139), .O(gate414inter4));
  nand2 gate1852(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1853(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1854(.a(N1447), .O(gate414inter7));
  inv1  gate1855(.a(N1489), .O(gate414inter8));
  nand2 gate1856(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1857(.a(s_139), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1858(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1859(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1860(.a(gate414inter12), .b(gate414inter1), .O(N1517));
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );

  xor2  gate1371(.a(N1494), .b(N1455), .O(gate417inter0));
  nand2 gate1372(.a(gate417inter0), .b(s_70), .O(gate417inter1));
  and2  gate1373(.a(N1494), .b(N1455), .O(gate417inter2));
  inv1  gate1374(.a(s_70), .O(gate417inter3));
  inv1  gate1375(.a(s_71), .O(gate417inter4));
  nand2 gate1376(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1377(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1378(.a(N1455), .O(gate417inter7));
  inv1  gate1379(.a(N1494), .O(gate417inter8));
  nand2 gate1380(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1381(.a(s_71), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1382(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1383(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1384(.a(gate417inter12), .b(gate417inter1), .O(N1522));
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate1665(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate1666(.a(gate421inter0), .b(s_112), .O(gate421inter1));
  and2  gate1667(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate1668(.a(s_112), .O(gate421inter3));
  inv1  gate1669(.a(s_113), .O(gate421inter4));
  nand2 gate1670(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1671(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1672(.a(N1462), .O(gate421inter7));
  inv1  gate1673(.a(N1498), .O(gate421inter8));
  nand2 gate1674(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1675(.a(s_113), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1676(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1677(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1678(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );

  xor2  gate1441(.a(N1531), .b(N1484), .O(gate432inter0));
  nand2 gate1442(.a(gate432inter0), .b(s_80), .O(gate432inter1));
  and2  gate1443(.a(N1531), .b(N1484), .O(gate432inter2));
  inv1  gate1444(.a(s_80), .O(gate432inter3));
  inv1  gate1445(.a(s_81), .O(gate432inter4));
  nand2 gate1446(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1447(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1448(.a(N1484), .O(gate432inter7));
  inv1  gate1449(.a(N1531), .O(gate432inter8));
  nand2 gate1450(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1451(.a(s_81), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1452(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1453(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1454(.a(gate432inter12), .b(gate432inter1), .O(N1567));
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );

  xor2  gate1469(.a(N1569), .b(N1576), .O(gate453inter0));
  nand2 gate1470(.a(gate453inter0), .b(s_84), .O(gate453inter1));
  and2  gate1471(.a(N1569), .b(N1576), .O(gate453inter2));
  inv1  gate1472(.a(s_84), .O(gate453inter3));
  inv1  gate1473(.a(s_85), .O(gate453inter4));
  nand2 gate1474(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1475(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1476(.a(N1576), .O(gate453inter7));
  inv1  gate1477(.a(N1569), .O(gate453inter8));
  nand2 gate1478(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1479(.a(s_85), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1480(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1481(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1482(.a(gate453inter12), .b(gate453inter1), .O(N1638));
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );

  xor2  gate1091(.a(N1217), .b(N1606), .O(gate466inter0));
  nand2 gate1092(.a(gate466inter0), .b(s_30), .O(gate466inter1));
  and2  gate1093(.a(N1217), .b(N1606), .O(gate466inter2));
  inv1  gate1094(.a(s_30), .O(gate466inter3));
  inv1  gate1095(.a(s_31), .O(gate466inter4));
  nand2 gate1096(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1097(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1098(.a(N1606), .O(gate466inter7));
  inv1  gate1099(.a(N1217), .O(gate466inter8));
  nand2 gate1100(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1101(.a(s_31), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1102(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1103(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1104(.a(gate466inter12), .b(gate466inter1), .O(N1678));
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );

  xor2  gate1245(.a(N1675), .b(N1647), .O(gate478inter0));
  nand2 gate1246(.a(gate478inter0), .b(s_52), .O(gate478inter1));
  and2  gate1247(.a(N1675), .b(N1647), .O(gate478inter2));
  inv1  gate1248(.a(s_52), .O(gate478inter3));
  inv1  gate1249(.a(s_53), .O(gate478inter4));
  nand2 gate1250(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1251(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1252(.a(N1647), .O(gate478inter7));
  inv1  gate1253(.a(N1675), .O(gate478inter8));
  nand2 gate1254(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1255(.a(s_53), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1256(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1257(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1258(.a(gate478inter12), .b(gate478inter1), .O(N1708));
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );

  xor2  gate1861(.a(N1713), .b(N1680), .O(gate500inter0));
  nand2 gate1862(.a(gate500inter0), .b(s_140), .O(gate500inter1));
  and2  gate1863(.a(N1713), .b(N1680), .O(gate500inter2));
  inv1  gate1864(.a(s_140), .O(gate500inter3));
  inv1  gate1865(.a(s_141), .O(gate500inter4));
  nand2 gate1866(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1867(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1868(.a(N1680), .O(gate500inter7));
  inv1  gate1869(.a(N1713), .O(gate500inter8));
  nand2 gate1870(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1871(.a(s_141), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1872(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1873(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1874(.a(gate500inter12), .b(gate500inter1), .O(N1751));

  xor2  gate1707(.a(N1721), .b(N1537), .O(gate501inter0));
  nand2 gate1708(.a(gate501inter0), .b(s_118), .O(gate501inter1));
  and2  gate1709(.a(N1721), .b(N1537), .O(gate501inter2));
  inv1  gate1710(.a(s_118), .O(gate501inter3));
  inv1  gate1711(.a(s_119), .O(gate501inter4));
  nand2 gate1712(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1713(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1714(.a(N1537), .O(gate501inter7));
  inv1  gate1715(.a(N1721), .O(gate501inter8));
  nand2 gate1716(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1717(.a(s_119), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1718(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1719(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1720(.a(gate501inter12), .b(gate501inter1), .O(N1759));
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate1931(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate1932(.a(gate503inter0), .b(s_150), .O(gate503inter1));
  and2  gate1933(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate1934(.a(s_150), .O(gate503inter3));
  inv1  gate1935(.a(s_151), .O(gate503inter4));
  nand2 gate1936(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1937(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1938(.a(N1697), .O(gate503inter7));
  inv1  gate1939(.a(N1727), .O(gate503inter8));
  nand2 gate1940(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1941(.a(s_151), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1942(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1943(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1944(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );

  xor2  gate1189(.a(N1730), .b(N1701), .O(gate505inter0));
  nand2 gate1190(.a(gate505inter0), .b(s_44), .O(gate505inter1));
  and2  gate1191(.a(N1730), .b(N1701), .O(gate505inter2));
  inv1  gate1192(.a(s_44), .O(gate505inter3));
  inv1  gate1193(.a(s_45), .O(gate505inter4));
  nand2 gate1194(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1195(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1196(.a(N1701), .O(gate505inter7));
  inv1  gate1197(.a(N1730), .O(gate505inter8));
  nand2 gate1198(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1199(.a(s_45), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1200(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1201(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1202(.a(gate505inter12), .b(gate505inter1), .O(N1764));
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );

  xor2  gate1623(.a(N1763), .b(N1664), .O(gate519inter0));
  nand2 gate1624(.a(gate519inter0), .b(s_106), .O(gate519inter1));
  and2  gate1625(.a(N1763), .b(N1664), .O(gate519inter2));
  inv1  gate1626(.a(s_106), .O(gate519inter3));
  inv1  gate1627(.a(s_107), .O(gate519inter4));
  nand2 gate1628(.a(gate519inter4), .b(gate519inter3), .O(gate519inter5));
  nor2  gate1629(.a(gate519inter5), .b(gate519inter2), .O(gate519inter6));
  inv1  gate1630(.a(N1664), .O(gate519inter7));
  inv1  gate1631(.a(N1763), .O(gate519inter8));
  nand2 gate1632(.a(gate519inter8), .b(gate519inter7), .O(gate519inter9));
  nand2 gate1633(.a(s_107), .b(gate519inter3), .O(gate519inter10));
  nor2  gate1634(.a(gate519inter10), .b(gate519inter9), .O(gate519inter11));
  nor2  gate1635(.a(gate519inter11), .b(gate519inter6), .O(gate519inter12));
  nand2 gate1636(.a(gate519inter12), .b(gate519inter1), .O(N1792));

  xor2  gate1525(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate1526(.a(gate520inter0), .b(s_92), .O(gate520inter1));
  and2  gate1527(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate1528(.a(s_92), .O(gate520inter3));
  inv1  gate1529(.a(s_93), .O(gate520inter4));
  nand2 gate1530(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate1531(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate1532(.a(N1751), .O(gate520inter7));
  inv1  gate1533(.a(N1155), .O(gate520inter8));
  nand2 gate1534(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate1535(.a(s_93), .b(gate520inter3), .O(gate520inter10));
  nor2  gate1536(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate1537(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate1538(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );

  xor2  gate1105(.a(N1218), .b(N1748), .O(gate526inter0));
  nand2 gate1106(.a(gate526inter0), .b(s_32), .O(gate526inter1));
  and2  gate1107(.a(N1218), .b(N1748), .O(gate526inter2));
  inv1  gate1108(.a(s_32), .O(gate526inter3));
  inv1  gate1109(.a(s_33), .O(gate526inter4));
  nand2 gate1110(.a(gate526inter4), .b(gate526inter3), .O(gate526inter5));
  nor2  gate1111(.a(gate526inter5), .b(gate526inter2), .O(gate526inter6));
  inv1  gate1112(.a(N1748), .O(gate526inter7));
  inv1  gate1113(.a(N1218), .O(gate526inter8));
  nand2 gate1114(.a(gate526inter8), .b(gate526inter7), .O(gate526inter9));
  nand2 gate1115(.a(s_33), .b(gate526inter3), .O(gate526inter10));
  nor2  gate1116(.a(gate526inter10), .b(gate526inter9), .O(gate526inter11));
  nor2  gate1117(.a(gate526inter11), .b(gate526inter6), .O(gate526inter12));
  nand2 gate1118(.a(gate526inter12), .b(gate526inter1), .O(N1808));

  xor2  gate1511(.a(N1783), .b(N1612), .O(gate527inter0));
  nand2 gate1512(.a(gate527inter0), .b(s_90), .O(gate527inter1));
  and2  gate1513(.a(N1783), .b(N1612), .O(gate527inter2));
  inv1  gate1514(.a(s_90), .O(gate527inter3));
  inv1  gate1515(.a(s_91), .O(gate527inter4));
  nand2 gate1516(.a(gate527inter4), .b(gate527inter3), .O(gate527inter5));
  nor2  gate1517(.a(gate527inter5), .b(gate527inter2), .O(gate527inter6));
  inv1  gate1518(.a(N1612), .O(gate527inter7));
  inv1  gate1519(.a(N1783), .O(gate527inter8));
  nand2 gate1520(.a(gate527inter8), .b(gate527inter7), .O(gate527inter9));
  nand2 gate1521(.a(s_91), .b(gate527inter3), .O(gate527inter10));
  nor2  gate1522(.a(gate527inter10), .b(gate527inter9), .O(gate527inter11));
  nor2  gate1523(.a(gate527inter11), .b(gate527inter6), .O(gate527inter12));
  nand2 gate1524(.a(gate527inter12), .b(gate527inter1), .O(N1809));
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );

  xor2  gate1035(.a(N1801), .b(N1772), .O(gate539inter0));
  nand2 gate1036(.a(gate539inter0), .b(s_22), .O(gate539inter1));
  and2  gate1037(.a(N1801), .b(N1772), .O(gate539inter2));
  inv1  gate1038(.a(s_22), .O(gate539inter3));
  inv1  gate1039(.a(s_23), .O(gate539inter4));
  nand2 gate1040(.a(gate539inter4), .b(gate539inter3), .O(gate539inter5));
  nor2  gate1041(.a(gate539inter5), .b(gate539inter2), .O(gate539inter6));
  inv1  gate1042(.a(N1772), .O(gate539inter7));
  inv1  gate1043(.a(N1801), .O(gate539inter8));
  nand2 gate1044(.a(gate539inter8), .b(gate539inter7), .O(gate539inter9));
  nand2 gate1045(.a(s_23), .b(gate539inter3), .O(gate539inter10));
  nor2  gate1046(.a(gate539inter10), .b(gate539inter9), .O(gate539inter11));
  nor2  gate1047(.a(gate539inter11), .b(gate539inter6), .O(gate539inter12));
  nand2 gate1048(.a(gate539inter12), .b(gate539inter1), .O(N1830));
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );

  xor2  gate1553(.a(N1787), .b(N1810), .O(gate542inter0));
  nand2 gate1554(.a(gate542inter0), .b(s_96), .O(gate542inter1));
  and2  gate1555(.a(N1787), .b(N1810), .O(gate542inter2));
  inv1  gate1556(.a(s_96), .O(gate542inter3));
  inv1  gate1557(.a(s_97), .O(gate542inter4));
  nand2 gate1558(.a(gate542inter4), .b(gate542inter3), .O(gate542inter5));
  nor2  gate1559(.a(gate542inter5), .b(gate542inter2), .O(gate542inter6));
  inv1  gate1560(.a(N1810), .O(gate542inter7));
  inv1  gate1561(.a(N1787), .O(gate542inter8));
  nand2 gate1562(.a(gate542inter8), .b(gate542inter7), .O(gate542inter9));
  nand2 gate1563(.a(s_97), .b(gate542inter3), .O(gate542inter10));
  nor2  gate1564(.a(gate542inter10), .b(gate542inter9), .O(gate542inter11));
  nor2  gate1565(.a(gate542inter11), .b(gate542inter6), .O(gate542inter12));
  nand2 gate1566(.a(gate542inter12), .b(gate542inter1), .O(N1841));
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );

  xor2  gate1203(.a(N290), .b(N1798), .O(gate550inter0));
  nand2 gate1204(.a(gate550inter0), .b(s_46), .O(gate550inter1));
  and2  gate1205(.a(N290), .b(N1798), .O(gate550inter2));
  inv1  gate1206(.a(s_46), .O(gate550inter3));
  inv1  gate1207(.a(s_47), .O(gate550inter4));
  nand2 gate1208(.a(gate550inter4), .b(gate550inter3), .O(gate550inter5));
  nor2  gate1209(.a(gate550inter5), .b(gate550inter2), .O(gate550inter6));
  inv1  gate1210(.a(N1798), .O(gate550inter7));
  inv1  gate1211(.a(N290), .O(gate550inter8));
  nand2 gate1212(.a(gate550inter8), .b(gate550inter7), .O(gate550inter9));
  nand2 gate1213(.a(s_47), .b(gate550inter3), .O(gate550inter10));
  nor2  gate1214(.a(gate550inter10), .b(gate550inter9), .O(gate550inter11));
  nor2  gate1215(.a(gate550inter11), .b(gate550inter6), .O(gate550inter12));
  nand2 gate1216(.a(gate550inter12), .b(gate550inter1), .O(N1858));
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );

  xor2  gate1693(.a(N1848), .b(N1821), .O(gate557inter0));
  nand2 gate1694(.a(gate557inter0), .b(s_116), .O(gate557inter1));
  and2  gate1695(.a(N1848), .b(N1821), .O(gate557inter2));
  inv1  gate1696(.a(s_116), .O(gate557inter3));
  inv1  gate1697(.a(s_117), .O(gate557inter4));
  nand2 gate1698(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate1699(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate1700(.a(N1821), .O(gate557inter7));
  inv1  gate1701(.a(N1848), .O(gate557inter8));
  nand2 gate1702(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate1703(.a(s_117), .b(gate557inter3), .O(gate557inter10));
  nor2  gate1704(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate1705(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate1706(.a(gate557inter12), .b(gate557inter1), .O(N1878));
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );

  xor2  gate1329(.a(N1852), .b(N1826), .O(gate561inter0));
  nand2 gate1330(.a(gate561inter0), .b(s_64), .O(gate561inter1));
  and2  gate1331(.a(N1852), .b(N1826), .O(gate561inter2));
  inv1  gate1332(.a(s_64), .O(gate561inter3));
  inv1  gate1333(.a(s_65), .O(gate561inter4));
  nand2 gate1334(.a(gate561inter4), .b(gate561inter3), .O(gate561inter5));
  nor2  gate1335(.a(gate561inter5), .b(gate561inter2), .O(gate561inter6));
  inv1  gate1336(.a(N1826), .O(gate561inter7));
  inv1  gate1337(.a(N1852), .O(gate561inter8));
  nand2 gate1338(.a(gate561inter8), .b(gate561inter7), .O(gate561inter9));
  nand2 gate1339(.a(s_65), .b(gate561inter3), .O(gate561inter10));
  nor2  gate1340(.a(gate561inter10), .b(gate561inter9), .O(gate561inter11));
  nor2  gate1341(.a(gate561inter11), .b(gate561inter6), .O(gate561inter12));
  nand2 gate1342(.a(gate561inter12), .b(gate561inter1), .O(N1884));
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );

  xor2  gate1721(.a(N1885), .b(N1855), .O(gate572inter0));
  nand2 gate1722(.a(gate572inter0), .b(s_120), .O(gate572inter1));
  and2  gate1723(.a(N1885), .b(N1855), .O(gate572inter2));
  inv1  gate1724(.a(s_120), .O(gate572inter3));
  inv1  gate1725(.a(s_121), .O(gate572inter4));
  nand2 gate1726(.a(gate572inter4), .b(gate572inter3), .O(gate572inter5));
  nor2  gate1727(.a(gate572inter5), .b(gate572inter2), .O(gate572inter6));
  inv1  gate1728(.a(N1855), .O(gate572inter7));
  inv1  gate1729(.a(N1885), .O(gate572inter8));
  nand2 gate1730(.a(gate572inter8), .b(gate572inter7), .O(gate572inter9));
  nand2 gate1731(.a(s_121), .b(gate572inter3), .O(gate572inter10));
  nor2  gate1732(.a(gate572inter10), .b(gate572inter9), .O(gate572inter11));
  nor2  gate1733(.a(gate572inter11), .b(gate572inter6), .O(gate572inter12));
  nand2 gate1734(.a(gate572inter12), .b(gate572inter1), .O(N1913));
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate1119(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate1120(.a(gate596inter0), .b(s_34), .O(gate596inter1));
  and2  gate1121(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate1122(.a(s_34), .O(gate596inter3));
  inv1  gate1123(.a(s_35), .O(gate596inter4));
  nand2 gate1124(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate1125(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate1126(.a(N1930), .O(gate596inter7));
  inv1  gate1127(.a(N917), .O(gate596inter8));
  nand2 gate1128(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate1129(.a(s_35), .b(gate596inter3), .O(gate596inter10));
  nor2  gate1130(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate1131(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate1132(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );

  xor2  gate1875(.a(N918), .b(N1927), .O(gate598inter0));
  nand2 gate1876(.a(gate598inter0), .b(s_142), .O(gate598inter1));
  and2  gate1877(.a(N918), .b(N1927), .O(gate598inter2));
  inv1  gate1878(.a(s_142), .O(gate598inter3));
  inv1  gate1879(.a(s_143), .O(gate598inter4));
  nand2 gate1880(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate1881(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate1882(.a(N1927), .O(gate598inter7));
  inv1  gate1883(.a(N918), .O(gate598inter8));
  nand2 gate1884(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate1885(.a(s_143), .b(gate598inter3), .O(gate598inter10));
  nor2  gate1886(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate1887(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate1888(.a(gate598inter12), .b(gate598inter1), .O(N1977));
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );

  xor2  gate1357(.a(N1937), .b(N1944), .O(gate605inter0));
  nand2 gate1358(.a(gate605inter0), .b(s_68), .O(gate605inter1));
  and2  gate1359(.a(N1937), .b(N1944), .O(gate605inter2));
  inv1  gate1360(.a(s_68), .O(gate605inter3));
  inv1  gate1361(.a(s_69), .O(gate605inter4));
  nand2 gate1362(.a(gate605inter4), .b(gate605inter3), .O(gate605inter5));
  nor2  gate1363(.a(gate605inter5), .b(gate605inter2), .O(gate605inter6));
  inv1  gate1364(.a(N1944), .O(gate605inter7));
  inv1  gate1365(.a(N1937), .O(gate605inter8));
  nand2 gate1366(.a(gate605inter8), .b(gate605inter7), .O(gate605inter9));
  nand2 gate1367(.a(s_69), .b(gate605inter3), .O(gate605inter10));
  nor2  gate1368(.a(gate605inter10), .b(gate605inter9), .O(gate605inter11));
  nor2  gate1369(.a(gate605inter11), .b(gate605inter6), .O(gate605inter12));
  nand2 gate1370(.a(gate605inter12), .b(gate605inter1), .O(N2000));
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate1077(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate1078(.a(gate612inter0), .b(s_28), .O(gate612inter1));
  and2  gate1079(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate1080(.a(s_28), .O(gate612inter3));
  inv1  gate1081(.a(s_29), .O(gate612inter4));
  nand2 gate1082(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate1083(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate1084(.a(N673), .O(gate612inter7));
  inv1  gate1085(.a(N1976), .O(gate612inter8));
  nand2 gate1086(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate1087(.a(s_29), .b(gate612inter3), .O(gate612inter10));
  nor2  gate1088(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate1089(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate1090(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );

  xor2  gate1385(.a(N2013), .b(N1875), .O(gate631inter0));
  nand2 gate1386(.a(gate631inter0), .b(s_72), .O(gate631inter1));
  and2  gate1387(.a(N2013), .b(N1875), .O(gate631inter2));
  inv1  gate1388(.a(s_72), .O(gate631inter3));
  inv1  gate1389(.a(s_73), .O(gate631inter4));
  nand2 gate1390(.a(gate631inter4), .b(gate631inter3), .O(gate631inter5));
  nor2  gate1391(.a(gate631inter5), .b(gate631inter2), .O(gate631inter6));
  inv1  gate1392(.a(N1875), .O(gate631inter7));
  inv1  gate1393(.a(N2013), .O(gate631inter8));
  nand2 gate1394(.a(gate631inter8), .b(gate631inter7), .O(gate631inter9));
  nand2 gate1395(.a(s_73), .b(gate631inter3), .O(gate631inter10));
  nor2  gate1396(.a(gate631inter10), .b(gate631inter9), .O(gate631inter11));
  nor2  gate1397(.a(gate631inter11), .b(gate631inter6), .O(gate631inter12));
  nand2 gate1398(.a(gate631inter12), .b(gate631inter1), .O(N2036));

  xor2  gate1917(.a(N2015), .b(N1571), .O(gate632inter0));
  nand2 gate1918(.a(gate632inter0), .b(s_148), .O(gate632inter1));
  and2  gate1919(.a(N2015), .b(N1571), .O(gate632inter2));
  inv1  gate1920(.a(s_148), .O(gate632inter3));
  inv1  gate1921(.a(s_149), .O(gate632inter4));
  nand2 gate1922(.a(gate632inter4), .b(gate632inter3), .O(gate632inter5));
  nor2  gate1923(.a(gate632inter5), .b(gate632inter2), .O(gate632inter6));
  inv1  gate1924(.a(N1571), .O(gate632inter7));
  inv1  gate1925(.a(N2015), .O(gate632inter8));
  nand2 gate1926(.a(gate632inter8), .b(gate632inter7), .O(gate632inter9));
  nand2 gate1927(.a(s_149), .b(gate632inter3), .O(gate632inter10));
  nor2  gate1928(.a(gate632inter10), .b(gate632inter9), .O(gate632inter11));
  nor2  gate1929(.a(gate632inter11), .b(gate632inter6), .O(gate632inter12));
  nand2 gate1930(.a(gate632inter12), .b(gate632inter1), .O(N2037));
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );

  xor2  gate923(.a(N2024), .b(N2004), .O(gate636inter0));
  nand2 gate924(.a(gate636inter0), .b(s_6), .O(gate636inter1));
  and2  gate925(.a(N2024), .b(N2004), .O(gate636inter2));
  inv1  gate926(.a(s_6), .O(gate636inter3));
  inv1  gate927(.a(s_7), .O(gate636inter4));
  nand2 gate928(.a(gate636inter4), .b(gate636inter3), .O(gate636inter5));
  nor2  gate929(.a(gate636inter5), .b(gate636inter2), .O(gate636inter6));
  inv1  gate930(.a(N2004), .O(gate636inter7));
  inv1  gate931(.a(N2024), .O(gate636inter8));
  nand2 gate932(.a(gate636inter8), .b(gate636inter7), .O(gate636inter9));
  nand2 gate933(.a(s_7), .b(gate636inter3), .O(gate636inter10));
  nor2  gate934(.a(gate636inter10), .b(gate636inter9), .O(gate636inter11));
  nor2  gate935(.a(gate636inter11), .b(gate636inter6), .O(gate636inter12));
  nand2 gate936(.a(gate636inter12), .b(gate636inter1), .O(N2041));
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );

  xor2  gate1483(.a(N534), .b(N2558), .O(gate750inter0));
  nand2 gate1484(.a(gate750inter0), .b(s_86), .O(gate750inter1));
  and2  gate1485(.a(N534), .b(N2558), .O(gate750inter2));
  inv1  gate1486(.a(s_86), .O(gate750inter3));
  inv1  gate1487(.a(s_87), .O(gate750inter4));
  nand2 gate1488(.a(gate750inter4), .b(gate750inter3), .O(gate750inter5));
  nor2  gate1489(.a(gate750inter5), .b(gate750inter2), .O(gate750inter6));
  inv1  gate1490(.a(N2558), .O(gate750inter7));
  inv1  gate1491(.a(N534), .O(gate750inter8));
  nand2 gate1492(.a(gate750inter8), .b(gate750inter7), .O(gate750inter9));
  nand2 gate1493(.a(s_87), .b(gate750inter3), .O(gate750inter10));
  nor2  gate1494(.a(gate750inter10), .b(gate750inter9), .O(gate750inter11));
  nor2  gate1495(.a(gate750inter11), .b(gate750inter6), .O(gate750inter12));
  nand2 gate1496(.a(gate750inter12), .b(gate750inter1), .O(N2669));
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );

  xor2  gate1273(.a(N543), .b(N2570), .O(gate758inter0));
  nand2 gate1274(.a(gate758inter0), .b(s_56), .O(gate758inter1));
  and2  gate1275(.a(N543), .b(N2570), .O(gate758inter2));
  inv1  gate1276(.a(s_56), .O(gate758inter3));
  inv1  gate1277(.a(s_57), .O(gate758inter4));
  nand2 gate1278(.a(gate758inter4), .b(gate758inter3), .O(gate758inter5));
  nor2  gate1279(.a(gate758inter5), .b(gate758inter2), .O(gate758inter6));
  inv1  gate1280(.a(N2570), .O(gate758inter7));
  inv1  gate1281(.a(N543), .O(gate758inter8));
  nand2 gate1282(.a(gate758inter8), .b(gate758inter7), .O(gate758inter9));
  nand2 gate1283(.a(s_57), .b(gate758inter3), .O(gate758inter10));
  nor2  gate1284(.a(gate758inter10), .b(gate758inter9), .O(gate758inter11));
  nor2  gate1285(.a(gate758inter11), .b(gate758inter6), .O(gate758inter12));
  nand2 gate1286(.a(gate758inter12), .b(gate758inter1), .O(N2682));
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate1763(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate1764(.a(gate773inter0), .b(s_126), .O(gate773inter1));
  and2  gate1765(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate1766(.a(s_126), .O(gate773inter3));
  inv1  gate1767(.a(s_127), .O(gate773inter4));
  nand2 gate1768(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate1769(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate1770(.a(N2645), .O(gate773inter7));
  inv1  gate1771(.a(N540), .O(gate773inter8));
  nand2 gate1772(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate1773(.a(s_127), .b(gate773inter3), .O(gate773inter10));
  nor2  gate1774(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate1775(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate1776(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );

  xor2  gate1609(.a(N541), .b(N2648), .O(gate775inter0));
  nand2 gate1610(.a(gate775inter0), .b(s_104), .O(gate775inter1));
  and2  gate1611(.a(N541), .b(N2648), .O(gate775inter2));
  inv1  gate1612(.a(s_104), .O(gate775inter3));
  inv1  gate1613(.a(s_105), .O(gate775inter4));
  nand2 gate1614(.a(gate775inter4), .b(gate775inter3), .O(gate775inter5));
  nor2  gate1615(.a(gate775inter5), .b(gate775inter2), .O(gate775inter6));
  inv1  gate1616(.a(N2648), .O(gate775inter7));
  inv1  gate1617(.a(N541), .O(gate775inter8));
  nand2 gate1618(.a(gate775inter8), .b(gate775inter7), .O(gate775inter9));
  nand2 gate1619(.a(s_105), .b(gate775inter3), .O(gate775inter10));
  nor2  gate1620(.a(gate775inter10), .b(gate775inter9), .O(gate775inter11));
  nor2  gate1621(.a(gate775inter11), .b(gate775inter6), .O(gate775inter12));
  nand2 gate1622(.a(gate775inter12), .b(gate775inter1), .O(N2730));
inv1 gate776( .a(N2648), .O(N2731) );

  xor2  gate1791(.a(N542), .b(N2651), .O(gate777inter0));
  nand2 gate1792(.a(gate777inter0), .b(s_130), .O(gate777inter1));
  and2  gate1793(.a(N542), .b(N2651), .O(gate777inter2));
  inv1  gate1794(.a(s_130), .O(gate777inter3));
  inv1  gate1795(.a(s_131), .O(gate777inter4));
  nand2 gate1796(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate1797(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate1798(.a(N2651), .O(gate777inter7));
  inv1  gate1799(.a(N542), .O(gate777inter8));
  nand2 gate1800(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate1801(.a(s_131), .b(gate777inter3), .O(gate777inter10));
  nor2  gate1802(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate1803(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate1804(.a(gate777inter12), .b(gate777inter1), .O(N2732));
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );

  xor2  gate1133(.a(N2691), .b(N388), .O(gate789inter0));
  nand2 gate1134(.a(gate789inter0), .b(s_36), .O(gate789inter1));
  and2  gate1135(.a(N2691), .b(N388), .O(gate789inter2));
  inv1  gate1136(.a(s_36), .O(gate789inter3));
  inv1  gate1137(.a(s_37), .O(gate789inter4));
  nand2 gate1138(.a(gate789inter4), .b(gate789inter3), .O(gate789inter5));
  nor2  gate1139(.a(gate789inter5), .b(gate789inter2), .O(gate789inter6));
  inv1  gate1140(.a(N388), .O(gate789inter7));
  inv1  gate1141(.a(N2691), .O(gate789inter8));
  nand2 gate1142(.a(gate789inter8), .b(gate789inter7), .O(gate789inter9));
  nand2 gate1143(.a(s_37), .b(gate789inter3), .O(gate789inter10));
  nor2  gate1144(.a(gate789inter10), .b(gate789inter9), .O(gate789inter11));
  nor2  gate1145(.a(gate789inter11), .b(gate789inter6), .O(gate789inter12));
  nand2 gate1146(.a(gate789inter12), .b(gate789inter1), .O(N2744));
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );

  xor2  gate1735(.a(N2733), .b(N367), .O(gate802inter0));
  nand2 gate1736(.a(gate802inter0), .b(s_122), .O(gate802inter1));
  and2  gate1737(.a(N2733), .b(N367), .O(gate802inter2));
  inv1  gate1738(.a(s_122), .O(gate802inter3));
  inv1  gate1739(.a(s_123), .O(gate802inter4));
  nand2 gate1740(.a(gate802inter4), .b(gate802inter3), .O(gate802inter5));
  nor2  gate1741(.a(gate802inter5), .b(gate802inter2), .O(gate802inter6));
  inv1  gate1742(.a(N367), .O(gate802inter7));
  inv1  gate1743(.a(N2733), .O(gate802inter8));
  nand2 gate1744(.a(gate802inter8), .b(gate802inter7), .O(gate802inter9));
  nand2 gate1745(.a(s_123), .b(gate802inter3), .O(gate802inter10));
  nor2  gate1746(.a(gate802inter10), .b(gate802inter9), .O(gate802inter11));
  nor2  gate1747(.a(gate802inter11), .b(gate802inter6), .O(gate802inter12));
  nand2 gate1748(.a(gate802inter12), .b(gate802inter1), .O(N2761));

  xor2  gate979(.a(N2734), .b(N2682), .O(gate803inter0));
  nand2 gate980(.a(gate803inter0), .b(s_14), .O(gate803inter1));
  and2  gate981(.a(N2734), .b(N2682), .O(gate803inter2));
  inv1  gate982(.a(s_14), .O(gate803inter3));
  inv1  gate983(.a(s_15), .O(gate803inter4));
  nand2 gate984(.a(gate803inter4), .b(gate803inter3), .O(gate803inter5));
  nor2  gate985(.a(gate803inter5), .b(gate803inter2), .O(gate803inter6));
  inv1  gate986(.a(N2682), .O(gate803inter7));
  inv1  gate987(.a(N2734), .O(gate803inter8));
  nand2 gate988(.a(gate803inter8), .b(gate803inter7), .O(gate803inter9));
  nand2 gate989(.a(s_15), .b(gate803inter3), .O(gate803inter10));
  nor2  gate990(.a(gate803inter10), .b(gate803inter9), .O(gate803inter11));
  nor2  gate991(.a(gate803inter11), .b(gate803inter6), .O(gate803inter12));
  nand2 gate992(.a(gate803inter12), .b(gate803inter1), .O(N2762));
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );

  xor2  gate1455(.a(N2744), .b(N2690), .O(gate809inter0));
  nand2 gate1456(.a(gate809inter0), .b(s_82), .O(gate809inter1));
  and2  gate1457(.a(N2744), .b(N2690), .O(gate809inter2));
  inv1  gate1458(.a(s_82), .O(gate809inter3));
  inv1  gate1459(.a(s_83), .O(gate809inter4));
  nand2 gate1460(.a(gate809inter4), .b(gate809inter3), .O(gate809inter5));
  nor2  gate1461(.a(gate809inter5), .b(gate809inter2), .O(gate809inter6));
  inv1  gate1462(.a(N2690), .O(gate809inter7));
  inv1  gate1463(.a(N2744), .O(gate809inter8));
  nand2 gate1464(.a(gate809inter8), .b(gate809inter7), .O(gate809inter9));
  nand2 gate1465(.a(s_83), .b(gate809inter3), .O(gate809inter10));
  nor2  gate1466(.a(gate809inter10), .b(gate809inter9), .O(gate809inter11));
  nor2  gate1467(.a(gate809inter11), .b(gate809inter6), .O(gate809inter12));
  nand2 gate1468(.a(gate809inter12), .b(gate809inter1), .O(N2768));
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );

  xor2  gate951(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate952(.a(gate815inter0), .b(s_10), .O(gate815inter1));
  and2  gate953(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate954(.a(s_10), .O(gate815inter3));
  inv1  gate955(.a(s_11), .O(gate815inter4));
  nand2 gate956(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate957(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate958(.a(N2730), .O(gate815inter7));
  inv1  gate959(.a(N2760), .O(gate815inter8));
  nand2 gate960(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate961(.a(s_11), .b(gate815inter3), .O(gate815inter10));
  nor2  gate962(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate963(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate964(.a(gate815inter12), .b(gate815inter1), .O(N2782));
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );

  xor2  gate909(.a(N2765), .b(N2739), .O(gate819inter0));
  nand2 gate910(.a(gate819inter0), .b(s_4), .O(gate819inter1));
  and2  gate911(.a(N2765), .b(N2739), .O(gate819inter2));
  inv1  gate912(.a(s_4), .O(gate819inter3));
  inv1  gate913(.a(s_5), .O(gate819inter4));
  nand2 gate914(.a(gate819inter4), .b(gate819inter3), .O(gate819inter5));
  nor2  gate915(.a(gate819inter5), .b(gate819inter2), .O(gate819inter6));
  inv1  gate916(.a(N2739), .O(gate819inter7));
  inv1  gate917(.a(N2765), .O(gate819inter8));
  nand2 gate918(.a(gate819inter8), .b(gate819inter7), .O(gate819inter9));
  nand2 gate919(.a(s_5), .b(gate819inter3), .O(gate819inter10));
  nor2  gate920(.a(gate819inter10), .b(gate819inter9), .O(gate819inter11));
  nor2  gate921(.a(gate819inter11), .b(gate819inter6), .O(gate819inter12));
  nand2 gate922(.a(gate819inter12), .b(gate819inter1), .O(N2786));

  xor2  gate1343(.a(N2766), .b(N2741), .O(gate820inter0));
  nand2 gate1344(.a(gate820inter0), .b(s_66), .O(gate820inter1));
  and2  gate1345(.a(N2766), .b(N2741), .O(gate820inter2));
  inv1  gate1346(.a(s_66), .O(gate820inter3));
  inv1  gate1347(.a(s_67), .O(gate820inter4));
  nand2 gate1348(.a(gate820inter4), .b(gate820inter3), .O(gate820inter5));
  nor2  gate1349(.a(gate820inter5), .b(gate820inter2), .O(gate820inter6));
  inv1  gate1350(.a(N2741), .O(gate820inter7));
  inv1  gate1351(.a(N2766), .O(gate820inter8));
  nand2 gate1352(.a(gate820inter8), .b(gate820inter7), .O(gate820inter9));
  nand2 gate1353(.a(s_67), .b(gate820inter3), .O(gate820inter10));
  nor2  gate1354(.a(gate820inter10), .b(gate820inter9), .O(gate820inter11));
  nor2  gate1355(.a(gate820inter11), .b(gate820inter6), .O(gate820inter12));
  nand2 gate1356(.a(gate820inter12), .b(gate820inter1), .O(N2787));
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );

  xor2  gate1175(.a(N2800), .b(N2384), .O(gate828inter0));
  nand2 gate1176(.a(gate828inter0), .b(s_42), .O(gate828inter1));
  and2  gate1177(.a(N2800), .b(N2384), .O(gate828inter2));
  inv1  gate1178(.a(s_42), .O(gate828inter3));
  inv1  gate1179(.a(s_43), .O(gate828inter4));
  nand2 gate1180(.a(gate828inter4), .b(gate828inter3), .O(gate828inter5));
  nor2  gate1181(.a(gate828inter5), .b(gate828inter2), .O(gate828inter6));
  inv1  gate1182(.a(N2384), .O(gate828inter7));
  inv1  gate1183(.a(N2800), .O(gate828inter8));
  nand2 gate1184(.a(gate828inter8), .b(gate828inter7), .O(gate828inter9));
  nand2 gate1185(.a(s_43), .b(gate828inter3), .O(gate828inter10));
  nor2  gate1186(.a(gate828inter10), .b(gate828inter9), .O(gate828inter11));
  nor2  gate1187(.a(gate828inter11), .b(gate828inter6), .O(gate828inter12));
  nand2 gate1188(.a(gate828inter12), .b(gate828inter1), .O(N2811));
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );

  xor2  gate1567(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate1568(.a(gate840inter0), .b(s_98), .O(gate840inter1));
  and2  gate1569(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate1570(.a(s_98), .O(gate840inter3));
  inv1  gate1571(.a(s_99), .O(gate840inter4));
  nand2 gate1572(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate1573(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate1574(.a(N2815), .O(gate840inter7));
  inv1  gate1575(.a(N2077), .O(gate840inter8));
  nand2 gate1576(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate1577(.a(s_99), .b(gate840inter3), .O(gate840inter10));
  nor2  gate1578(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate1579(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate1580(.a(gate840inter12), .b(gate840inter1), .O(N2851));
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );

  xor2  gate1651(.a(N1985), .b(N2829), .O(gate850inter0));
  nand2 gate1652(.a(gate850inter0), .b(s_110), .O(gate850inter1));
  and2  gate1653(.a(N1985), .b(N2829), .O(gate850inter2));
  inv1  gate1654(.a(s_110), .O(gate850inter3));
  inv1  gate1655(.a(s_111), .O(gate850inter4));
  nand2 gate1656(.a(gate850inter4), .b(gate850inter3), .O(gate850inter5));
  nor2  gate1657(.a(gate850inter5), .b(gate850inter2), .O(gate850inter6));
  inv1  gate1658(.a(N2829), .O(gate850inter7));
  inv1  gate1659(.a(N1985), .O(gate850inter8));
  nand2 gate1660(.a(gate850inter8), .b(gate850inter7), .O(gate850inter9));
  nand2 gate1661(.a(s_111), .b(gate850inter3), .O(gate850inter10));
  nor2  gate1662(.a(gate850inter10), .b(gate850inter9), .O(gate850inter11));
  nor2  gate1663(.a(gate850inter11), .b(gate850inter6), .O(gate850inter12));
  nand2 gate1664(.a(gate850inter12), .b(gate850inter1), .O(N2863));
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );

  xor2  gate1315(.a(N2860), .b(N1818), .O(gate854inter0));
  nand2 gate1316(.a(gate854inter0), .b(s_62), .O(gate854inter1));
  and2  gate1317(.a(N2860), .b(N1818), .O(gate854inter2));
  inv1  gate1318(.a(s_62), .O(gate854inter3));
  inv1  gate1319(.a(s_63), .O(gate854inter4));
  nand2 gate1320(.a(gate854inter4), .b(gate854inter3), .O(gate854inter5));
  nor2  gate1321(.a(gate854inter5), .b(gate854inter2), .O(gate854inter6));
  inv1  gate1322(.a(N1818), .O(gate854inter7));
  inv1  gate1323(.a(N2860), .O(gate854inter8));
  nand2 gate1324(.a(gate854inter8), .b(gate854inter7), .O(gate854inter9));
  nand2 gate1325(.a(s_63), .b(gate854inter3), .O(gate854inter10));
  nor2  gate1326(.a(gate854inter10), .b(gate854inter9), .O(gate854inter11));
  nor2  gate1327(.a(gate854inter11), .b(gate854inter6), .O(gate854inter12));
  nand2 gate1328(.a(gate854inter12), .b(gate854inter1), .O(N2869));
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );

  xor2  gate1007(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1008(.a(gate856inter0), .b(s_18), .O(gate856inter1));
  and2  gate1009(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1010(.a(s_18), .O(gate856inter3));
  inv1  gate1011(.a(s_19), .O(gate856inter4));
  nand2 gate1012(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1013(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1014(.a(N2843), .O(gate856inter7));
  inv1  gate1015(.a(N886), .O(gate856inter8));
  nand2 gate1016(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1017(.a(s_19), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1018(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1019(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1020(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );

  xor2  gate881(.a(N887), .b(N2846), .O(gate858inter0));
  nand2 gate882(.a(gate858inter0), .b(s_0), .O(gate858inter1));
  and2  gate883(.a(N887), .b(N2846), .O(gate858inter2));
  inv1  gate884(.a(s_0), .O(gate858inter3));
  inv1  gate885(.a(s_1), .O(gate858inter4));
  nand2 gate886(.a(gate858inter4), .b(gate858inter3), .O(gate858inter5));
  nor2  gate887(.a(gate858inter5), .b(gate858inter2), .O(gate858inter6));
  inv1  gate888(.a(N2846), .O(gate858inter7));
  inv1  gate889(.a(N887), .O(gate858inter8));
  nand2 gate890(.a(gate858inter8), .b(gate858inter7), .O(gate858inter9));
  nand2 gate891(.a(s_1), .b(gate858inter3), .O(gate858inter10));
  nor2  gate892(.a(gate858inter10), .b(gate858inter9), .O(gate858inter11));
  nor2  gate893(.a(gate858inter11), .b(gate858inter6), .O(gate858inter12));
  nand2 gate894(.a(gate858inter12), .b(gate858inter1), .O(N2873));
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );

  xor2  gate1637(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate1638(.a(gate865inter0), .b(s_108), .O(gate865inter1));
  and2  gate1639(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate1640(.a(s_108), .O(gate865inter3));
  inv1  gate1641(.a(s_109), .O(gate865inter4));
  nand2 gate1642(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate1643(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate1644(.a(N2870), .O(gate865inter7));
  inv1  gate1645(.a(N2854), .O(gate865inter8));
  nand2 gate1646(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate1647(.a(s_109), .b(gate865inter3), .O(gate865inter10));
  nor2  gate1648(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate1649(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate1650(.a(gate865inter12), .b(gate865inter1), .O(N2880));
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );

  xor2  gate1497(.a(N2874), .b(N685), .O(gate867inter0));
  nand2 gate1498(.a(gate867inter0), .b(s_88), .O(gate867inter1));
  and2  gate1499(.a(N2874), .b(N685), .O(gate867inter2));
  inv1  gate1500(.a(s_88), .O(gate867inter3));
  inv1  gate1501(.a(s_89), .O(gate867inter4));
  nand2 gate1502(.a(gate867inter4), .b(gate867inter3), .O(gate867inter5));
  nor2  gate1503(.a(gate867inter5), .b(gate867inter2), .O(gate867inter6));
  inv1  gate1504(.a(N685), .O(gate867inter7));
  inv1  gate1505(.a(N2874), .O(gate867inter8));
  nand2 gate1506(.a(gate867inter8), .b(gate867inter7), .O(gate867inter9));
  nand2 gate1507(.a(s_89), .b(gate867inter3), .O(gate867inter10));
  nor2  gate1508(.a(gate867inter10), .b(gate867inter9), .O(gate867inter11));
  nor2  gate1509(.a(gate867inter11), .b(gate867inter6), .O(gate867inter12));
  nand2 gate1510(.a(gate867inter12), .b(gate867inter1), .O(N2882));
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );

  xor2  gate895(.a(N2882), .b(N2873), .O(gate875inter0));
  nand2 gate896(.a(gate875inter0), .b(s_2), .O(gate875inter1));
  and2  gate897(.a(N2882), .b(N2873), .O(gate875inter2));
  inv1  gate898(.a(s_2), .O(gate875inter3));
  inv1  gate899(.a(s_3), .O(gate875inter4));
  nand2 gate900(.a(gate875inter4), .b(gate875inter3), .O(gate875inter5));
  nor2  gate901(.a(gate875inter5), .b(gate875inter2), .O(gate875inter6));
  inv1  gate902(.a(N2873), .O(gate875inter7));
  inv1  gate903(.a(N2882), .O(gate875inter8));
  nand2 gate904(.a(gate875inter8), .b(gate875inter7), .O(gate875inter9));
  nand2 gate905(.a(s_3), .b(gate875inter3), .O(gate875inter10));
  nor2  gate906(.a(gate875inter10), .b(gate875inter9), .O(gate875inter11));
  nor2  gate907(.a(gate875inter11), .b(gate875inter6), .O(gate875inter12));
  nand2 gate908(.a(gate875inter12), .b(gate875inter1), .O(N2892));

  xor2  gate1259(.a(N1461), .b(N2883), .O(gate876inter0));
  nand2 gate1260(.a(gate876inter0), .b(s_54), .O(gate876inter1));
  and2  gate1261(.a(N1461), .b(N2883), .O(gate876inter2));
  inv1  gate1262(.a(s_54), .O(gate876inter3));
  inv1  gate1263(.a(s_55), .O(gate876inter4));
  nand2 gate1264(.a(gate876inter4), .b(gate876inter3), .O(gate876inter5));
  nor2  gate1265(.a(gate876inter5), .b(gate876inter2), .O(gate876inter6));
  inv1  gate1266(.a(N2883), .O(gate876inter7));
  inv1  gate1267(.a(N1461), .O(gate876inter8));
  nand2 gate1268(.a(gate876inter8), .b(gate876inter7), .O(gate876inter9));
  nand2 gate1269(.a(s_55), .b(gate876inter3), .O(gate876inter10));
  nor2  gate1270(.a(gate876inter10), .b(gate876inter9), .O(gate876inter11));
  nor2  gate1271(.a(gate876inter11), .b(gate876inter6), .O(gate876inter12));
  nand2 gate1272(.a(gate876inter12), .b(gate876inter1), .O(N2895));
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule