module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate245(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate246(.a(gate19inter0), .b(s_12), .O(gate19inter1));
  and2  gate247(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate248(.a(s_12), .O(gate19inter3));
  inv1  gate249(.a(s_13), .O(gate19inter4));
  nand2 gate250(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate251(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate252(.a(N118), .O(gate19inter7));
  inv1  gate253(.a(N4), .O(gate19inter8));
  nand2 gate254(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate255(.a(s_13), .b(gate19inter3), .O(gate19inter10));
  nor2  gate256(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate257(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate258(.a(gate19inter12), .b(gate19inter1), .O(N154));
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate273(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate274(.a(gate22inter0), .b(s_16), .O(gate22inter1));
  and2  gate275(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate276(.a(s_16), .O(gate22inter3));
  inv1  gate277(.a(s_17), .O(gate22inter4));
  nand2 gate278(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate279(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate280(.a(N122), .O(gate22inter7));
  inv1  gate281(.a(N17), .O(gate22inter8));
  nand2 gate282(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate283(.a(s_17), .b(gate22inter3), .O(gate22inter10));
  nor2  gate284(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate285(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate286(.a(gate22inter12), .b(gate22inter1), .O(N159));

  xor2  gate399(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate400(.a(gate23inter0), .b(s_34), .O(gate23inter1));
  and2  gate401(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate402(.a(s_34), .O(gate23inter3));
  inv1  gate403(.a(s_35), .O(gate23inter4));
  nand2 gate404(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate405(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate406(.a(N126), .O(gate23inter7));
  inv1  gate407(.a(N30), .O(gate23inter8));
  nand2 gate408(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate409(.a(s_35), .b(gate23inter3), .O(gate23inter10));
  nor2  gate410(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate411(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate412(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate189(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate190(.a(gate27inter0), .b(s_4), .O(gate27inter1));
  and2  gate191(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate192(.a(s_4), .O(gate27inter3));
  inv1  gate193(.a(s_5), .O(gate27inter4));
  nand2 gate194(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate195(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate196(.a(N142), .O(gate27inter7));
  inv1  gate197(.a(N82), .O(gate27inter8));
  nand2 gate198(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate199(.a(s_5), .b(gate27inter3), .O(gate27inter10));
  nor2  gate200(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate201(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate202(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate525(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate526(.a(gate32inter0), .b(s_52), .O(gate32inter1));
  and2  gate527(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate528(.a(s_52), .O(gate32inter3));
  inv1  gate529(.a(s_53), .O(gate32inter4));
  nand2 gate530(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate531(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate532(.a(N34), .O(gate32inter7));
  inv1  gate533(.a(N127), .O(gate32inter8));
  nand2 gate534(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate535(.a(s_53), .b(gate32inter3), .O(gate32inter10));
  nor2  gate536(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate537(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate538(.a(gate32inter12), .b(gate32inter1), .O(N185));

  xor2  gate357(.a(N127), .b(N40), .O(gate33inter0));
  nand2 gate358(.a(gate33inter0), .b(s_28), .O(gate33inter1));
  and2  gate359(.a(N127), .b(N40), .O(gate33inter2));
  inv1  gate360(.a(s_28), .O(gate33inter3));
  inv1  gate361(.a(s_29), .O(gate33inter4));
  nand2 gate362(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate363(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate364(.a(N40), .O(gate33inter7));
  inv1  gate365(.a(N127), .O(gate33inter8));
  nand2 gate366(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate367(.a(s_29), .b(gate33inter3), .O(gate33inter10));
  nor2  gate368(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate369(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate370(.a(gate33inter12), .b(gate33inter1), .O(N186));
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate231(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate232(.a(gate36inter0), .b(s_10), .O(gate36inter1));
  and2  gate233(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate234(.a(s_10), .O(gate36inter3));
  inv1  gate235(.a(s_11), .O(gate36inter4));
  nand2 gate236(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate237(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate238(.a(N60), .O(gate36inter7));
  inv1  gate239(.a(N135), .O(gate36inter8));
  nand2 gate240(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate241(.a(s_11), .b(gate36inter3), .O(gate36inter10));
  nor2  gate242(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate243(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate244(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );

  xor2  gate161(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate162(.a(gate39inter0), .b(s_0), .O(gate39inter1));
  and2  gate163(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate164(.a(s_0), .O(gate39inter3));
  inv1  gate165(.a(s_1), .O(gate39inter4));
  nand2 gate166(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate167(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate168(.a(N79), .O(gate39inter7));
  inv1  gate169(.a(N139), .O(gate39inter8));
  nand2 gate170(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate171(.a(s_1), .b(gate39inter3), .O(gate39inter10));
  nor2  gate172(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate173(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate174(.a(gate39inter12), .b(gate39inter1), .O(N192));
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );

  xor2  gate371(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate372(.a(gate53inter0), .b(s_30), .O(gate53inter1));
  and2  gate373(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate374(.a(s_30), .O(gate53inter3));
  inv1  gate375(.a(s_31), .O(gate53inter4));
  nand2 gate376(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate377(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate378(.a(N203), .O(gate53inter7));
  inv1  gate379(.a(N165), .O(gate53inter8));
  nand2 gate380(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate381(.a(s_31), .b(gate53inter3), .O(gate53inter10));
  nor2  gate382(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate383(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate384(.a(gate53inter12), .b(gate53inter1), .O(N233));
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );

  xor2  gate329(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate330(.a(gate56inter0), .b(s_24), .O(gate56inter1));
  and2  gate331(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate332(.a(s_24), .O(gate56inter3));
  inv1  gate333(.a(s_25), .O(gate56inter4));
  nand2 gate334(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate335(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate336(.a(N1), .O(gate56inter7));
  inv1  gate337(.a(N213), .O(gate56inter8));
  nand2 gate338(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate339(.a(s_25), .b(gate56inter3), .O(gate56inter10));
  nor2  gate340(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate341(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate342(.a(gate56inter12), .b(gate56inter1), .O(N242));
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate511(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate512(.a(gate62inter0), .b(s_50), .O(gate62inter1));
  and2  gate513(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate514(.a(s_50), .O(gate62inter3));
  inv1  gate515(.a(s_51), .O(gate62inter4));
  nand2 gate516(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate517(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate518(.a(N213), .O(gate62inter7));
  inv1  gate519(.a(N37), .O(gate62inter8));
  nand2 gate520(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate521(.a(s_51), .b(gate62inter3), .O(gate62inter10));
  nor2  gate522(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate523(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate524(.a(gate62inter12), .b(gate62inter1), .O(N254));
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );

  xor2  gate441(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate442(.a(gate66inter0), .b(s_40), .O(gate66inter1));
  and2  gate443(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate444(.a(s_40), .O(gate66inter3));
  inv1  gate445(.a(s_41), .O(gate66inter4));
  nand2 gate446(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate447(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate448(.a(N213), .O(gate66inter7));
  inv1  gate449(.a(N89), .O(gate66inter8));
  nand2 gate450(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate451(.a(s_41), .b(gate66inter3), .O(gate66inter10));
  nor2  gate452(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate453(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate454(.a(gate66inter12), .b(gate66inter1), .O(N258));

  xor2  gate581(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate582(.a(gate67inter0), .b(s_60), .O(gate67inter1));
  and2  gate583(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate584(.a(s_60), .O(gate67inter3));
  inv1  gate585(.a(s_61), .O(gate67inter4));
  nand2 gate586(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate587(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate588(.a(N213), .O(gate67inter7));
  inv1  gate589(.a(N102), .O(gate67inter8));
  nand2 gate590(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate591(.a(s_61), .b(gate67inter3), .O(gate67inter10));
  nor2  gate592(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate593(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate594(.a(gate67inter12), .b(gate67inter1), .O(N259));
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate385(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate386(.a(gate70inter0), .b(s_32), .O(gate70inter1));
  and2  gate387(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate388(.a(s_32), .O(gate70inter3));
  inv1  gate389(.a(s_33), .O(gate70inter4));
  nand2 gate390(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate391(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate392(.a(N227), .O(gate70inter7));
  inv1  gate393(.a(N183), .O(gate70inter8));
  nand2 gate394(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate395(.a(s_33), .b(gate70inter3), .O(gate70inter10));
  nor2  gate396(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate397(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate398(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate427(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate428(.a(gate72inter0), .b(s_38), .O(gate72inter1));
  and2  gate429(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate430(.a(s_38), .O(gate72inter3));
  inv1  gate431(.a(s_39), .O(gate72inter4));
  nand2 gate432(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate433(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate434(.a(N233), .O(gate72inter7));
  inv1  gate435(.a(N187), .O(gate72inter8));
  nand2 gate436(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate437(.a(s_39), .b(gate72inter3), .O(gate72inter10));
  nor2  gate438(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate439(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate440(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate343(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate344(.a(gate77inter0), .b(s_26), .O(gate77inter1));
  and2  gate345(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate346(.a(s_26), .O(gate77inter3));
  inv1  gate347(.a(s_27), .O(gate77inter4));
  nand2 gate348(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate349(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate350(.a(N251), .O(gate77inter7));
  inv1  gate351(.a(N197), .O(gate77inter8));
  nand2 gate352(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate353(.a(s_27), .b(gate77inter3), .O(gate77inter10));
  nor2  gate354(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate355(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate356(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate469(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate470(.a(gate80inter0), .b(s_44), .O(gate80inter1));
  and2  gate471(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate472(.a(s_44), .O(gate80inter3));
  inv1  gate473(.a(s_45), .O(gate80inter4));
  nand2 gate474(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate475(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate476(.a(N233), .O(gate80inter7));
  inv1  gate477(.a(N188), .O(gate80inter8));
  nand2 gate478(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate479(.a(s_45), .b(gate80inter3), .O(gate80inter10));
  nor2  gate480(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate481(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate482(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );

  xor2  gate287(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate288(.a(gate84inter0), .b(s_18), .O(gate84inter1));
  and2  gate289(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate290(.a(s_18), .O(gate84inter3));
  inv1  gate291(.a(s_19), .O(gate84inter4));
  nand2 gate292(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate293(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate294(.a(N247), .O(gate84inter7));
  inv1  gate295(.a(N196), .O(gate84inter8));
  nand2 gate296(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate297(.a(s_19), .b(gate84inter3), .O(gate84inter10));
  nor2  gate298(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate299(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate300(.a(gate84inter12), .b(gate84inter1), .O(N294));
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate483(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate484(.a(gate99inter0), .b(s_46), .O(gate99inter1));
  and2  gate485(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate486(.a(s_46), .O(gate99inter3));
  inv1  gate487(.a(s_47), .O(gate99inter4));
  nand2 gate488(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate489(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate490(.a(N309), .O(gate99inter7));
  inv1  gate491(.a(N260), .O(gate99inter8));
  nand2 gate492(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate493(.a(s_47), .b(gate99inter3), .O(gate99inter10));
  nor2  gate494(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate495(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate496(.a(gate99inter12), .b(gate99inter1), .O(N330));

  xor2  gate497(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate498(.a(gate100inter0), .b(s_48), .O(gate100inter1));
  and2  gate499(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate500(.a(s_48), .O(gate100inter3));
  inv1  gate501(.a(s_49), .O(gate100inter4));
  nand2 gate502(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate503(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate504(.a(N309), .O(gate100inter7));
  inv1  gate505(.a(N264), .O(gate100inter8));
  nand2 gate506(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate507(.a(s_49), .b(gate100inter3), .O(gate100inter10));
  nor2  gate508(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate509(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate510(.a(gate100inter12), .b(gate100inter1), .O(N331));
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );

  xor2  gate413(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate414(.a(gate106inter0), .b(s_36), .O(gate106inter1));
  and2  gate415(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate416(.a(s_36), .O(gate106inter3));
  inv1  gate417(.a(s_37), .O(gate106inter4));
  nand2 gate418(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate419(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate420(.a(N309), .O(gate106inter7));
  inv1  gate421(.a(N276), .O(gate106inter8));
  nand2 gate422(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate423(.a(s_37), .b(gate106inter3), .O(gate106inter10));
  nor2  gate424(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate425(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate426(.a(gate106inter12), .b(gate106inter1), .O(N337));

  xor2  gate217(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate218(.a(gate107inter0), .b(s_8), .O(gate107inter1));
  and2  gate219(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate220(.a(s_8), .O(gate107inter3));
  inv1  gate221(.a(s_9), .O(gate107inter4));
  nand2 gate222(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate223(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate224(.a(N319), .O(gate107inter7));
  inv1  gate225(.a(N34), .O(gate107inter8));
  nand2 gate226(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate227(.a(s_9), .b(gate107inter3), .O(gate107inter10));
  nor2  gate228(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate229(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate230(.a(gate107inter12), .b(gate107inter1), .O(N338));

  xor2  gate539(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate540(.a(gate108inter0), .b(s_54), .O(gate108inter1));
  and2  gate541(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate542(.a(s_54), .O(gate108inter3));
  inv1  gate543(.a(s_55), .O(gate108inter4));
  nand2 gate544(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate545(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate546(.a(N309), .O(gate108inter7));
  inv1  gate547(.a(N279), .O(gate108inter8));
  nand2 gate548(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate549(.a(s_55), .b(gate108inter3), .O(gate108inter10));
  nor2  gate550(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate551(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate552(.a(gate108inter12), .b(gate108inter1), .O(N339));
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate315(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate316(.a(gate111inter0), .b(s_22), .O(gate111inter1));
  and2  gate317(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate318(.a(s_22), .O(gate111inter3));
  inv1  gate319(.a(s_23), .O(gate111inter4));
  nand2 gate320(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate321(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate322(.a(N319), .O(gate111inter7));
  inv1  gate323(.a(N60), .O(gate111inter8));
  nand2 gate324(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate325(.a(s_23), .b(gate111inter3), .O(gate111inter10));
  nor2  gate326(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate327(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate328(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate175(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate176(.a(gate113inter0), .b(s_2), .O(gate113inter1));
  and2  gate177(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate178(.a(s_2), .O(gate113inter3));
  inv1  gate179(.a(s_3), .O(gate113inter4));
  nand2 gate180(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate181(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate182(.a(N319), .O(gate113inter7));
  inv1  gate183(.a(N73), .O(gate113inter8));
  nand2 gate184(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate185(.a(s_3), .b(gate113inter3), .O(gate113inter10));
  nor2  gate186(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate187(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate188(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate259(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate260(.a(gate119inter0), .b(s_14), .O(gate119inter1));
  and2  gate261(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate262(.a(s_14), .O(gate119inter3));
  inv1  gate263(.a(s_15), .O(gate119inter4));
  nand2 gate264(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate265(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate266(.a(N332), .O(gate119inter7));
  inv1  gate267(.a(N302), .O(gate119inter8));
  nand2 gate268(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate269(.a(s_15), .b(gate119inter3), .O(gate119inter10));
  nor2  gate270(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate271(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate272(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate567(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate568(.a(gate121inter0), .b(s_58), .O(gate121inter1));
  and2  gate569(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate570(.a(s_58), .O(gate121inter3));
  inv1  gate571(.a(s_59), .O(gate121inter4));
  nand2 gate572(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate573(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate574(.a(N335), .O(gate121inter7));
  inv1  gate575(.a(N304), .O(gate121inter8));
  nand2 gate576(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate577(.a(s_59), .b(gate121inter3), .O(gate121inter10));
  nor2  gate578(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate579(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate580(.a(gate121inter12), .b(gate121inter1), .O(N352));
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );

  xor2  gate203(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate204(.a(gate125inter0), .b(s_6), .O(gate125inter1));
  and2  gate205(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate206(.a(s_6), .O(gate125inter3));
  inv1  gate207(.a(s_7), .O(gate125inter4));
  nand2 gate208(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate209(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate210(.a(N343), .O(gate125inter7));
  inv1  gate211(.a(N308), .O(gate125inter8));
  nand2 gate212(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate213(.a(s_7), .b(gate125inter3), .O(gate125inter10));
  nor2  gate214(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate215(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate216(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate553(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate554(.a(gate131inter0), .b(s_56), .O(gate131inter1));
  and2  gate555(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate556(.a(s_56), .O(gate131inter3));
  inv1  gate557(.a(s_57), .O(gate131inter4));
  nand2 gate558(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate559(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate560(.a(N360), .O(gate131inter7));
  inv1  gate561(.a(N40), .O(gate131inter8));
  nand2 gate562(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate563(.a(s_57), .b(gate131inter3), .O(gate131inter10));
  nor2  gate564(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate565(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate566(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );

  xor2  gate301(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate302(.a(gate133inter0), .b(s_20), .O(gate133inter1));
  and2  gate303(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate304(.a(s_20), .O(gate133inter3));
  inv1  gate305(.a(s_21), .O(gate133inter4));
  nand2 gate306(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate307(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate308(.a(N360), .O(gate133inter7));
  inv1  gate309(.a(N66), .O(gate133inter8));
  nand2 gate310(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate311(.a(s_21), .b(gate133inter3), .O(gate133inter10));
  nor2  gate312(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate313(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate314(.a(gate133inter12), .b(gate133inter1), .O(N375));
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate455(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate456(.a(gate135inter0), .b(s_42), .O(gate135inter1));
  and2  gate457(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate458(.a(s_42), .O(gate135inter3));
  inv1  gate459(.a(s_43), .O(gate135inter4));
  nand2 gate460(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate461(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate462(.a(N360), .O(gate135inter7));
  inv1  gate463(.a(N92), .O(gate135inter8));
  nand2 gate464(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate465(.a(s_43), .b(gate135inter3), .O(gate135inter10));
  nor2  gate466(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate467(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate468(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule