module c5315 (N1,N4,N11,N14,N17,N20,N23,N24,N25,N26,
              N27,N31,N34,N37,N40,N43,N46,N49,N52,N53,
              N54,N61,N64,N67,N70,N73,N76,N79,N80,N81,
              N82,N83,N86,N87,N88,N91,N94,N97,N100,N103,
              N106,N109,N112,N113,N114,N115,N116,N117,N118,N119,
              N120,N121,N122,N123,N126,N127,N128,N129,N130,N131,
              N132,N135,N136,N137,N140,N141,N145,N146,N149,N152,
              N155,N158,N161,N164,N167,N170,N173,N176,N179,N182,
              N185,N188,N191,N194,N197,N200,N203,N206,N209,N210,
              N217,N218,N225,N226,N233,N234,N241,N242,N245,N248,
              N251,N254,N257,N264,N265,N272,N273,N280,N281,N288,
              N289,N292,N293,N299,N302,N307,N308,N315,N316,N323,
              N324,N331,N332,N335,N338,N341,N348,N351,N358,N361,
              N366,N369,N372,N373,N374,N386,N389,N400,N411,N422,
              N435,N446,N457,N468,N479,N490,N503,N514,N523,N534,
              N545,N549,N552,N556,N559,N562,N566,N571,N574,N577,
              N580,N583,N588,N591,N592,N595,N596,N597,N598,N599,
              N603,N607,N610,N613,N616,N619,N625,N631,N709,N816,
              N1066,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,
              N1147,N1152,N1153,N1154,N1155,N1972,N2054,N2060,N2061,N2139,
              N2142,N2309,N2387,N2527,N2584,N2590,N2623,N3357,N3358,N3359,
              N3360,N3604,N3613,N4272,N4275,N4278,N4279,N4737,N4738,N4739,
              N4740,N5240,N5388,N6641,N6643,N6646,N6648,N6716,N6877,N6924,
              N6925,N6926,N6927,N7015,N7363,N7365,N7432,N7449,N7465,N7466,
              N7467,N7469,N7470,N7471,N7472,N7473,N7474,N7476,N7503,N7504,
              N7506,N7511,N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,
              N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7626,N7698,
              N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7735,
              N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7754,N7755,N7756,
              N7757,N7758,N7759,N7760,N7761,N8075,N8076,N8123,N8124,N8127,
              N8128);

input N1,N4,N11,N14,N17,N20,N23,N24,N25,N26,
      N27,N31,N34,N37,N40,N43,N46,N49,N52,N53,
      N54,N61,N64,N67,N70,N73,N76,N79,N80,N81,
      N82,N83,N86,N87,N88,N91,N94,N97,N100,N103,
      N106,N109,N112,N113,N114,N115,N116,N117,N118,N119,
      N120,N121,N122,N123,N126,N127,N128,N129,N130,N131,
      N132,N135,N136,N137,N140,N141,N145,N146,N149,N152,
      N155,N158,N161,N164,N167,N170,N173,N176,N179,N182,
      N185,N188,N191,N194,N197,N200,N203,N206,N209,N210,
      N217,N218,N225,N226,N233,N234,N241,N242,N245,N248,
      N251,N254,N257,N264,N265,N272,N273,N280,N281,N288,
      N289,N292,N293,N299,N302,N307,N308,N315,N316,N323,
      N324,N331,N332,N335,N338,N341,N348,N351,N358,N361,
      N366,N369,N372,N373,N374,N386,N389,N400,N411,N422,
      N435,N446,N457,N468,N479,N490,N503,N514,N523,N534,
      N545,N549,N552,N556,N559,N562,N566,N571,N574,N577,
      N580,N583,N588,N591,N592,N595,N596,N597,N598,N599,
      N603,N607,N610,N613,N616,N619,N625,N631;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
output N709,N816,N1066,N1137,N1138,N1139,N1140,N1141,N1142,N1143,
       N1144,N1145,N1147,N1152,N1153,N1154,N1155,N1972,N2054,N2060,
       N2061,N2139,N2142,N2309,N2387,N2527,N2584,N2590,N2623,N3357,
       N3358,N3359,N3360,N3604,N3613,N4272,N4275,N4278,N4279,N4737,
       N4738,N4739,N4740,N5240,N5388,N6641,N6643,N6646,N6648,N6716,
       N6877,N6924,N6925,N6926,N6927,N7015,N7363,N7365,N7432,N7449,
       N7465,N7466,N7467,N7469,N7470,N7471,N7472,N7473,N7474,N7476,
       N7503,N7504,N7506,N7511,N7515,N7516,N7517,N7518,N7519,N7520,
       N7521,N7522,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,
       N7626,N7698,N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,
       N7707,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7754,
       N7755,N7756,N7757,N7758,N7759,N7760,N7761,N8075,N8076,N8123,
       N8124,N8127,N8128;

wire N1042,N1043,N1067,N1080,N1092,N1104,N1146,N1148,N1149,N1150,
     N1151,N1156,N1157,N1161,N1173,N1185,N1197,N1209,N1213,N1216,
     N1219,N1223,N1235,N1247,N1259,N1271,N1280,N1292,N1303,N1315,
     N1327,N1339,N1351,N1363,N1375,N1378,N1381,N1384,N1387,N1390,
     N1393,N1396,N1415,N1418,N1421,N1424,N1427,N1430,N1433,N1436,
     N1455,N1462,N1469,N1475,N1479,N1482,N1492,N1495,N1498,N1501,
     N1504,N1507,N1510,N1513,N1516,N1519,N1522,N1525,N1542,N1545,
     N1548,N1551,N1554,N1557,N1560,N1563,N1566,N1573,N1580,N1583,
     N1588,N1594,N1597,N1600,N1603,N1606,N1609,N1612,N1615,N1618,
     N1621,N1624,N1627,N1630,N1633,N1636,N1639,N1642,N1645,N1648,
     N1651,N1654,N1657,N1660,N1663,N1675,N1685,N1697,N1709,N1721,
     N1727,N1731,N1743,N1755,N1758,N1761,N1769,N1777,N1785,N1793,
     N1800,N1807,N1814,N1821,N1824,N1827,N1830,N1833,N1836,N1839,
     N1842,N1845,N1848,N1851,N1854,N1857,N1860,N1863,N1866,N1869,
     N1872,N1875,N1878,N1881,N1884,N1887,N1890,N1893,N1896,N1899,
     N1902,N1905,N1908,N1911,N1914,N1917,N1920,N1923,N1926,N1929,
     N1932,N1935,N1938,N1941,N1944,N1947,N1950,N1953,N1956,N1959,
     N1962,N1965,N1968,N2349,N2350,N2585,N2586,N2587,N2588,N2589,
     N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,
     N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
     N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,
     N2621,N2622,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,
     N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,
     N2642,N2643,N2644,N2645,N2646,N2647,N2653,N2664,N2675,N2681,
     N2692,N2703,N2704,N2709,N2710,N2711,N2712,N2713,N2714,N2715,
     N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2728,N2739,N2750,
     N2756,N2767,N2778,N2779,N2790,N2801,N2812,N2823,N2824,N2825,
     N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,
     N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,
     N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,
     N2861,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,
     N2876,N2877,N2882,N2891,N2901,N2902,N2903,N2904,N2905,N2906,
     N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,
     N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,
     N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,
     N2937,N2938,N2939,N2940,N2941,N2942,N2948,N2954,N2955,N2956,
     N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2969,N2970,
     N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,
     N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,
     N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,
     N3003,N3006,N3007,N3010,N3013,N3014,N3015,N3016,N3017,N3018,
     N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,
     N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3038,N3041,N3052,
     N3063,N3068,N3071,N3072,N3073,N3074,N3075,N3086,N3097,N3108,
     N3119,N3130,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3158,
     N3169,N3180,N3191,N3194,N3195,N3196,N3197,N3198,N3199,N3200,
     N3203,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,
     N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3444,N3445,N3446,
     N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,
     N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3481,N3482,
     N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,
     N3493,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,
     N3511,N3512,N3513,N3514,N3515,N3558,N3559,N3560,N3561,N3562,
     N3563,N3605,N3606,N3607,N3608,N3609,N3610,N3614,N3615,N3616,
     N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,
     N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,
     N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,
     N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,
     N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,
     N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,
     N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,
     N3687,N3688,N3689,N3691,N3700,N3701,N3702,N3703,N3704,N3705,
     N3708,N3709,N3710,N3711,N3712,N3713,N3715,N3716,N3717,N3718,
     N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,
     N3729,N3730,N3731,N3732,N3738,N3739,N3740,N3741,N3742,N3743,
     N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,
     N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,
     N3764,N3765,N3766,N3767,N3768,N3769,N3770,N3771,N3775,N3779,
     N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,
     N3793,N3797,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,
     N3808,N3809,N3810,N3813,N3816,N3819,N3822,N3823,N3824,N3827,
     N3828,N3829,N3830,N3831,N3834,N3835,N3836,N3837,N3838,N3839,
     N3840,N3841,N3842,N3849,N3855,N3861,N3867,N3873,N3881,N3887,
     N3893,N3908,N3909,N3911,N3914,N3915,N3916,N3917,N3918,N3919,
     N3920,N3921,N3927,N3933,N3942,N3948,N3956,N3962,N3968,N3975,
     N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,N3987,
     N3988,N3989,N3990,N3991,N3998,N4008,N4011,N4021,N4024,N4027,
     N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,
     N4041,N4042,N4067,N4080,N4088,N4091,N4094,N4097,N4100,N4103,
     N4106,N4109,N4144,N4147,N4150,N4153,N4156,N4159,N4183,N4184,
     N4185,N4186,N4188,N4191,N4196,N4197,N4198,N4199,N4200,N4203,
     N4206,N4209,N4212,N4215,N4219,N4223,N4224,N4225,N4228,N4231,
     N4234,N4237,N4240,N4243,N4246,N4249,N4252,N4255,N4258,N4263,
     N4264,N4267,N4268,N4269,N4270,N4271,N4273,N4274,N4276,N4277,
     N4280,N4284,N4290,N4297,N4298,N4301,N4305,N4310,N4316,N4320,
     N4325,N4331,N4332,N4336,N4342,N4349,N4357,N4364,N4375,N4379,
     N4385,N4392,N4396,N4400,N4405,N4412,N4418,N4425,N4436,N4440,
     N4445,N4451,N4456,N4462,N4469,N4477,N4512,N4515,N4516,N4521,
     N4523,N4524,N4532,N4547,N4548,N4551,N4554,N4557,N4560,N4563,
     N4566,N4569,N4572,N4575,N4578,N4581,N4584,N4587,N4590,N4593,
     N4596,N4599,N4602,N4605,N4608,N4611,N4614,N4617,N4621,N4624,
     N4627,N4630,N4633,N4637,N4640,N4643,N4646,N4649,N4652,N4655,
     N4658,N4662,N4665,N4668,N4671,N4674,N4677,N4680,N4683,N4686,
     N4689,N4692,N4695,N4698,N4701,N4702,N4720,N4721,N4724,N4725,
     N4726,N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,
     N4736,N4741,N4855,N4856,N4908,N4909,N4939,N4942,N4947,N4953,
     N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4965,N4966,
     N4967,N4968,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,
     N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N5049,N5052,
     N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,
     N5063,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,
     N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,
     N5084,N5085,N5086,N5087,N5088,N5089,N5090,N5091,N5092,N5093,
     N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,
     N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,
     N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,
     N5124,N5125,N5126,N5127,N5128,N5129,N5130,N5131,N5132,N5133,
     N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,N5144,
     N5145,N5146,N5147,N5148,N5150,N5153,N5154,N5155,N5156,N5157,
     N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5169,N5172,N5173,
     N5176,N5177,N5180,N5183,N5186,N5189,N5192,N5195,N5198,N5199,
     N5202,N5205,N5208,N5211,N5214,N5217,N5220,N5223,N5224,N5225,
     N5226,N5227,N5228,N5229,N5230,N5232,N5233,N5234,N5235,N5236,
     N5239,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,
     N5250,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,
     N5261,N5262,N5263,N5264,N5274,N5275,N5282,N5283,N5284,N5298,
     N5299,N5300,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,
     N5311,N5312,N5315,N5319,N5324,N5328,N5331,N5332,N5346,N5363,
     N5364,N5365,N5366,N5367,N5368,N5369,N5370,N5371,N5374,N5377,
     N5382,N5385,N5389,N5396,N5407,N5418,N5424,N5431,N5441,N5452,
     N5462,N5469,N5470,N5477,N5488,N5498,N5506,N5520,N5536,N5549,
     N5555,N5562,N5573,N5579,N5595,N5606,N5616,N5617,N5618,N5619,
     N5620,N5621,N5622,N5624,N5634,N5655,N5671,N5684,N5690,N5691,
     N5692,N5696,N5700,N5703,N5707,N5711,N5726,N5727,N5728,N5730,
     N5731,N5732,N5733,N5734,N5735,N5736,N5739,N5742,N5745,N5755,
     N5756,N5954,N5955,N5956,N6005,N6006,N6023,N6024,N6025,N6028,
     N6031,N6034,N6037,N6040,N6044,N6045,N6048,N6051,N6054,N6065,
     N6066,N6067,N6068,N6069,N6071,N6072,N6073,N6074,N6075,N6076,
     N6077,N6078,N6079,N6080,N6083,N6084,N6085,N6086,N6087,N6088,
     N6089,N6090,N6091,N6094,N6095,N6096,N6097,N6098,N6099,N6100,
     N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6111,N6112,
     N6113,N6114,N6115,N6116,N6117,N6120,N6121,N6122,N6123,N6124,
     N6125,N6126,N6127,N6128,N6129,N6130,N6131,N6132,N6133,N6134,
     N6135,N6136,N6137,N6138,N6139,N6140,N6143,N6144,N6145,N6146,
     N6147,N6148,N6149,N6152,N6153,N6154,N6155,N6156,N6157,N6158,
     N6159,N6160,N6161,N6162,N6163,N6164,N6168,N6171,N6172,N6173,
     N6174,N6175,N6178,N6179,N6180,N6181,N6182,N6183,N6184,N6185,
     N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6197,
     N6200,N6203,N6206,N6209,N6212,N6215,N6218,N6221,N6234,N6235,
     N6238,N6241,N6244,N6247,N6250,N6253,N6256,N6259,N6262,N6265,
     N6268,N6271,N6274,N6277,N6280,N6283,N6286,N6289,N6292,N6295,
     N6298,N6301,N6304,N6307,N6310,N6313,N6316,N6319,N6322,N6325,
     N6328,N6331,N6335,N6338,N6341,N6344,N6347,N6350,N6353,N6356,
     N6359,N6364,N6367,N6370,N6373,N6374,N6375,N6376,N6377,N6378,
     N6382,N6386,N6388,N6392,N6397,N6411,N6415,N6419,N6427,N6434,
     N6437,N6441,N6445,N6448,N6449,N6466,N6469,N6470,N6471,N6472,
     N6473,N6474,N6475,N6476,N6477,N6478,N6482,N6486,N6490,N6494,
     N6500,N6504,N6508,N6512,N6516,N6526,N6536,N6539,N6553,N6556,
     N6566,N6569,N6572,N6575,N6580,N6584,N6587,N6592,N6599,N6606,
     N6609,N6619,N6622,N6630,N6631,N6632,N6633,N6634,N6637,N6640,
     N6650,N6651,N6653,N6655,N6657,N6659,N6660,N6661,N6662,N6663,
     N6664,N6666,N6668,N6670,N6672,N6675,N6680,N6681,N6682,N6683,
     N6689,N6690,N6691,N6692,N6693,N6695,N6698,N6699,N6700,N6703,
     N6708,N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6718,N6719,
     N6720,N6721,N6722,N6724,N6739,N6740,N6741,N6744,N6745,N6746,
     N6751,N6752,N6753,N6754,N6755,N6760,N6761,N6762,N6772,N6773,
     N6776,N6777,N6782,N6783,N6784,N6785,N6790,N6791,N6792,N6795,
     N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,N6810,
     N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6823,N6824,N6825,
     N6826,N6827,N6828,N6829,N6830,N6831,N6834,N6835,N6836,N6837,
     N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6850,N6851,N6852,
     N6853,N6854,N6855,N6856,N6857,N6860,N6861,N6862,N6863,N6866,
     N6872,N6873,N6874,N6875,N6876,N6879,N6880,N6881,N6884,N6885,
     N6888,N6889,N6890,N6891,N6894,N6895,N6896,N6897,N6900,N6901,
     N6904,N6905,N6908,N6909,N6912,N6913,N6914,N6915,N6916,N6919,
     N6922,N6923,N6930,N6932,N6935,N6936,N6937,N6938,N6939,N6940,
     N6946,N6947,N6948,N6949,N6953,N6954,N6955,N6956,N6957,N6958,
     N6964,N6965,N6966,N6967,N6973,N6974,N6975,N6976,N6977,N6978,
     N6979,N6987,N6990,N6999,N7002,N7003,N7006,N7011,N7012,N7013,
     N7016,N7018,N7019,N7020,N7021,N7022,N7023,N7028,N7031,N7034,
     N7037,N7040,N7041,N7044,N7045,N7046,N7047,N7048,N7049,N7054,
     N7057,N7060,N7064,N7065,N7072,N7073,N7074,N7075,N7076,N7079,
     N7080,N7083,N7084,N7085,N7086,N7087,N7088,N7089,N7090,N7093,
     N7094,N7097,N7101,N7105,N7110,N7114,N7115,N7116,N7125,N7126,
     N7127,N7130,N7131,N7139,N7140,N7141,N7146,N7147,N7149,N7150,
     N7151,N7152,N7153,N7158,N7159,N7160,N7166,N7167,N7168,N7169,
     N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,
     N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,N7189,
     N7190,N7196,N7197,N7198,N7204,N7205,N7206,N7207,N7208,N7209,
     N7212,N7215,N7216,N7217,N7218,N7219,N7222,N7225,N7228,N7229,
     N7236,N7239,N7242,N7245,N7250,N7257,N7260,N7263,N7268,N7269,
     N7270,N7276,N7282,N7288,N7294,N7300,N7301,N7304,N7310,N7320,
     N7321,N7328,N7338,N7339,N7340,N7341,N7342,N7349,N7357,N7364,
     N7394,N7397,N7402,N7405,N7406,N7407,N7408,N7409,N7412,N7415,
     N7416,N7417,N7418,N7419,N7420,N7421,N7424,N7425,N7426,N7427,
     N7428,N7429,N7430,N7431,N7433,N7434,N7435,N7436,N7437,N7438,
     N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,
     N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,
     N7460,N7461,N7462,N7463,N7464,N7468,N7479,N7481,N7482,N7483,
     N7484,N7485,N7486,N7487,N7488,N7489,N7492,N7493,N7498,N7499,
     N7500,N7505,N7507,N7508,N7509,N7510,N7512,N7513,N7514,N7525,
     N7526,N7527,N7528,N7529,N7530,N7531,N7537,N7543,N7549,N7555,
     N7561,N7567,N7573,N7579,N7582,N7585,N7586,N7587,N7588,N7589,
     N7592,N7595,N7598,N7599,N7624,N7625,N7631,N7636,N7657,N7658,
     N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,N7674,
     N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,
     N7685,N7686,N7687,N7688,N7689,N7690,N7691,N7692,N7693,N7694,
     N7695,N7696,N7697,N7708,N7709,N7710,N7711,N7712,N7715,N7718,
     N7719,N7720,N7721,N7722,N7723,N7724,N7727,N7728,N7729,N7730,
     N7731,N7732,N7733,N7734,N7743,N7744,N7749,N7750,N7751,N7762,
     N7765,N7768,N7769,N7770,N7771,N7772,N7775,N7778,N7781,N7782,
     N7787,N7788,N7795,N7796,N7797,N7798,N7799,N7800,N7803,N7806,
     N7807,N7808,N7809,N7810,N7811,N7812,N7815,N7816,N7821,N7822,
     N7823,N7826,N7829,N7832,N7833,N7834,N7835,N7836,N7839,N7842,
     N7845,N7846,N7851,N7852,N7859,N7860,N7861,N7862,N7863,N7864,
     N7867,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7879,N7880,
     N7885,N7886,N7887,N7890,N7893,N7896,N7897,N7898,N7899,N7900,
     N7903,N7906,N7909,N7910,N7917,N7918,N7923,N7924,N7925,N7926,
     N7927,N7928,N7929,N7930,N7931,N7932,N7935,N7938,N7939,N7940,
     N7943,N7944,N7945,N7946,N7951,N7954,N7957,N7960,N7963,N7966,
     N7967,N7968,N7969,N7970,N7973,N7974,N7984,N7985,N7987,N7988,
     N7989,N7990,N7991,N7992,N7993,N7994,N7995,N7996,N7997,N7998,
     N8001,N8004,N8009,N8013,N8017,N8020,N8021,N8022,N8023,N8025,
     N8026,N8027,N8031,N8032,N8033,N8034,N8035,N8036,N8037,N8038,
     N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8048,N8055,N8056,
     N8057,N8058,N8059,N8060,N8061,N8064,N8071,N8072,N8073,N8074,
     N8077,N8078,N8079,N8082,N8089,N8090,N8091,N8092,N8093,N8096,
     N8099,N8102,N8113,N8114,N8115,N8116,N8117,N8118,N8119,N8120,
     N8121,N8122,N8125,N8126, gate1401inter0, gate1401inter1, gate1401inter2, gate1401inter3, gate1401inter4, gate1401inter5, gate1401inter6, gate1401inter7, gate1401inter8, gate1401inter9, gate1401inter10, gate1401inter11, gate1401inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate555inter0, gate555inter1, gate555inter2, gate555inter3, gate555inter4, gate555inter5, gate555inter6, gate555inter7, gate555inter8, gate555inter9, gate555inter10, gate555inter11, gate555inter12, gate1650inter0, gate1650inter1, gate1650inter2, gate1650inter3, gate1650inter4, gate1650inter5, gate1650inter6, gate1650inter7, gate1650inter8, gate1650inter9, gate1650inter10, gate1650inter11, gate1650inter12, gate2249inter0, gate2249inter1, gate2249inter2, gate2249inter3, gate2249inter4, gate2249inter5, gate2249inter6, gate2249inter7, gate2249inter8, gate2249inter9, gate2249inter10, gate2249inter11, gate2249inter12, gate1087inter0, gate1087inter1, gate1087inter2, gate1087inter3, gate1087inter4, gate1087inter5, gate1087inter6, gate1087inter7, gate1087inter8, gate1087inter9, gate1087inter10, gate1087inter11, gate1087inter12, gate1720inter0, gate1720inter1, gate1720inter2, gate1720inter3, gate1720inter4, gate1720inter5, gate1720inter6, gate1720inter7, gate1720inter8, gate1720inter9, gate1720inter10, gate1720inter11, gate1720inter12, gate2216inter0, gate2216inter1, gate2216inter2, gate2216inter3, gate2216inter4, gate2216inter5, gate2216inter6, gate2216inter7, gate2216inter8, gate2216inter9, gate2216inter10, gate2216inter11, gate2216inter12, gate1130inter0, gate1130inter1, gate1130inter2, gate1130inter3, gate1130inter4, gate1130inter5, gate1130inter6, gate1130inter7, gate1130inter8, gate1130inter9, gate1130inter10, gate1130inter11, gate1130inter12, gate2032inter0, gate2032inter1, gate2032inter2, gate2032inter3, gate2032inter4, gate2032inter5, gate2032inter6, gate2032inter7, gate2032inter8, gate2032inter9, gate2032inter10, gate2032inter11, gate2032inter12, gate2226inter0, gate2226inter1, gate2226inter2, gate2226inter3, gate2226inter4, gate2226inter5, gate2226inter6, gate2226inter7, gate2226inter8, gate2226inter9, gate2226inter10, gate2226inter11, gate2226inter12, gate1968inter0, gate1968inter1, gate1968inter2, gate1968inter3, gate1968inter4, gate1968inter5, gate1968inter6, gate1968inter7, gate1968inter8, gate1968inter9, gate1968inter10, gate1968inter11, gate1968inter12, gate1219inter0, gate1219inter1, gate1219inter2, gate1219inter3, gate1219inter4, gate1219inter5, gate1219inter6, gate1219inter7, gate1219inter8, gate1219inter9, gate1219inter10, gate1219inter11, gate1219inter12, gate977inter0, gate977inter1, gate977inter2, gate977inter3, gate977inter4, gate977inter5, gate977inter6, gate977inter7, gate977inter8, gate977inter9, gate977inter10, gate977inter11, gate977inter12, gate1716inter0, gate1716inter1, gate1716inter2, gate1716inter3, gate1716inter4, gate1716inter5, gate1716inter6, gate1716inter7, gate1716inter8, gate1716inter9, gate1716inter10, gate1716inter11, gate1716inter12, gate1296inter0, gate1296inter1, gate1296inter2, gate1296inter3, gate1296inter4, gate1296inter5, gate1296inter6, gate1296inter7, gate1296inter8, gate1296inter9, gate1296inter10, gate1296inter11, gate1296inter12, gate2140inter0, gate2140inter1, gate2140inter2, gate2140inter3, gate2140inter4, gate2140inter5, gate2140inter6, gate2140inter7, gate2140inter8, gate2140inter9, gate2140inter10, gate2140inter11, gate2140inter12, gate1721inter0, gate1721inter1, gate1721inter2, gate1721inter3, gate1721inter4, gate1721inter5, gate1721inter6, gate1721inter7, gate1721inter8, gate1721inter9, gate1721inter10, gate1721inter11, gate1721inter12, gate1179inter0, gate1179inter1, gate1179inter2, gate1179inter3, gate1179inter4, gate1179inter5, gate1179inter6, gate1179inter7, gate1179inter8, gate1179inter9, gate1179inter10, gate1179inter11, gate1179inter12, gate2200inter0, gate2200inter1, gate2200inter2, gate2200inter3, gate2200inter4, gate2200inter5, gate2200inter6, gate2200inter7, gate2200inter8, gate2200inter9, gate2200inter10, gate2200inter11, gate2200inter12, gate1872inter0, gate1872inter1, gate1872inter2, gate1872inter3, gate1872inter4, gate1872inter5, gate1872inter6, gate1872inter7, gate1872inter8, gate1872inter9, gate1872inter10, gate1872inter11, gate1872inter12, gate1757inter0, gate1757inter1, gate1757inter2, gate1757inter3, gate1757inter4, gate1757inter5, gate1757inter6, gate1757inter7, gate1757inter8, gate1757inter9, gate1757inter10, gate1757inter11, gate1757inter12, gate1213inter0, gate1213inter1, gate1213inter2, gate1213inter3, gate1213inter4, gate1213inter5, gate1213inter6, gate1213inter7, gate1213inter8, gate1213inter9, gate1213inter10, gate1213inter11, gate1213inter12, gate2157inter0, gate2157inter1, gate2157inter2, gate2157inter3, gate2157inter4, gate2157inter5, gate2157inter6, gate2157inter7, gate2157inter8, gate2157inter9, gate2157inter10, gate2157inter11, gate2157inter12, gate1056inter0, gate1056inter1, gate1056inter2, gate1056inter3, gate1056inter4, gate1056inter5, gate1056inter6, gate1056inter7, gate1056inter8, gate1056inter9, gate1056inter10, gate1056inter11, gate1056inter12, gate1319inter0, gate1319inter1, gate1319inter2, gate1319inter3, gate1319inter4, gate1319inter5, gate1319inter6, gate1319inter7, gate1319inter8, gate1319inter9, gate1319inter10, gate1319inter11, gate1319inter12, gate571inter0, gate571inter1, gate571inter2, gate571inter3, gate571inter4, gate571inter5, gate571inter6, gate571inter7, gate571inter8, gate571inter9, gate571inter10, gate571inter11, gate571inter12, gate1788inter0, gate1788inter1, gate1788inter2, gate1788inter3, gate1788inter4, gate1788inter5, gate1788inter6, gate1788inter7, gate1788inter8, gate1788inter9, gate1788inter10, gate1788inter11, gate1788inter12, gate2176inter0, gate2176inter1, gate2176inter2, gate2176inter3, gate2176inter4, gate2176inter5, gate2176inter6, gate2176inter7, gate2176inter8, gate2176inter9, gate2176inter10, gate2176inter11, gate2176inter12, gate1970inter0, gate1970inter1, gate1970inter2, gate1970inter3, gate1970inter4, gate1970inter5, gate1970inter6, gate1970inter7, gate1970inter8, gate1970inter9, gate1970inter10, gate1970inter11, gate1970inter12, gate1232inter0, gate1232inter1, gate1232inter2, gate1232inter3, gate1232inter4, gate1232inter5, gate1232inter6, gate1232inter7, gate1232inter8, gate1232inter9, gate1232inter10, gate1232inter11, gate1232inter12, gate866inter0, gate866inter1, gate866inter2, gate866inter3, gate866inter4, gate866inter5, gate866inter6, gate866inter7, gate866inter8, gate866inter9, gate866inter10, gate866inter11, gate866inter12, gate1635inter0, gate1635inter1, gate1635inter2, gate1635inter3, gate1635inter4, gate1635inter5, gate1635inter6, gate1635inter7, gate1635inter8, gate1635inter9, gate1635inter10, gate1635inter11, gate1635inter12, gate2215inter0, gate2215inter1, gate2215inter2, gate2215inter3, gate2215inter4, gate2215inter5, gate2215inter6, gate2215inter7, gate2215inter8, gate2215inter9, gate2215inter10, gate2215inter11, gate2215inter12, gate2161inter0, gate2161inter1, gate2161inter2, gate2161inter3, gate2161inter4, gate2161inter5, gate2161inter6, gate2161inter7, gate2161inter8, gate2161inter9, gate2161inter10, gate2161inter11, gate2161inter12, gate1252inter0, gate1252inter1, gate1252inter2, gate1252inter3, gate1252inter4, gate1252inter5, gate1252inter6, gate1252inter7, gate1252inter8, gate1252inter9, gate1252inter10, gate1252inter11, gate1252inter12, gate1078inter0, gate1078inter1, gate1078inter2, gate1078inter3, gate1078inter4, gate1078inter5, gate1078inter6, gate1078inter7, gate1078inter8, gate1078inter9, gate1078inter10, gate1078inter11, gate1078inter12, gate2253inter0, gate2253inter1, gate2253inter2, gate2253inter3, gate2253inter4, gate2253inter5, gate2253inter6, gate2253inter7, gate2253inter8, gate2253inter9, gate2253inter10, gate2253inter11, gate2253inter12, gate2251inter0, gate2251inter1, gate2251inter2, gate2251inter3, gate2251inter4, gate2251inter5, gate2251inter6, gate2251inter7, gate2251inter8, gate2251inter9, gate2251inter10, gate2251inter11, gate2251inter12, gate1810inter0, gate1810inter1, gate1810inter2, gate1810inter3, gate1810inter4, gate1810inter5, gate1810inter6, gate1810inter7, gate1810inter8, gate1810inter9, gate1810inter10, gate1810inter11, gate1810inter12, gate2209inter0, gate2209inter1, gate2209inter2, gate2209inter3, gate2209inter4, gate2209inter5, gate2209inter6, gate2209inter7, gate2209inter8, gate2209inter9, gate2209inter10, gate2209inter11, gate2209inter12, gate2031inter0, gate2031inter1, gate2031inter2, gate2031inter3, gate2031inter4, gate2031inter5, gate2031inter6, gate2031inter7, gate2031inter8, gate2031inter9, gate2031inter10, gate2031inter11, gate2031inter12, gate2123inter0, gate2123inter1, gate2123inter2, gate2123inter3, gate2123inter4, gate2123inter5, gate2123inter6, gate2123inter7, gate2123inter8, gate2123inter9, gate2123inter10, gate2123inter11, gate2123inter12, gate1228inter0, gate1228inter1, gate1228inter2, gate1228inter3, gate1228inter4, gate1228inter5, gate1228inter6, gate1228inter7, gate1228inter8, gate1228inter9, gate1228inter10, gate1228inter11, gate1228inter12, gate1774inter0, gate1774inter1, gate1774inter2, gate1774inter3, gate1774inter4, gate1774inter5, gate1774inter6, gate1774inter7, gate1774inter8, gate1774inter9, gate1774inter10, gate1774inter11, gate1774inter12, gate1058inter0, gate1058inter1, gate1058inter2, gate1058inter3, gate1058inter4, gate1058inter5, gate1058inter6, gate1058inter7, gate1058inter8, gate1058inter9, gate1058inter10, gate1058inter11, gate1058inter12, gate1849inter0, gate1849inter1, gate1849inter2, gate1849inter3, gate1849inter4, gate1849inter5, gate1849inter6, gate1849inter7, gate1849inter8, gate1849inter9, gate1849inter10, gate1849inter11, gate1849inter12, gate1866inter0, gate1866inter1, gate1866inter2, gate1866inter3, gate1866inter4, gate1866inter5, gate1866inter6, gate1866inter7, gate1866inter8, gate1866inter9, gate1866inter10, gate1866inter11, gate1866inter12, gate1292inter0, gate1292inter1, gate1292inter2, gate1292inter3, gate1292inter4, gate1292inter5, gate1292inter6, gate1292inter7, gate1292inter8, gate1292inter9, gate1292inter10, gate1292inter11, gate1292inter12, gate1674inter0, gate1674inter1, gate1674inter2, gate1674inter3, gate1674inter4, gate1674inter5, gate1674inter6, gate1674inter7, gate1674inter8, gate1674inter9, gate1674inter10, gate1674inter11, gate1674inter12, gate2143inter0, gate2143inter1, gate2143inter2, gate2143inter3, gate2143inter4, gate2143inter5, gate2143inter6, gate2143inter7, gate2143inter8, gate2143inter9, gate2143inter10, gate2143inter11, gate2143inter12, gate1197inter0, gate1197inter1, gate1197inter2, gate1197inter3, gate1197inter4, gate1197inter5, gate1197inter6, gate1197inter7, gate1197inter8, gate1197inter9, gate1197inter10, gate1197inter11, gate1197inter12, gate2079inter0, gate2079inter1, gate2079inter2, gate2079inter3, gate2079inter4, gate2079inter5, gate2079inter6, gate2079inter7, gate2079inter8, gate2079inter9, gate2079inter10, gate2079inter11, gate2079inter12, gate2189inter0, gate2189inter1, gate2189inter2, gate2189inter3, gate2189inter4, gate2189inter5, gate2189inter6, gate2189inter7, gate2189inter8, gate2189inter9, gate2189inter10, gate2189inter11, gate2189inter12, gate1244inter0, gate1244inter1, gate1244inter2, gate1244inter3, gate1244inter4, gate1244inter5, gate1244inter6, gate1244inter7, gate1244inter8, gate1244inter9, gate1244inter10, gate1244inter11, gate1244inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12, gate2167inter0, gate2167inter1, gate2167inter2, gate2167inter3, gate2167inter4, gate2167inter5, gate2167inter6, gate2167inter7, gate2167inter8, gate2167inter9, gate2167inter10, gate2167inter11, gate2167inter12, gate2138inter0, gate2138inter1, gate2138inter2, gate2138inter3, gate2138inter4, gate2138inter5, gate2138inter6, gate2138inter7, gate2138inter8, gate2138inter9, gate2138inter10, gate2138inter11, gate2138inter12, gate2172inter0, gate2172inter1, gate2172inter2, gate2172inter3, gate2172inter4, gate2172inter5, gate2172inter6, gate2172inter7, gate2172inter8, gate2172inter9, gate2172inter10, gate2172inter11, gate2172inter12, gate2170inter0, gate2170inter1, gate2170inter2, gate2170inter3, gate2170inter4, gate2170inter5, gate2170inter6, gate2170inter7, gate2170inter8, gate2170inter9, gate2170inter10, gate2170inter11, gate2170inter12, gate739inter0, gate739inter1, gate739inter2, gate739inter3, gate739inter4, gate739inter5, gate739inter6, gate739inter7, gate739inter8, gate739inter9, gate739inter10, gate739inter11, gate739inter12, gate1255inter0, gate1255inter1, gate1255inter2, gate1255inter3, gate1255inter4, gate1255inter5, gate1255inter6, gate1255inter7, gate1255inter8, gate1255inter9, gate1255inter10, gate1255inter11, gate1255inter12, gate1096inter0, gate1096inter1, gate1096inter2, gate1096inter3, gate1096inter4, gate1096inter5, gate1096inter6, gate1096inter7, gate1096inter8, gate1096inter9, gate1096inter10, gate1096inter11, gate1096inter12, gate569inter0, gate569inter1, gate569inter2, gate569inter3, gate569inter4, gate569inter5, gate569inter6, gate569inter7, gate569inter8, gate569inter9, gate569inter10, gate569inter11, gate569inter12, gate1971inter0, gate1971inter1, gate1971inter2, gate1971inter3, gate1971inter4, gate1971inter5, gate1971inter6, gate1971inter7, gate1971inter8, gate1971inter9, gate1971inter10, gate1971inter11, gate1971inter12, gate744inter0, gate744inter1, gate744inter2, gate744inter3, gate744inter4, gate744inter5, gate744inter6, gate744inter7, gate744inter8, gate744inter9, gate744inter10, gate744inter11, gate744inter12, gate1889inter0, gate1889inter1, gate1889inter2, gate1889inter3, gate1889inter4, gate1889inter5, gate1889inter6, gate1889inter7, gate1889inter8, gate1889inter9, gate1889inter10, gate1889inter11, gate1889inter12, gate2186inter0, gate2186inter1, gate2186inter2, gate2186inter3, gate2186inter4, gate2186inter5, gate2186inter6, gate2186inter7, gate2186inter8, gate2186inter9, gate2186inter10, gate2186inter11, gate2186inter12, gate1294inter0, gate1294inter1, gate1294inter2, gate1294inter3, gate1294inter4, gate1294inter5, gate1294inter6, gate1294inter7, gate1294inter8, gate1294inter9, gate1294inter10, gate1294inter11, gate1294inter12, gate1856inter0, gate1856inter1, gate1856inter2, gate1856inter3, gate1856inter4, gate1856inter5, gate1856inter6, gate1856inter7, gate1856inter8, gate1856inter9, gate1856inter10, gate1856inter11, gate1856inter12, gate1772inter0, gate1772inter1, gate1772inter2, gate1772inter3, gate1772inter4, gate1772inter5, gate1772inter6, gate1772inter7, gate1772inter8, gate1772inter9, gate1772inter10, gate1772inter11, gate1772inter12, gate1062inter0, gate1062inter1, gate1062inter2, gate1062inter3, gate1062inter4, gate1062inter5, gate1062inter6, gate1062inter7, gate1062inter8, gate1062inter9, gate1062inter10, gate1062inter11, gate1062inter12, gate1904inter0, gate1904inter1, gate1904inter2, gate1904inter3, gate1904inter4, gate1904inter5, gate1904inter6, gate1904inter7, gate1904inter8, gate1904inter9, gate1904inter10, gate1904inter11, gate1904inter12, gate2223inter0, gate2223inter1, gate2223inter2, gate2223inter3, gate2223inter4, gate2223inter5, gate2223inter6, gate2223inter7, gate2223inter8, gate2223inter9, gate2223inter10, gate2223inter11, gate2223inter12, gate2187inter0, gate2187inter1, gate2187inter2, gate2187inter3, gate2187inter4, gate2187inter5, gate2187inter6, gate2187inter7, gate2187inter8, gate2187inter9, gate2187inter10, gate2187inter11, gate2187inter12, gate2270inter0, gate2270inter1, gate2270inter2, gate2270inter3, gate2270inter4, gate2270inter5, gate2270inter6, gate2270inter7, gate2270inter8, gate2270inter9, gate2270inter10, gate2270inter11, gate2270inter12, gate1775inter0, gate1775inter1, gate1775inter2, gate1775inter3, gate1775inter4, gate1775inter5, gate1775inter6, gate1775inter7, gate1775inter8, gate1775inter9, gate1775inter10, gate1775inter11, gate1775inter12, gate2013inter0, gate2013inter1, gate2013inter2, gate2013inter3, gate2013inter4, gate2013inter5, gate2013inter6, gate2013inter7, gate2013inter8, gate2013inter9, gate2013inter10, gate2013inter11, gate2013inter12, gate2016inter0, gate2016inter1, gate2016inter2, gate2016inter3, gate2016inter4, gate2016inter5, gate2016inter6, gate2016inter7, gate2016inter8, gate2016inter9, gate2016inter10, gate2016inter11, gate2016inter12, gate2155inter0, gate2155inter1, gate2155inter2, gate2155inter3, gate2155inter4, gate2155inter5, gate2155inter6, gate2155inter7, gate2155inter8, gate2155inter9, gate2155inter10, gate2155inter11, gate2155inter12, gate2179inter0, gate2179inter1, gate2179inter2, gate2179inter3, gate2179inter4, gate2179inter5, gate2179inter6, gate2179inter7, gate2179inter8, gate2179inter9, gate2179inter10, gate2179inter11, gate2179inter12, gate1189inter0, gate1189inter1, gate1189inter2, gate1189inter3, gate1189inter4, gate1189inter5, gate1189inter6, gate1189inter7, gate1189inter8, gate1189inter9, gate1189inter10, gate1189inter11, gate1189inter12, gate2106inter0, gate2106inter1, gate2106inter2, gate2106inter3, gate2106inter4, gate2106inter5, gate2106inter6, gate2106inter7, gate2106inter8, gate2106inter9, gate2106inter10, gate2106inter11, gate2106inter12, gate1119inter0, gate1119inter1, gate1119inter2, gate1119inter3, gate1119inter4, gate1119inter5, gate1119inter6, gate1119inter7, gate1119inter8, gate1119inter9, gate1119inter10, gate1119inter11, gate1119inter12, gate2192inter0, gate2192inter1, gate2192inter2, gate2192inter3, gate2192inter4, gate2192inter5, gate2192inter6, gate2192inter7, gate2192inter8, gate2192inter9, gate2192inter10, gate2192inter11, gate2192inter12, gate2159inter0, gate2159inter1, gate2159inter2, gate2159inter3, gate2159inter4, gate2159inter5, gate2159inter6, gate2159inter7, gate2159inter8, gate2159inter9, gate2159inter10, gate2159inter11, gate2159inter12, gate1108inter0, gate1108inter1, gate1108inter2, gate1108inter3, gate1108inter4, gate1108inter5, gate1108inter6, gate1108inter7, gate1108inter8, gate1108inter9, gate1108inter10, gate1108inter11, gate1108inter12, gate1038inter0, gate1038inter1, gate1038inter2, gate1038inter3, gate1038inter4, gate1038inter5, gate1038inter6, gate1038inter7, gate1038inter8, gate1038inter9, gate1038inter10, gate1038inter11, gate1038inter12, gate1671inter0, gate1671inter1, gate1671inter2, gate1671inter3, gate1671inter4, gate1671inter5, gate1671inter6, gate1671inter7, gate1671inter8, gate1671inter9, gate1671inter10, gate1671inter11, gate1671inter12, gate2191inter0, gate2191inter1, gate2191inter2, gate2191inter3, gate2191inter4, gate2191inter5, gate2191inter6, gate2191inter7, gate2191inter8, gate2191inter9, gate2191inter10, gate2191inter11, gate2191inter12, gate1741inter0, gate1741inter1, gate1741inter2, gate1741inter3, gate1741inter4, gate1741inter5, gate1741inter6, gate1741inter7, gate1741inter8, gate1741inter9, gate1741inter10, gate1741inter11, gate1741inter12, gate1269inter0, gate1269inter1, gate1269inter2, gate1269inter3, gate1269inter4, gate1269inter5, gate1269inter6, gate1269inter7, gate1269inter8, gate1269inter9, gate1269inter10, gate1269inter11, gate1269inter12, gate1089inter0, gate1089inter1, gate1089inter2, gate1089inter3, gate1089inter4, gate1089inter5, gate1089inter6, gate1089inter7, gate1089inter8, gate1089inter9, gate1089inter10, gate1089inter11, gate1089inter12, gate2244inter0, gate2244inter1, gate2244inter2, gate2244inter3, gate2244inter4, gate2244inter5, gate2244inter6, gate2244inter7, gate2244inter8, gate2244inter9, gate2244inter10, gate2244inter11, gate2244inter12, gate1091inter0, gate1091inter1, gate1091inter2, gate1091inter3, gate1091inter4, gate1091inter5, gate1091inter6, gate1091inter7, gate1091inter8, gate1091inter9, gate1091inter10, gate1091inter11, gate1091inter12, gate2124inter0, gate2124inter1, gate2124inter2, gate2124inter3, gate2124inter4, gate2124inter5, gate2124inter6, gate2124inter7, gate2124inter8, gate2124inter9, gate2124inter10, gate2124inter11, gate2124inter12, gate1732inter0, gate1732inter1, gate1732inter2, gate1732inter3, gate1732inter4, gate1732inter5, gate1732inter6, gate1732inter7, gate1732inter8, gate1732inter9, gate1732inter10, gate1732inter11, gate1732inter12, gate2193inter0, gate2193inter1, gate2193inter2, gate2193inter3, gate2193inter4, gate2193inter5, gate2193inter6, gate2193inter7, gate2193inter8, gate2193inter9, gate2193inter10, gate2193inter11, gate2193inter12, gate2012inter0, gate2012inter1, gate2012inter2, gate2012inter3, gate2012inter4, gate2012inter5, gate2012inter6, gate2012inter7, gate2012inter8, gate2012inter9, gate2012inter10, gate2012inter11, gate2012inter12, gate2014inter0, gate2014inter1, gate2014inter2, gate2014inter3, gate2014inter4, gate2014inter5, gate2014inter6, gate2014inter7, gate2014inter8, gate2014inter9, gate2014inter10, gate2014inter11, gate2014inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate1558inter0, gate1558inter1, gate1558inter2, gate1558inter3, gate1558inter4, gate1558inter5, gate1558inter6, gate1558inter7, gate1558inter8, gate1558inter9, gate1558inter10, gate1558inter11, gate1558inter12, gate1050inter0, gate1050inter1, gate1050inter2, gate1050inter3, gate1050inter4, gate1050inter5, gate1050inter6, gate1050inter7, gate1050inter8, gate1050inter9, gate1050inter10, gate1050inter11, gate1050inter12, gate975inter0, gate975inter1, gate975inter2, gate975inter3, gate975inter4, gate975inter5, gate975inter6, gate975inter7, gate975inter8, gate975inter9, gate975inter10, gate975inter11, gate975inter12, gate1784inter0, gate1784inter1, gate1784inter2, gate1784inter3, gate1784inter4, gate1784inter5, gate1784inter6, gate1784inter7, gate1784inter8, gate1784inter9, gate1784inter10, gate1784inter11, gate1784inter12, gate2203inter0, gate2203inter1, gate2203inter2, gate2203inter3, gate2203inter4, gate2203inter5, gate2203inter6, gate2203inter7, gate2203inter8, gate2203inter9, gate2203inter10, gate2203inter11, gate2203inter12, gate1068inter0, gate1068inter1, gate1068inter2, gate1068inter3, gate1068inter4, gate1068inter5, gate1068inter6, gate1068inter7, gate1068inter8, gate1068inter9, gate1068inter10, gate1068inter11, gate1068inter12, gate2134inter0, gate2134inter1, gate2134inter2, gate2134inter3, gate2134inter4, gate2134inter5, gate2134inter6, gate2134inter7, gate2134inter8, gate2134inter9, gate2134inter10, gate2134inter11, gate2134inter12, gate2006inter0, gate2006inter1, gate2006inter2, gate2006inter3, gate2006inter4, gate2006inter5, gate2006inter6, gate2006inter7, gate2006inter8, gate2006inter9, gate2006inter10, gate2006inter11, gate2006inter12, gate1865inter0, gate1865inter1, gate1865inter2, gate1865inter3, gate1865inter4, gate1865inter5, gate1865inter6, gate1865inter7, gate1865inter8, gate1865inter9, gate1865inter10, gate1865inter11, gate1865inter12, gate2007inter0, gate2007inter1, gate2007inter2, gate2007inter3, gate2007inter4, gate2007inter5, gate2007inter6, gate2007inter7, gate2007inter8, gate2007inter9, gate2007inter10, gate2007inter11, gate2007inter12, gate1173inter0, gate1173inter1, gate1173inter2, gate1173inter3, gate1173inter4, gate1173inter5, gate1173inter6, gate1173inter7, gate1173inter8, gate1173inter9, gate1173inter10, gate1173inter11, gate1173inter12, gate2108inter0, gate2108inter1, gate2108inter2, gate2108inter3, gate2108inter4, gate2108inter5, gate2108inter6, gate2108inter7, gate2108inter8, gate2108inter9, gate2108inter10, gate2108inter11, gate2108inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate1854inter0, gate1854inter1, gate1854inter2, gate1854inter3, gate1854inter4, gate1854inter5, gate1854inter6, gate1854inter7, gate1854inter8, gate1854inter9, gate1854inter10, gate1854inter11, gate1854inter12, gate1226inter0, gate1226inter1, gate1226inter2, gate1226inter3, gate1226inter4, gate1226inter5, gate1226inter6, gate1226inter7, gate1226inter8, gate1226inter9, gate1226inter10, gate1226inter11, gate1226inter12, gate1293inter0, gate1293inter1, gate1293inter2, gate1293inter3, gate1293inter4, gate1293inter5, gate1293inter6, gate1293inter7, gate1293inter8, gate1293inter9, gate1293inter10, gate1293inter11, gate1293inter12, gate1280inter0, gate1280inter1, gate1280inter2, gate1280inter3, gate1280inter4, gate1280inter5, gate1280inter6, gate1280inter7, gate1280inter8, gate1280inter9, gate1280inter10, gate1280inter11, gate1280inter12, gate1186inter0, gate1186inter1, gate1186inter2, gate1186inter3, gate1186inter4, gate1186inter5, gate1186inter6, gate1186inter7, gate1186inter8, gate1186inter9, gate1186inter10, gate1186inter11, gate1186inter12, gate1182inter0, gate1182inter1, gate1182inter2, gate1182inter3, gate1182inter4, gate1182inter5, gate1182inter6, gate1182inter7, gate1182inter8, gate1182inter9, gate1182inter10, gate1182inter11, gate1182inter12, gate2107inter0, gate2107inter1, gate2107inter2, gate2107inter3, gate2107inter4, gate2107inter5, gate2107inter6, gate2107inter7, gate2107inter8, gate2107inter9, gate2107inter10, gate2107inter11, gate2107inter12;



buf1 gate1( .a(N141), .O(N709) );
buf1 gate2( .a(N293), .O(N816) );
and2 gate3( .a(N135), .b(N631), .O(N1042) );
inv1 gate4( .a(N591), .O(N1043) );
buf1 gate5( .a(N592), .O(N1066) );
inv1 gate6( .a(N595), .O(N1067) );
inv1 gate7( .a(N596), .O(N1080) );
inv1 gate8( .a(N597), .O(N1092) );
inv1 gate9( .a(N598), .O(N1104) );
inv1 gate10( .a(N545), .O(N1137) );
inv1 gate11( .a(N348), .O(N1138) );
inv1 gate12( .a(N366), .O(N1139) );
and2 gate13( .a(N552), .b(N562), .O(N1140) );
inv1 gate14( .a(N549), .O(N1141) );
inv1 gate15( .a(N545), .O(N1142) );
inv1 gate16( .a(N545), .O(N1143) );
inv1 gate17( .a(N338), .O(N1144) );
inv1 gate18( .a(N358), .O(N1145) );
nand2 gate19( .a(N373), .b(N1), .O(N1146) );
and2 gate20( .a(N141), .b(N145), .O(N1147) );
inv1 gate21( .a(N592), .O(N1148) );
inv1 gate22( .a(N1042), .O(N1149) );
and2 gate23( .a(N1043), .b(N27), .O(N1150) );
and2 gate24( .a(N386), .b(N556), .O(N1151) );
inv1 gate25( .a(N245), .O(N1152) );
inv1 gate26( .a(N552), .O(N1153) );
inv1 gate27( .a(N562), .O(N1154) );
inv1 gate28( .a(N559), .O(N1155) );
and4 gate29( .a(N386), .b(N559), .c(N556), .d(N552), .O(N1156) );
inv1 gate30( .a(N566), .O(N1157) );
buf1 gate31( .a(N571), .O(N1161) );
buf1 gate32( .a(N574), .O(N1173) );
buf1 gate33( .a(N571), .O(N1185) );
buf1 gate34( .a(N574), .O(N1197) );
buf1 gate35( .a(N137), .O(N1209) );
buf1 gate36( .a(N137), .O(N1213) );
buf1 gate37( .a(N141), .O(N1216) );
inv1 gate38( .a(N583), .O(N1219) );
buf1 gate39( .a(N577), .O(N1223) );
buf1 gate40( .a(N580), .O(N1235) );
buf1 gate41( .a(N577), .O(N1247) );
buf1 gate42( .a(N580), .O(N1259) );
buf1 gate43( .a(N254), .O(N1271) );
buf1 gate44( .a(N251), .O(N1280) );
buf1 gate45( .a(N251), .O(N1292) );
buf1 gate46( .a(N248), .O(N1303) );
buf1 gate47( .a(N248), .O(N1315) );
buf1 gate48( .a(N610), .O(N1327) );
buf1 gate49( .a(N607), .O(N1339) );
buf1 gate50( .a(N613), .O(N1351) );
buf1 gate51( .a(N616), .O(N1363) );
buf1 gate52( .a(N210), .O(N1375) );
buf1 gate53( .a(N210), .O(N1378) );
buf1 gate54( .a(N218), .O(N1381) );
buf1 gate55( .a(N218), .O(N1384) );
buf1 gate56( .a(N226), .O(N1387) );
buf1 gate57( .a(N226), .O(N1390) );
buf1 gate58( .a(N234), .O(N1393) );
buf1 gate59( .a(N234), .O(N1396) );
buf1 gate60( .a(N257), .O(N1415) );
buf1 gate61( .a(N257), .O(N1418) );
buf1 gate62( .a(N265), .O(N1421) );
buf1 gate63( .a(N265), .O(N1424) );
buf1 gate64( .a(N273), .O(N1427) );
buf1 gate65( .a(N273), .O(N1430) );
buf1 gate66( .a(N281), .O(N1433) );
buf1 gate67( .a(N281), .O(N1436) );
buf1 gate68( .a(N335), .O(N1455) );
buf1 gate69( .a(N335), .O(N1462) );
buf1 gate70( .a(N206), .O(N1469) );
and2 gate71( .a(N27), .b(N31), .O(N1475) );
buf1 gate72( .a(N1), .O(N1479) );
buf1 gate73( .a(N588), .O(N1482) );
buf1 gate74( .a(N293), .O(N1492) );
buf1 gate75( .a(N302), .O(N1495) );
buf1 gate76( .a(N308), .O(N1498) );
buf1 gate77( .a(N308), .O(N1501) );
buf1 gate78( .a(N316), .O(N1504) );
buf1 gate79( .a(N316), .O(N1507) );
buf1 gate80( .a(N324), .O(N1510) );
buf1 gate81( .a(N324), .O(N1513) );
buf1 gate82( .a(N341), .O(N1516) );
buf1 gate83( .a(N341), .O(N1519) );
buf1 gate84( .a(N351), .O(N1522) );
buf1 gate85( .a(N351), .O(N1525) );
buf1 gate86( .a(N257), .O(N1542) );
buf1 gate87( .a(N257), .O(N1545) );
buf1 gate88( .a(N265), .O(N1548) );
buf1 gate89( .a(N265), .O(N1551) );
buf1 gate90( .a(N273), .O(N1554) );
buf1 gate91( .a(N273), .O(N1557) );
buf1 gate92( .a(N281), .O(N1560) );
buf1 gate93( .a(N281), .O(N1563) );
buf1 gate94( .a(N332), .O(N1566) );
buf1 gate95( .a(N332), .O(N1573) );
buf1 gate96( .a(N549), .O(N1580) );
and2 gate97( .a(N31), .b(N27), .O(N1583) );
inv1 gate98( .a(N588), .O(N1588) );
buf1 gate99( .a(N324), .O(N1594) );
buf1 gate100( .a(N324), .O(N1597) );
buf1 gate101( .a(N341), .O(N1600) );
buf1 gate102( .a(N341), .O(N1603) );
buf1 gate103( .a(N351), .O(N1606) );
buf1 gate104( .a(N351), .O(N1609) );
buf1 gate105( .a(N293), .O(N1612) );
buf1 gate106( .a(N302), .O(N1615) );
buf1 gate107( .a(N308), .O(N1618) );
buf1 gate108( .a(N308), .O(N1621) );
buf1 gate109( .a(N316), .O(N1624) );
buf1 gate110( .a(N316), .O(N1627) );
buf1 gate111( .a(N361), .O(N1630) );
buf1 gate112( .a(N361), .O(N1633) );
buf1 gate113( .a(N210), .O(N1636) );
buf1 gate114( .a(N210), .O(N1639) );
buf1 gate115( .a(N218), .O(N1642) );
buf1 gate116( .a(N218), .O(N1645) );
buf1 gate117( .a(N226), .O(N1648) );
buf1 gate118( .a(N226), .O(N1651) );
buf1 gate119( .a(N234), .O(N1654) );
buf1 gate120( .a(N234), .O(N1657) );
inv1 gate121( .a(N324), .O(N1660) );
buf1 gate122( .a(N242), .O(N1663) );
buf1 gate123( .a(N242), .O(N1675) );
buf1 gate124( .a(N254), .O(N1685) );
buf1 gate125( .a(N610), .O(N1697) );
buf1 gate126( .a(N607), .O(N1709) );
buf1 gate127( .a(N625), .O(N1721) );
buf1 gate128( .a(N619), .O(N1727) );
buf1 gate129( .a(N613), .O(N1731) );
buf1 gate130( .a(N616), .O(N1743) );
inv1 gate131( .a(N599), .O(N1755) );
inv1 gate132( .a(N603), .O(N1758) );
buf1 gate133( .a(N619), .O(N1761) );
buf1 gate134( .a(N625), .O(N1769) );
buf1 gate135( .a(N619), .O(N1777) );
buf1 gate136( .a(N625), .O(N1785) );
buf1 gate137( .a(N619), .O(N1793) );
buf1 gate138( .a(N625), .O(N1800) );
buf1 gate139( .a(N619), .O(N1807) );
buf1 gate140( .a(N625), .O(N1814) );
buf1 gate141( .a(N299), .O(N1821) );
buf1 gate142( .a(N446), .O(N1824) );
buf1 gate143( .a(N457), .O(N1827) );
buf1 gate144( .a(N468), .O(N1830) );
buf1 gate145( .a(N422), .O(N1833) );
buf1 gate146( .a(N435), .O(N1836) );
buf1 gate147( .a(N389), .O(N1839) );
buf1 gate148( .a(N400), .O(N1842) );
buf1 gate149( .a(N411), .O(N1845) );
buf1 gate150( .a(N374), .O(N1848) );
buf1 gate151( .a(N4), .O(N1851) );
buf1 gate152( .a(N446), .O(N1854) );
buf1 gate153( .a(N457), .O(N1857) );
buf1 gate154( .a(N468), .O(N1860) );
buf1 gate155( .a(N435), .O(N1863) );
buf1 gate156( .a(N389), .O(N1866) );
buf1 gate157( .a(N400), .O(N1869) );
buf1 gate158( .a(N411), .O(N1872) );
buf1 gate159( .a(N422), .O(N1875) );
buf1 gate160( .a(N374), .O(N1878) );
buf1 gate161( .a(N479), .O(N1881) );
buf1 gate162( .a(N490), .O(N1884) );
buf1 gate163( .a(N503), .O(N1887) );
buf1 gate164( .a(N514), .O(N1890) );
buf1 gate165( .a(N523), .O(N1893) );
buf1 gate166( .a(N534), .O(N1896) );
buf1 gate167( .a(N54), .O(N1899) );
buf1 gate168( .a(N479), .O(N1902) );
buf1 gate169( .a(N503), .O(N1905) );
buf1 gate170( .a(N514), .O(N1908) );
buf1 gate171( .a(N523), .O(N1911) );
buf1 gate172( .a(N534), .O(N1914) );
buf1 gate173( .a(N490), .O(N1917) );
buf1 gate174( .a(N361), .O(N1920) );
buf1 gate175( .a(N369), .O(N1923) );
buf1 gate176( .a(N341), .O(N1926) );
buf1 gate177( .a(N351), .O(N1929) );
buf1 gate178( .a(N308), .O(N1932) );
buf1 gate179( .a(N316), .O(N1935) );
buf1 gate180( .a(N293), .O(N1938) );
buf1 gate181( .a(N302), .O(N1941) );
buf1 gate182( .a(N281), .O(N1944) );
buf1 gate183( .a(N289), .O(N1947) );
buf1 gate184( .a(N265), .O(N1950) );
buf1 gate185( .a(N273), .O(N1953) );
buf1 gate186( .a(N234), .O(N1956) );
buf1 gate187( .a(N257), .O(N1959) );
buf1 gate188( .a(N218), .O(N1962) );
buf1 gate189( .a(N226), .O(N1965) );
buf1 gate190( .a(N210), .O(N1968) );
inv1 gate191( .a(N1146), .O(N1972) );
and2 gate192( .a(N136), .b(N1148), .O(N2054) );
inv1 gate193( .a(N1150), .O(N2060) );
inv1 gate194( .a(N1151), .O(N2061) );
buf1 gate195( .a(N1209), .O(N2139) );
buf1 gate196( .a(N1216), .O(N2142) );
buf1 gate197( .a(N1479), .O(N2309) );
and2 gate198( .a(N1104), .b(N514), .O(N2349) );
or2 gate199( .a(N1067), .b(N514), .O(N2350) );
buf1 gate200( .a(N1580), .O(N2387) );
buf1 gate201( .a(N1821), .O(N2527) );
inv1 gate202( .a(N1580), .O(N2584) );
and3 gate203( .a(N170), .b(N1161), .c(N1173), .O(N2585) );
and3 gate204( .a(N173), .b(N1161), .c(N1173), .O(N2586) );
and3 gate205( .a(N167), .b(N1161), .c(N1173), .O(N2587) );
and3 gate206( .a(N164), .b(N1161), .c(N1173), .O(N2588) );
and3 gate207( .a(N161), .b(N1161), .c(N1173), .O(N2589) );
nand2 gate208( .a(N1475), .b(N140), .O(N2590) );
and3 gate209( .a(N185), .b(N1185), .c(N1197), .O(N2591) );
and3 gate210( .a(N158), .b(N1185), .c(N1197), .O(N2592) );
and3 gate211( .a(N152), .b(N1185), .c(N1197), .O(N2593) );
and3 gate212( .a(N146), .b(N1185), .c(N1197), .O(N2594) );
and3 gate213( .a(N170), .b(N1223), .c(N1235), .O(N2595) );
and3 gate214( .a(N173), .b(N1223), .c(N1235), .O(N2596) );
and3 gate215( .a(N167), .b(N1223), .c(N1235), .O(N2597) );
and3 gate216( .a(N164), .b(N1223), .c(N1235), .O(N2598) );
and3 gate217( .a(N161), .b(N1223), .c(N1235), .O(N2599) );
and3 gate218( .a(N185), .b(N1247), .c(N1259), .O(N2600) );
and3 gate219( .a(N158), .b(N1247), .c(N1259), .O(N2601) );
and3 gate220( .a(N152), .b(N1247), .c(N1259), .O(N2602) );
and3 gate221( .a(N146), .b(N1247), .c(N1259), .O(N2603) );
and3 gate222( .a(N106), .b(N1731), .c(N1743), .O(N2604) );
and3 gate223( .a(N61), .b(N1327), .c(N1339), .O(N2605) );
and3 gate224( .a(N106), .b(N1697), .c(N1709), .O(N2606) );
and3 gate225( .a(N49), .b(N1697), .c(N1709), .O(N2607) );
and3 gate226( .a(N103), .b(N1697), .c(N1709), .O(N2608) );
and3 gate227( .a(N40), .b(N1697), .c(N1709), .O(N2609) );
and3 gate228( .a(N37), .b(N1697), .c(N1709), .O(N2610) );
and3 gate229( .a(N20), .b(N1327), .c(N1339), .O(N2611) );
and3 gate230( .a(N17), .b(N1327), .c(N1339), .O(N2612) );
and3 gate231( .a(N70), .b(N1327), .c(N1339), .O(N2613) );
and3 gate232( .a(N64), .b(N1327), .c(N1339), .O(N2614) );
and3 gate233( .a(N49), .b(N1731), .c(N1743), .O(N2615) );
and3 gate234( .a(N103), .b(N1731), .c(N1743), .O(N2616) );
and3 gate235( .a(N40), .b(N1731), .c(N1743), .O(N2617) );
and3 gate236( .a(N37), .b(N1731), .c(N1743), .O(N2618) );
and3 gate237( .a(N20), .b(N1351), .c(N1363), .O(N2619) );
and3 gate238( .a(N17), .b(N1351), .c(N1363), .O(N2620) );
and3 gate239( .a(N70), .b(N1351), .c(N1363), .O(N2621) );
and3 gate240( .a(N64), .b(N1351), .c(N1363), .O(N2622) );
inv1 gate241( .a(N1475), .O(N2623) );
and3 gate242( .a(N123), .b(N1758), .c(N599), .O(N2624) );
and2 gate243( .a(N1777), .b(N1785), .O(N2625) );
and3 gate244( .a(N61), .b(N1351), .c(N1363), .O(N2626) );
and2 gate245( .a(N1761), .b(N1769), .O(N2627) );
inv1 gate246( .a(N1824), .O(N2628) );
inv1 gate247( .a(N1827), .O(N2629) );
inv1 gate248( .a(N1830), .O(N2630) );
inv1 gate249( .a(N1833), .O(N2631) );
inv1 gate250( .a(N1836), .O(N2632) );
inv1 gate251( .a(N1839), .O(N2633) );
inv1 gate252( .a(N1842), .O(N2634) );
inv1 gate253( .a(N1845), .O(N2635) );
inv1 gate254( .a(N1848), .O(N2636) );
inv1 gate255( .a(N1851), .O(N2637) );
inv1 gate256( .a(N1854), .O(N2638) );
inv1 gate257( .a(N1857), .O(N2639) );
inv1 gate258( .a(N1860), .O(N2640) );
inv1 gate259( .a(N1863), .O(N2641) );
inv1 gate260( .a(N1866), .O(N2642) );
inv1 gate261( .a(N1869), .O(N2643) );
inv1 gate262( .a(N1872), .O(N2644) );
inv1 gate263( .a(N1875), .O(N2645) );
inv1 gate264( .a(N1878), .O(N2646) );
buf1 gate265( .a(N1209), .O(N2647) );
inv1 gate266( .a(N1161), .O(N2653) );
inv1 gate267( .a(N1173), .O(N2664) );
buf1 gate268( .a(N1209), .O(N2675) );
inv1 gate269( .a(N1185), .O(N2681) );
inv1 gate270( .a(N1197), .O(N2692) );
and3 gate271( .a(N179), .b(N1185), .c(N1197), .O(N2703) );
buf1 gate272( .a(N1479), .O(N2704) );
inv1 gate273( .a(N1881), .O(N2709) );
inv1 gate274( .a(N1884), .O(N2710) );
inv1 gate275( .a(N1887), .O(N2711) );
inv1 gate276( .a(N1890), .O(N2712) );
inv1 gate277( .a(N1893), .O(N2713) );
inv1 gate278( .a(N1896), .O(N2714) );
inv1 gate279( .a(N1899), .O(N2715) );
inv1 gate280( .a(N1902), .O(N2716) );
inv1 gate281( .a(N1905), .O(N2717) );
inv1 gate282( .a(N1908), .O(N2718) );
inv1 gate283( .a(N1911), .O(N2719) );
inv1 gate284( .a(N1914), .O(N2720) );
inv1 gate285( .a(N1917), .O(N2721) );
buf1 gate286( .a(N1213), .O(N2722) );
inv1 gate287( .a(N1223), .O(N2728) );
inv1 gate288( .a(N1235), .O(N2739) );
buf1 gate289( .a(N1213), .O(N2750) );
inv1 gate290( .a(N1247), .O(N2756) );
inv1 gate291( .a(N1259), .O(N2767) );
and3 gate292( .a(N179), .b(N1247), .c(N1259), .O(N2778) );
inv1 gate293( .a(N1327), .O(N2779) );
inv1 gate294( .a(N1339), .O(N2790) );
inv1 gate295( .a(N1351), .O(N2801) );
inv1 gate296( .a(N1363), .O(N2812) );
inv1 gate297( .a(N1375), .O(N2823) );
inv1 gate298( .a(N1378), .O(N2824) );
inv1 gate299( .a(N1381), .O(N2825) );
inv1 gate300( .a(N1384), .O(N2826) );
inv1 gate301( .a(N1387), .O(N2827) );
inv1 gate302( .a(N1390), .O(N2828) );
inv1 gate303( .a(N1393), .O(N2829) );
inv1 gate304( .a(N1396), .O(N2830) );
and3 gate305( .a(N1104), .b(N457), .c(N1378), .O(N2831) );
and3 gate306( .a(N1104), .b(N468), .c(N1384), .O(N2832) );
and3 gate307( .a(N1104), .b(N422), .c(N1390), .O(N2833) );
and3 gate308( .a(N1104), .b(N435), .c(N1396), .O(N2834) );
and2 gate309( .a(N1067), .b(N1375), .O(N2835) );
and2 gate310( .a(N1067), .b(N1381), .O(N2836) );
and2 gate311( .a(N1067), .b(N1387), .O(N2837) );
and2 gate312( .a(N1067), .b(N1393), .O(N2838) );
inv1 gate313( .a(N1415), .O(N2839) );
inv1 gate314( .a(N1418), .O(N2840) );
inv1 gate315( .a(N1421), .O(N2841) );
inv1 gate316( .a(N1424), .O(N2842) );
inv1 gate317( .a(N1427), .O(N2843) );
inv1 gate318( .a(N1430), .O(N2844) );
inv1 gate319( .a(N1433), .O(N2845) );
inv1 gate320( .a(N1436), .O(N2846) );
and3 gate321( .a(N1104), .b(N389), .c(N1418), .O(N2847) );
and3 gate322( .a(N1104), .b(N400), .c(N1424), .O(N2848) );
and3 gate323( .a(N1104), .b(N411), .c(N1430), .O(N2849) );
and3 gate324( .a(N1104), .b(N374), .c(N1436), .O(N2850) );
and2 gate325( .a(N1067), .b(N1415), .O(N2851) );
and2 gate326( .a(N1067), .b(N1421), .O(N2852) );
and2 gate327( .a(N1067), .b(N1427), .O(N2853) );
and2 gate328( .a(N1067), .b(N1433), .O(N2854) );
inv1 gate329( .a(N1455), .O(N2855) );
inv1 gate330( .a(N1462), .O(N2861) );
and2 gate331( .a(N292), .b(N1455), .O(N2867) );
and2 gate332( .a(N288), .b(N1455), .O(N2868) );
and2 gate333( .a(N280), .b(N1455), .O(N2869) );
and2 gate334( .a(N272), .b(N1455), .O(N2870) );
and2 gate335( .a(N264), .b(N1455), .O(N2871) );
and2 gate336( .a(N241), .b(N1462), .O(N2872) );
and2 gate337( .a(N233), .b(N1462), .O(N2873) );
and2 gate338( .a(N225), .b(N1462), .O(N2874) );
and2 gate339( .a(N217), .b(N1462), .O(N2875) );
and2 gate340( .a(N209), .b(N1462), .O(N2876) );
buf1 gate341( .a(N1216), .O(N2877) );
inv1 gate342( .a(N1482), .O(N2882) );
inv1 gate343( .a(N1475), .O(N2891) );
inv1 gate344( .a(N1492), .O(N2901) );
inv1 gate345( .a(N1495), .O(N2902) );
inv1 gate346( .a(N1498), .O(N2903) );
inv1 gate347( .a(N1501), .O(N2904) );
inv1 gate348( .a(N1504), .O(N2905) );
inv1 gate349( .a(N1507), .O(N2906) );
and2 gate350( .a(N1303), .b(N1495), .O(N2907) );
and3 gate351( .a(N1303), .b(N479), .c(N1501), .O(N2908) );
and3 gate352( .a(N1303), .b(N490), .c(N1507), .O(N2909) );
and2 gate353( .a(N1663), .b(N1492), .O(N2910) );
and2 gate354( .a(N1663), .b(N1498), .O(N2911) );
and2 gate355( .a(N1663), .b(N1504), .O(N2912) );
inv1 gate356( .a(N1510), .O(N2913) );
inv1 gate357( .a(N1513), .O(N2914) );
inv1 gate358( .a(N1516), .O(N2915) );
inv1 gate359( .a(N1519), .O(N2916) );
inv1 gate360( .a(N1522), .O(N2917) );
inv1 gate361( .a(N1525), .O(N2918) );
and3 gate362( .a(N1104), .b(N503), .c(N1513), .O(N2919) );
inv1 gate363( .a(N2349), .O(N2920) );
and3 gate364( .a(N1104), .b(N523), .c(N1519), .O(N2921) );
and3 gate365( .a(N1104), .b(N534), .c(N1525), .O(N2922) );
and2 gate366( .a(N1067), .b(N1510), .O(N2923) );
and2 gate367( .a(N1067), .b(N1516), .O(N2924) );
and2 gate368( .a(N1067), .b(N1522), .O(N2925) );
inv1 gate369( .a(N1542), .O(N2926) );
inv1 gate370( .a(N1545), .O(N2927) );
inv1 gate371( .a(N1548), .O(N2928) );
inv1 gate372( .a(N1551), .O(N2929) );
inv1 gate373( .a(N1554), .O(N2930) );
inv1 gate374( .a(N1557), .O(N2931) );
inv1 gate375( .a(N1560), .O(N2932) );
inv1 gate376( .a(N1563), .O(N2933) );
and3 gate377( .a(N1303), .b(N389), .c(N1545), .O(N2934) );
and3 gate378( .a(N1303), .b(N400), .c(N1551), .O(N2935) );
and3 gate379( .a(N1303), .b(N411), .c(N1557), .O(N2936) );
and3 gate380( .a(N1303), .b(N374), .c(N1563), .O(N2937) );
and2 gate381( .a(N1663), .b(N1542), .O(N2938) );
and2 gate382( .a(N1663), .b(N1548), .O(N2939) );
and2 gate383( .a(N1663), .b(N1554), .O(N2940) );
and2 gate384( .a(N1663), .b(N1560), .O(N2941) );
inv1 gate385( .a(N1566), .O(N2942) );
inv1 gate386( .a(N1573), .O(N2948) );
and2 gate387( .a(N372), .b(N1566), .O(N2954) );
and2 gate388( .a(N366), .b(N1566), .O(N2955) );
and2 gate389( .a(N358), .b(N1566), .O(N2956) );
and2 gate390( .a(N348), .b(N1566), .O(N2957) );
and2 gate391( .a(N338), .b(N1566), .O(N2958) );
and2 gate392( .a(N331), .b(N1573), .O(N2959) );
and2 gate393( .a(N323), .b(N1573), .O(N2960) );
and2 gate394( .a(N315), .b(N1573), .O(N2961) );
and2 gate395( .a(N307), .b(N1573), .O(N2962) );
and2 gate396( .a(N299), .b(N1573), .O(N2963) );
inv1 gate397( .a(N1588), .O(N2964) );
and2 gate398( .a(N83), .b(N1588), .O(N2969) );
and2 gate399( .a(N86), .b(N1588), .O(N2970) );
and2 gate400( .a(N88), .b(N1588), .O(N2971) );
and2 gate401( .a(N88), .b(N1588), .O(N2972) );
inv1 gate402( .a(N1594), .O(N2973) );
inv1 gate403( .a(N1597), .O(N2974) );
inv1 gate404( .a(N1600), .O(N2975) );
inv1 gate405( .a(N1603), .O(N2976) );
inv1 gate406( .a(N1606), .O(N2977) );
inv1 gate407( .a(N1609), .O(N2978) );
and3 gate408( .a(N1315), .b(N503), .c(N1597), .O(N2979) );
and2 gate409( .a(N1315), .b(N514), .O(N2980) );
and3 gate410( .a(N1315), .b(N523), .c(N1603), .O(N2981) );
and3 gate411( .a(N1315), .b(N534), .c(N1609), .O(N2982) );
and2 gate412( .a(N1675), .b(N1594), .O(N2983) );
or2 gate413( .a(N1675), .b(N514), .O(N2984) );
and2 gate414( .a(N1675), .b(N1600), .O(N2985) );
and2 gate415( .a(N1675), .b(N1606), .O(N2986) );
inv1 gate416( .a(N1612), .O(N2987) );
inv1 gate417( .a(N1615), .O(N2988) );
inv1 gate418( .a(N1618), .O(N2989) );
inv1 gate419( .a(N1621), .O(N2990) );
inv1 gate420( .a(N1624), .O(N2991) );
inv1 gate421( .a(N1627), .O(N2992) );
and2 gate422( .a(N1315), .b(N1615), .O(N2993) );
and3 gate423( .a(N1315), .b(N479), .c(N1621), .O(N2994) );
and3 gate424( .a(N1315), .b(N490), .c(N1627), .O(N2995) );
and2 gate425( .a(N1675), .b(N1612), .O(N2996) );
and2 gate426( .a(N1675), .b(N1618), .O(N2997) );
and2 gate427( .a(N1675), .b(N1624), .O(N2998) );
inv1 gate428( .a(N1630), .O(N2999) );
buf1 gate429( .a(N1469), .O(N3000) );
buf1 gate430( .a(N1469), .O(N3003) );
inv1 gate431( .a(N1633), .O(N3006) );
buf1 gate432( .a(N1469), .O(N3007) );
buf1 gate433( .a(N1469), .O(N3010) );
and2 gate434( .a(N1315), .b(N1630), .O(N3013) );
and2 gate435( .a(N1315), .b(N1633), .O(N3014) );
inv1 gate436( .a(N1636), .O(N3015) );
inv1 gate437( .a(N1639), .O(N3016) );
inv1 gate438( .a(N1642), .O(N3017) );
inv1 gate439( .a(N1645), .O(N3018) );
inv1 gate440( .a(N1648), .O(N3019) );
inv1 gate441( .a(N1651), .O(N3020) );
inv1 gate442( .a(N1654), .O(N3021) );
inv1 gate443( .a(N1657), .O(N3022) );
and3 gate444( .a(N1303), .b(N457), .c(N1639), .O(N3023) );
and3 gate445( .a(N1303), .b(N468), .c(N1645), .O(N3024) );
and3 gate446( .a(N1303), .b(N422), .c(N1651), .O(N3025) );
and3 gate447( .a(N1303), .b(N435), .c(N1657), .O(N3026) );
and2 gate448( .a(N1663), .b(N1636), .O(N3027) );
and2 gate449( .a(N1663), .b(N1642), .O(N3028) );
and2 gate450( .a(N1663), .b(N1648), .O(N3029) );
and2 gate451( .a(N1663), .b(N1654), .O(N3030) );
inv1 gate452( .a(N1920), .O(N3031) );
inv1 gate453( .a(N1923), .O(N3032) );
inv1 gate454( .a(N1926), .O(N3033) );
inv1 gate455( .a(N1929), .O(N3034) );
buf1 gate456( .a(N1660), .O(N3035) );
buf1 gate457( .a(N1660), .O(N3038) );
inv1 gate458( .a(N1697), .O(N3041) );
inv1 gate459( .a(N1709), .O(N3052) );
inv1 gate460( .a(N1721), .O(N3063) );
inv1 gate461( .a(N1727), .O(N3068) );
and2 gate462( .a(N97), .b(N1721), .O(N3071) );
and2 gate463( .a(N94), .b(N1721), .O(N3072) );
and2 gate464( .a(N97), .b(N1721), .O(N3073) );
and2 gate465( .a(N94), .b(N1721), .O(N3074) );
inv1 gate466( .a(N1731), .O(N3075) );
inv1 gate467( .a(N1743), .O(N3086) );
inv1 gate468( .a(N1761), .O(N3097) );
inv1 gate469( .a(N1769), .O(N3108) );
inv1 gate470( .a(N1777), .O(N3119) );
inv1 gate471( .a(N1785), .O(N3130) );
inv1 gate472( .a(N1944), .O(N3141) );
inv1 gate473( .a(N1947), .O(N3142) );
inv1 gate474( .a(N1950), .O(N3143) );
inv1 gate475( .a(N1953), .O(N3144) );
inv1 gate476( .a(N1956), .O(N3145) );
inv1 gate477( .a(N1959), .O(N3146) );
inv1 gate478( .a(N1793), .O(N3147) );
inv1 gate479( .a(N1800), .O(N3158) );
inv1 gate480( .a(N1807), .O(N3169) );
inv1 gate481( .a(N1814), .O(N3180) );
buf1 gate482( .a(N1821), .O(N3191) );
inv1 gate483( .a(N1932), .O(N3194) );
inv1 gate484( .a(N1935), .O(N3195) );
inv1 gate485( .a(N1938), .O(N3196) );
inv1 gate486( .a(N1941), .O(N3197) );
inv1 gate487( .a(N1962), .O(N3198) );
inv1 gate488( .a(N1965), .O(N3199) );
buf1 gate489( .a(N1469), .O(N3200) );
inv1 gate490( .a(N1968), .O(N3203) );
buf1 gate491( .a(N2704), .O(N3357) );
buf1 gate492( .a(N2704), .O(N3358) );
buf1 gate493( .a(N2704), .O(N3359) );
buf1 gate494( .a(N2704), .O(N3360) );
and3 gate495( .a(N457), .b(N1092), .c(N2824), .O(N3401) );
and3 gate496( .a(N468), .b(N1092), .c(N2826), .O(N3402) );
and3 gate497( .a(N422), .b(N1092), .c(N2828), .O(N3403) );
and3 gate498( .a(N435), .b(N1092), .c(N2830), .O(N3404) );
and2 gate499( .a(N1080), .b(N2823), .O(N3405) );
and2 gate500( .a(N1080), .b(N2825), .O(N3406) );
and2 gate501( .a(N1080), .b(N2827), .O(N3407) );
and2 gate502( .a(N1080), .b(N2829), .O(N3408) );
and3 gate503( .a(N389), .b(N1092), .c(N2840), .O(N3409) );
and3 gate504( .a(N400), .b(N1092), .c(N2842), .O(N3410) );
and3 gate505( .a(N411), .b(N1092), .c(N2844), .O(N3411) );
and3 gate506( .a(N374), .b(N1092), .c(N2846), .O(N3412) );
and2 gate507( .a(N1080), .b(N2839), .O(N3413) );
and2 gate508( .a(N1080), .b(N2841), .O(N3414) );
and2 gate509( .a(N1080), .b(N2843), .O(N3415) );
and2 gate510( .a(N1080), .b(N2845), .O(N3416) );
and2 gate511( .a(N1280), .b(N2902), .O(N3444) );
and3 gate512( .a(N479), .b(N1280), .c(N2904), .O(N3445) );
and3 gate513( .a(N490), .b(N1280), .c(N2906), .O(N3446) );
and2 gate514( .a(N1685), .b(N2901), .O(N3447) );
and2 gate515( .a(N1685), .b(N2903), .O(N3448) );
and2 gate516( .a(N1685), .b(N2905), .O(N3449) );
and3 gate517( .a(N503), .b(N1092), .c(N2914), .O(N3450) );
and3 gate518( .a(N523), .b(N1092), .c(N2916), .O(N3451) );
and3 gate519( .a(N534), .b(N1092), .c(N2918), .O(N3452) );
and2 gate520( .a(N1080), .b(N2913), .O(N3453) );
and2 gate521( .a(N1080), .b(N2915), .O(N3454) );
and2 gate522( .a(N1080), .b(N2917), .O(N3455) );
and2 gate523( .a(N2920), .b(N2350), .O(N3456) );
and3 gate524( .a(N389), .b(N1280), .c(N2927), .O(N3459) );
and3 gate525( .a(N400), .b(N1280), .c(N2929), .O(N3460) );
and3 gate526( .a(N411), .b(N1280), .c(N2931), .O(N3461) );
and3 gate527( .a(N374), .b(N1280), .c(N2933), .O(N3462) );
and2 gate528( .a(N1685), .b(N2926), .O(N3463) );
and2 gate529( .a(N1685), .b(N2928), .O(N3464) );
and2 gate530( .a(N1685), .b(N2930), .O(N3465) );
and2 gate531( .a(N1685), .b(N2932), .O(N3466) );
and3 gate532( .a(N503), .b(N1292), .c(N2974), .O(N3481) );
inv1 gate533( .a(N2980), .O(N3482) );
and3 gate534( .a(N523), .b(N1292), .c(N2976), .O(N3483) );
and3 gate535( .a(N534), .b(N1292), .c(N2978), .O(N3484) );
and2 gate536( .a(N1271), .b(N2973), .O(N3485) );
and2 gate537( .a(N1271), .b(N2975), .O(N3486) );
and2 gate538( .a(N1271), .b(N2977), .O(N3487) );
and2 gate539( .a(N1292), .b(N2988), .O(N3488) );
and3 gate540( .a(N479), .b(N1292), .c(N2990), .O(N3489) );
and3 gate541( .a(N490), .b(N1292), .c(N2992), .O(N3490) );
and2 gate542( .a(N1271), .b(N2987), .O(N3491) );
and2 gate543( .a(N1271), .b(N2989), .O(N3492) );
and2 gate544( .a(N1271), .b(N2991), .O(N3493) );
and2 gate545( .a(N1292), .b(N2999), .O(N3502) );
and2 gate546( .a(N1292), .b(N3006), .O(N3503) );
and3 gate547( .a(N457), .b(N1280), .c(N3016), .O(N3504) );
and3 gate548( .a(N468), .b(N1280), .c(N3018), .O(N3505) );
and3 gate549( .a(N422), .b(N1280), .c(N3020), .O(N3506) );
and3 gate550( .a(N435), .b(N1280), .c(N3022), .O(N3507) );
and2 gate551( .a(N1685), .b(N3015), .O(N3508) );
and2 gate552( .a(N1685), .b(N3017), .O(N3509) );
and2 gate553( .a(N1685), .b(N3019), .O(N3510) );
and2 gate554( .a(N1685), .b(N3021), .O(N3511) );

  xor2  gate2336(.a(N3031), .b(N1923), .O(gate555inter0));
  nand2 gate2337(.a(gate555inter0), .b(s_4), .O(gate555inter1));
  and2  gate2338(.a(N3031), .b(N1923), .O(gate555inter2));
  inv1  gate2339(.a(s_4), .O(gate555inter3));
  inv1  gate2340(.a(s_5), .O(gate555inter4));
  nand2 gate2341(.a(gate555inter4), .b(gate555inter3), .O(gate555inter5));
  nor2  gate2342(.a(gate555inter5), .b(gate555inter2), .O(gate555inter6));
  inv1  gate2343(.a(N1923), .O(gate555inter7));
  inv1  gate2344(.a(N3031), .O(gate555inter8));
  nand2 gate2345(.a(gate555inter8), .b(gate555inter7), .O(gate555inter9));
  nand2 gate2346(.a(s_5), .b(gate555inter3), .O(gate555inter10));
  nor2  gate2347(.a(gate555inter10), .b(gate555inter9), .O(gate555inter11));
  nor2  gate2348(.a(gate555inter11), .b(gate555inter6), .O(gate555inter12));
  nand2 gate2349(.a(gate555inter12), .b(gate555inter1), .O(N3512));
nand2 gate556( .a(N1920), .b(N3032), .O(N3513) );

  xor2  gate3890(.a(N3033), .b(N1929), .O(gate557inter0));
  nand2 gate3891(.a(gate557inter0), .b(s_226), .O(gate557inter1));
  and2  gate3892(.a(N3033), .b(N1929), .O(gate557inter2));
  inv1  gate3893(.a(s_226), .O(gate557inter3));
  inv1  gate3894(.a(s_227), .O(gate557inter4));
  nand2 gate3895(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate3896(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate3897(.a(N1929), .O(gate557inter7));
  inv1  gate3898(.a(N3033), .O(gate557inter8));
  nand2 gate3899(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate3900(.a(s_227), .b(gate557inter3), .O(gate557inter10));
  nor2  gate3901(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate3902(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate3903(.a(gate557inter12), .b(gate557inter1), .O(N3514));

  xor2  gate3708(.a(N3034), .b(N1926), .O(gate558inter0));
  nand2 gate3709(.a(gate558inter0), .b(s_200), .O(gate558inter1));
  and2  gate3710(.a(N3034), .b(N1926), .O(gate558inter2));
  inv1  gate3711(.a(s_200), .O(gate558inter3));
  inv1  gate3712(.a(s_201), .O(gate558inter4));
  nand2 gate3713(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate3714(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate3715(.a(N1926), .O(gate558inter7));
  inv1  gate3716(.a(N3034), .O(gate558inter8));
  nand2 gate3717(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate3718(.a(s_201), .b(gate558inter3), .O(gate558inter10));
  nor2  gate3719(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate3720(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate3721(.a(gate558inter12), .b(gate558inter1), .O(N3515));

  xor2  gate3078(.a(N3141), .b(N1947), .O(gate559inter0));
  nand2 gate3079(.a(gate559inter0), .b(s_110), .O(gate559inter1));
  and2  gate3080(.a(N3141), .b(N1947), .O(gate559inter2));
  inv1  gate3081(.a(s_110), .O(gate559inter3));
  inv1  gate3082(.a(s_111), .O(gate559inter4));
  nand2 gate3083(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate3084(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate3085(.a(N1947), .O(gate559inter7));
  inv1  gate3086(.a(N3141), .O(gate559inter8));
  nand2 gate3087(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate3088(.a(s_111), .b(gate559inter3), .O(gate559inter10));
  nor2  gate3089(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate3090(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate3091(.a(gate559inter12), .b(gate559inter1), .O(N3558));
nand2 gate560( .a(N1944), .b(N3142), .O(N3559) );
nand2 gate561( .a(N1953), .b(N3143), .O(N3560) );
nand2 gate562( .a(N1950), .b(N3144), .O(N3561) );
nand2 gate563( .a(N1959), .b(N3145), .O(N3562) );
nand2 gate564( .a(N1956), .b(N3146), .O(N3563) );
buf1 gate565( .a(N3191), .O(N3604) );

  xor2  gate2322(.a(N3194), .b(N1935), .O(gate566inter0));
  nand2 gate2323(.a(gate566inter0), .b(s_2), .O(gate566inter1));
  and2  gate2324(.a(N3194), .b(N1935), .O(gate566inter2));
  inv1  gate2325(.a(s_2), .O(gate566inter3));
  inv1  gate2326(.a(s_3), .O(gate566inter4));
  nand2 gate2327(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate2328(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate2329(.a(N1935), .O(gate566inter7));
  inv1  gate2330(.a(N3194), .O(gate566inter8));
  nand2 gate2331(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate2332(.a(s_3), .b(gate566inter3), .O(gate566inter10));
  nor2  gate2333(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate2334(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate2335(.a(gate566inter12), .b(gate566inter1), .O(N3605));
nand2 gate567( .a(N1932), .b(N3195), .O(N3606) );
nand2 gate568( .a(N1941), .b(N3196), .O(N3607) );

  xor2  gate3190(.a(N3197), .b(N1938), .O(gate569inter0));
  nand2 gate3191(.a(gate569inter0), .b(s_126), .O(gate569inter1));
  and2  gate3192(.a(N3197), .b(N1938), .O(gate569inter2));
  inv1  gate3193(.a(s_126), .O(gate569inter3));
  inv1  gate3194(.a(s_127), .O(gate569inter4));
  nand2 gate3195(.a(gate569inter4), .b(gate569inter3), .O(gate569inter5));
  nor2  gate3196(.a(gate569inter5), .b(gate569inter2), .O(gate569inter6));
  inv1  gate3197(.a(N1938), .O(gate569inter7));
  inv1  gate3198(.a(N3197), .O(gate569inter8));
  nand2 gate3199(.a(gate569inter8), .b(gate569inter7), .O(gate569inter9));
  nand2 gate3200(.a(s_127), .b(gate569inter3), .O(gate569inter10));
  nor2  gate3201(.a(gate569inter10), .b(gate569inter9), .O(gate569inter11));
  nor2  gate3202(.a(gate569inter11), .b(gate569inter6), .O(gate569inter12));
  nand2 gate3203(.a(gate569inter12), .b(gate569inter1), .O(N3608));
nand2 gate570( .a(N1965), .b(N3198), .O(N3609) );

  xor2  gate2672(.a(N3199), .b(N1962), .O(gate571inter0));
  nand2 gate2673(.a(gate571inter0), .b(s_52), .O(gate571inter1));
  and2  gate2674(.a(N3199), .b(N1962), .O(gate571inter2));
  inv1  gate2675(.a(s_52), .O(gate571inter3));
  inv1  gate2676(.a(s_53), .O(gate571inter4));
  nand2 gate2677(.a(gate571inter4), .b(gate571inter3), .O(gate571inter5));
  nor2  gate2678(.a(gate571inter5), .b(gate571inter2), .O(gate571inter6));
  inv1  gate2679(.a(N1962), .O(gate571inter7));
  inv1  gate2680(.a(N3199), .O(gate571inter8));
  nand2 gate2681(.a(gate571inter8), .b(gate571inter7), .O(gate571inter9));
  nand2 gate2682(.a(s_53), .b(gate571inter3), .O(gate571inter10));
  nor2  gate2683(.a(gate571inter10), .b(gate571inter9), .O(gate571inter11));
  nor2  gate2684(.a(gate571inter11), .b(gate571inter6), .O(gate571inter12));
  nand2 gate2685(.a(gate571inter12), .b(gate571inter1), .O(N3610));
inv1 gate572( .a(N3191), .O(N3613) );
and2 gate573( .a(N2882), .b(N2891), .O(N3614) );
and2 gate574( .a(N1482), .b(N2891), .O(N3615) );
and3 gate575( .a(N200), .b(N2653), .c(N1173), .O(N3616) );
and3 gate576( .a(N203), .b(N2653), .c(N1173), .O(N3617) );
and3 gate577( .a(N197), .b(N2653), .c(N1173), .O(N3618) );
and3 gate578( .a(N194), .b(N2653), .c(N1173), .O(N3619) );
and3 gate579( .a(N191), .b(N2653), .c(N1173), .O(N3620) );
and3 gate580( .a(N182), .b(N2681), .c(N1197), .O(N3621) );
and3 gate581( .a(N188), .b(N2681), .c(N1197), .O(N3622) );
and3 gate582( .a(N155), .b(N2681), .c(N1197), .O(N3623) );
and3 gate583( .a(N149), .b(N2681), .c(N1197), .O(N3624) );
and2 gate584( .a(N2882), .b(N2891), .O(N3625) );
and2 gate585( .a(N1482), .b(N2891), .O(N3626) );
and3 gate586( .a(N200), .b(N2728), .c(N1235), .O(N3627) );
and3 gate587( .a(N203), .b(N2728), .c(N1235), .O(N3628) );
and3 gate588( .a(N197), .b(N2728), .c(N1235), .O(N3629) );
and3 gate589( .a(N194), .b(N2728), .c(N1235), .O(N3630) );
and3 gate590( .a(N191), .b(N2728), .c(N1235), .O(N3631) );
and3 gate591( .a(N182), .b(N2756), .c(N1259), .O(N3632) );
and3 gate592( .a(N188), .b(N2756), .c(N1259), .O(N3633) );
and3 gate593( .a(N155), .b(N2756), .c(N1259), .O(N3634) );
and3 gate594( .a(N149), .b(N2756), .c(N1259), .O(N3635) );
and2 gate595( .a(N2882), .b(N2891), .O(N3636) );
and2 gate596( .a(N1482), .b(N2891), .O(N3637) );
and3 gate597( .a(N109), .b(N3075), .c(N1743), .O(N3638) );
and2 gate598( .a(N2882), .b(N2891), .O(N3639) );
and2 gate599( .a(N1482), .b(N2891), .O(N3640) );
and3 gate600( .a(N11), .b(N2779), .c(N1339), .O(N3641) );
and3 gate601( .a(N109), .b(N3041), .c(N1709), .O(N3642) );
and3 gate602( .a(N46), .b(N3041), .c(N1709), .O(N3643) );
and3 gate603( .a(N100), .b(N3041), .c(N1709), .O(N3644) );
and3 gate604( .a(N91), .b(N3041), .c(N1709), .O(N3645) );
and3 gate605( .a(N43), .b(N3041), .c(N1709), .O(N3646) );
and3 gate606( .a(N76), .b(N2779), .c(N1339), .O(N3647) );
and3 gate607( .a(N73), .b(N2779), .c(N1339), .O(N3648) );
and3 gate608( .a(N67), .b(N2779), .c(N1339), .O(N3649) );
and3 gate609( .a(N14), .b(N2779), .c(N1339), .O(N3650) );
and3 gate610( .a(N46), .b(N3075), .c(N1743), .O(N3651) );
and3 gate611( .a(N100), .b(N3075), .c(N1743), .O(N3652) );
and3 gate612( .a(N91), .b(N3075), .c(N1743), .O(N3653) );
and3 gate613( .a(N43), .b(N3075), .c(N1743), .O(N3654) );
and3 gate614( .a(N76), .b(N2801), .c(N1363), .O(N3655) );
and3 gate615( .a(N73), .b(N2801), .c(N1363), .O(N3656) );
and3 gate616( .a(N67), .b(N2801), .c(N1363), .O(N3657) );
and3 gate617( .a(N14), .b(N2801), .c(N1363), .O(N3658) );
and3 gate618( .a(N120), .b(N3119), .c(N1785), .O(N3659) );
and3 gate619( .a(N11), .b(N2801), .c(N1363), .O(N3660) );
and3 gate620( .a(N118), .b(N3097), .c(N1769), .O(N3661) );
and3 gate621( .a(N176), .b(N2681), .c(N1197), .O(N3662) );
and3 gate622( .a(N176), .b(N2756), .c(N1259), .O(N3663) );
or2 gate623( .a(N2831), .b(N3401), .O(N3664) );
or2 gate624( .a(N2832), .b(N3402), .O(N3665) );
or2 gate625( .a(N2833), .b(N3403), .O(N3666) );
or2 gate626( .a(N2834), .b(N3404), .O(N3667) );
or3 gate627( .a(N2835), .b(N3405), .c(N457), .O(N3668) );
or3 gate628( .a(N2836), .b(N3406), .c(N468), .O(N3669) );
or3 gate629( .a(N2837), .b(N3407), .c(N422), .O(N3670) );
or3 gate630( .a(N2838), .b(N3408), .c(N435), .O(N3671) );
or2 gate631( .a(N2847), .b(N3409), .O(N3672) );
or2 gate632( .a(N2848), .b(N3410), .O(N3673) );
or2 gate633( .a(N2849), .b(N3411), .O(N3674) );
or2 gate634( .a(N2850), .b(N3412), .O(N3675) );
or3 gate635( .a(N2851), .b(N3413), .c(N389), .O(N3676) );
or3 gate636( .a(N2852), .b(N3414), .c(N400), .O(N3677) );
or3 gate637( .a(N2853), .b(N3415), .c(N411), .O(N3678) );
or3 gate638( .a(N2854), .b(N3416), .c(N374), .O(N3679) );
and2 gate639( .a(N289), .b(N2855), .O(N3680) );
and2 gate640( .a(N281), .b(N2855), .O(N3681) );
and2 gate641( .a(N273), .b(N2855), .O(N3682) );
and2 gate642( .a(N265), .b(N2855), .O(N3683) );
and2 gate643( .a(N257), .b(N2855), .O(N3684) );
and2 gate644( .a(N234), .b(N2861), .O(N3685) );
and2 gate645( .a(N226), .b(N2861), .O(N3686) );
and2 gate646( .a(N218), .b(N2861), .O(N3687) );
and2 gate647( .a(N210), .b(N2861), .O(N3688) );
and2 gate648( .a(N206), .b(N2861), .O(N3689) );
inv1 gate649( .a(N2891), .O(N3691) );
or2 gate650( .a(N2907), .b(N3444), .O(N3700) );
or2 gate651( .a(N2908), .b(N3445), .O(N3701) );
or2 gate652( .a(N2909), .b(N3446), .O(N3702) );
or3 gate653( .a(N2911), .b(N3448), .c(N479), .O(N3703) );
or3 gate654( .a(N2912), .b(N3449), .c(N490), .O(N3704) );
or2 gate655( .a(N2910), .b(N3447), .O(N3705) );
or2 gate656( .a(N2919), .b(N3450), .O(N3708) );
or2 gate657( .a(N2921), .b(N3451), .O(N3709) );
or2 gate658( .a(N2922), .b(N3452), .O(N3710) );
or3 gate659( .a(N2923), .b(N3453), .c(N503), .O(N3711) );
or3 gate660( .a(N2924), .b(N3454), .c(N523), .O(N3712) );
or3 gate661( .a(N2925), .b(N3455), .c(N534), .O(N3713) );
or2 gate662( .a(N2934), .b(N3459), .O(N3715) );
or2 gate663( .a(N2935), .b(N3460), .O(N3716) );
or2 gate664( .a(N2936), .b(N3461), .O(N3717) );
or2 gate665( .a(N2937), .b(N3462), .O(N3718) );
or3 gate666( .a(N2938), .b(N3463), .c(N389), .O(N3719) );
or3 gate667( .a(N2939), .b(N3464), .c(N400), .O(N3720) );
or3 gate668( .a(N2940), .b(N3465), .c(N411), .O(N3721) );
or3 gate669( .a(N2941), .b(N3466), .c(N374), .O(N3722) );
and2 gate670( .a(N369), .b(N2942), .O(N3723) );
and2 gate671( .a(N361), .b(N2942), .O(N3724) );
and2 gate672( .a(N351), .b(N2942), .O(N3725) );
and2 gate673( .a(N341), .b(N2942), .O(N3726) );
and2 gate674( .a(N324), .b(N2948), .O(N3727) );
and2 gate675( .a(N316), .b(N2948), .O(N3728) );
and2 gate676( .a(N308), .b(N2948), .O(N3729) );
and2 gate677( .a(N302), .b(N2948), .O(N3730) );
and2 gate678( .a(N293), .b(N2948), .O(N3731) );
or2 gate679( .a(N2942), .b(N2958), .O(N3732) );
and2 gate680( .a(N83), .b(N2964), .O(N3738) );
and2 gate681( .a(N87), .b(N2964), .O(N3739) );
and2 gate682( .a(N34), .b(N2964), .O(N3740) );
and2 gate683( .a(N34), .b(N2964), .O(N3741) );
or2 gate684( .a(N2979), .b(N3481), .O(N3742) );
or2 gate685( .a(N2981), .b(N3483), .O(N3743) );
or2 gate686( .a(N2982), .b(N3484), .O(N3744) );
or3 gate687( .a(N2983), .b(N3485), .c(N503), .O(N3745) );
or3 gate688( .a(N2985), .b(N3486), .c(N523), .O(N3746) );
or3 gate689( .a(N2986), .b(N3487), .c(N534), .O(N3747) );
or2 gate690( .a(N2993), .b(N3488), .O(N3748) );
or2 gate691( .a(N2994), .b(N3489), .O(N3749) );
or2 gate692( .a(N2995), .b(N3490), .O(N3750) );
or3 gate693( .a(N2997), .b(N3492), .c(N479), .O(N3751) );
or3 gate694( .a(N2998), .b(N3493), .c(N490), .O(N3752) );
inv1 gate695( .a(N3000), .O(N3753) );
inv1 gate696( .a(N3003), .O(N3754) );
inv1 gate697( .a(N3007), .O(N3755) );
inv1 gate698( .a(N3010), .O(N3756) );
or2 gate699( .a(N3013), .b(N3502), .O(N3757) );
and3 gate700( .a(N1315), .b(N446), .c(N3003), .O(N3758) );
or2 gate701( .a(N3014), .b(N3503), .O(N3759) );
and3 gate702( .a(N1315), .b(N446), .c(N3010), .O(N3760) );
and2 gate703( .a(N1675), .b(N3000), .O(N3761) );
and2 gate704( .a(N1675), .b(N3007), .O(N3762) );
or2 gate705( .a(N3023), .b(N3504), .O(N3763) );
or2 gate706( .a(N3024), .b(N3505), .O(N3764) );
or2 gate707( .a(N3025), .b(N3506), .O(N3765) );
or2 gate708( .a(N3026), .b(N3507), .O(N3766) );
or3 gate709( .a(N3027), .b(N3508), .c(N457), .O(N3767) );
or3 gate710( .a(N3028), .b(N3509), .c(N468), .O(N3768) );
or3 gate711( .a(N3029), .b(N3510), .c(N422), .O(N3769) );
or3 gate712( .a(N3030), .b(N3511), .c(N435), .O(N3770) );
nand2 gate713( .a(N3512), .b(N3513), .O(N3771) );
nand2 gate714( .a(N3514), .b(N3515), .O(N3775) );
inv1 gate715( .a(N3035), .O(N3779) );
inv1 gate716( .a(N3038), .O(N3780) );
and3 gate717( .a(N117), .b(N3097), .c(N1769), .O(N3781) );
and3 gate718( .a(N126), .b(N3097), .c(N1769), .O(N3782) );
and3 gate719( .a(N127), .b(N3097), .c(N1769), .O(N3783) );
and3 gate720( .a(N128), .b(N3097), .c(N1769), .O(N3784) );
and3 gate721( .a(N131), .b(N3119), .c(N1785), .O(N3785) );
and3 gate722( .a(N129), .b(N3119), .c(N1785), .O(N3786) );
and3 gate723( .a(N119), .b(N3119), .c(N1785), .O(N3787) );
and3 gate724( .a(N130), .b(N3119), .c(N1785), .O(N3788) );
nand2 gate725( .a(N3558), .b(N3559), .O(N3789) );
nand2 gate726( .a(N3560), .b(N3561), .O(N3793) );
nand2 gate727( .a(N3562), .b(N3563), .O(N3797) );
and3 gate728( .a(N122), .b(N3147), .c(N1800), .O(N3800) );
and3 gate729( .a(N113), .b(N3147), .c(N1800), .O(N3801) );
and3 gate730( .a(N53), .b(N3147), .c(N1800), .O(N3802) );
and3 gate731( .a(N114), .b(N3147), .c(N1800), .O(N3803) );
and3 gate732( .a(N115), .b(N3147), .c(N1800), .O(N3804) );
and3 gate733( .a(N52), .b(N3169), .c(N1814), .O(N3805) );
and3 gate734( .a(N112), .b(N3169), .c(N1814), .O(N3806) );
and3 gate735( .a(N116), .b(N3169), .c(N1814), .O(N3807) );
and3 gate736( .a(N121), .b(N3169), .c(N1814), .O(N3808) );
and3 gate737( .a(N123), .b(N3169), .c(N1814), .O(N3809) );
nand2 gate738( .a(N3607), .b(N3608), .O(N3810) );

  xor2  gate3148(.a(N3606), .b(N3605), .O(gate739inter0));
  nand2 gate3149(.a(gate739inter0), .b(s_120), .O(gate739inter1));
  and2  gate3150(.a(N3606), .b(N3605), .O(gate739inter2));
  inv1  gate3151(.a(s_120), .O(gate739inter3));
  inv1  gate3152(.a(s_121), .O(gate739inter4));
  nand2 gate3153(.a(gate739inter4), .b(gate739inter3), .O(gate739inter5));
  nor2  gate3154(.a(gate739inter5), .b(gate739inter2), .O(gate739inter6));
  inv1  gate3155(.a(N3605), .O(gate739inter7));
  inv1  gate3156(.a(N3606), .O(gate739inter8));
  nand2 gate3157(.a(gate739inter8), .b(gate739inter7), .O(gate739inter9));
  nand2 gate3158(.a(s_121), .b(gate739inter3), .O(gate739inter10));
  nor2  gate3159(.a(gate739inter10), .b(gate739inter9), .O(gate739inter11));
  nor2  gate3160(.a(gate739inter11), .b(gate739inter6), .O(gate739inter12));
  nand2 gate3161(.a(gate739inter12), .b(gate739inter1), .O(N3813));
and2 gate740( .a(N3482), .b(N2984), .O(N3816) );
or2 gate741( .a(N2996), .b(N3491), .O(N3819) );
inv1 gate742( .a(N3200), .O(N3822) );
nand2 gate743( .a(N3200), .b(N3203), .O(N3823) );

  xor2  gate3218(.a(N3610), .b(N3609), .O(gate744inter0));
  nand2 gate3219(.a(gate744inter0), .b(s_130), .O(gate744inter1));
  and2  gate3220(.a(N3610), .b(N3609), .O(gate744inter2));
  inv1  gate3221(.a(s_130), .O(gate744inter3));
  inv1  gate3222(.a(s_131), .O(gate744inter4));
  nand2 gate3223(.a(gate744inter4), .b(gate744inter3), .O(gate744inter5));
  nor2  gate3224(.a(gate744inter5), .b(gate744inter2), .O(gate744inter6));
  inv1  gate3225(.a(N3609), .O(gate744inter7));
  inv1  gate3226(.a(N3610), .O(gate744inter8));
  nand2 gate3227(.a(gate744inter8), .b(gate744inter7), .O(gate744inter9));
  nand2 gate3228(.a(s_131), .b(gate744inter3), .O(gate744inter10));
  nor2  gate3229(.a(gate744inter10), .b(gate744inter9), .O(gate744inter11));
  nor2  gate3230(.a(gate744inter11), .b(gate744inter6), .O(gate744inter12));
  nand2 gate3231(.a(gate744inter12), .b(gate744inter1), .O(N3824));
inv1 gate745( .a(N3456), .O(N3827) );
or2 gate746( .a(N3739), .b(N2970), .O(N3828) );
or2 gate747( .a(N3740), .b(N2971), .O(N3829) );
or2 gate748( .a(N3741), .b(N2972), .O(N3830) );
or2 gate749( .a(N3738), .b(N2969), .O(N3831) );
inv1 gate750( .a(N3664), .O(N3834) );
inv1 gate751( .a(N3665), .O(N3835) );
inv1 gate752( .a(N3666), .O(N3836) );
inv1 gate753( .a(N3667), .O(N3837) );
inv1 gate754( .a(N3672), .O(N3838) );
inv1 gate755( .a(N3673), .O(N3839) );
inv1 gate756( .a(N3674), .O(N3840) );
inv1 gate757( .a(N3675), .O(N3841) );
or2 gate758( .a(N3681), .b(N2868), .O(N3842) );
or2 gate759( .a(N3682), .b(N2869), .O(N3849) );
or2 gate760( .a(N3683), .b(N2870), .O(N3855) );
or2 gate761( .a(N3684), .b(N2871), .O(N3861) );
or2 gate762( .a(N3685), .b(N2872), .O(N3867) );
or2 gate763( .a(N3686), .b(N2873), .O(N3873) );
or2 gate764( .a(N3687), .b(N2874), .O(N3881) );
or2 gate765( .a(N3688), .b(N2875), .O(N3887) );
or2 gate766( .a(N3689), .b(N2876), .O(N3893) );
inv1 gate767( .a(N3701), .O(N3908) );
inv1 gate768( .a(N3702), .O(N3909) );
inv1 gate769( .a(N3700), .O(N3911) );
inv1 gate770( .a(N3708), .O(N3914) );
inv1 gate771( .a(N3709), .O(N3915) );
inv1 gate772( .a(N3710), .O(N3916) );
inv1 gate773( .a(N3715), .O(N3917) );
inv1 gate774( .a(N3716), .O(N3918) );
inv1 gate775( .a(N3717), .O(N3919) );
inv1 gate776( .a(N3718), .O(N3920) );
or2 gate777( .a(N3724), .b(N2955), .O(N3921) );
or2 gate778( .a(N3725), .b(N2956), .O(N3927) );
or2 gate779( .a(N3726), .b(N2957), .O(N3933) );
or2 gate780( .a(N3727), .b(N2959), .O(N3942) );
or2 gate781( .a(N3728), .b(N2960), .O(N3948) );
or2 gate782( .a(N3729), .b(N2961), .O(N3956) );
or2 gate783( .a(N3730), .b(N2962), .O(N3962) );
or2 gate784( .a(N3731), .b(N2963), .O(N3968) );
inv1 gate785( .a(N3742), .O(N3975) );
inv1 gate786( .a(N3743), .O(N3976) );
inv1 gate787( .a(N3744), .O(N3977) );
inv1 gate788( .a(N3749), .O(N3978) );
inv1 gate789( .a(N3750), .O(N3979) );
and3 gate790( .a(N446), .b(N1292), .c(N3754), .O(N3980) );
and3 gate791( .a(N446), .b(N1292), .c(N3756), .O(N3981) );
and2 gate792( .a(N1271), .b(N3753), .O(N3982) );
and2 gate793( .a(N1271), .b(N3755), .O(N3983) );
inv1 gate794( .a(N3757), .O(N3984) );
inv1 gate795( .a(N3759), .O(N3987) );
inv1 gate796( .a(N3763), .O(N3988) );
inv1 gate797( .a(N3764), .O(N3989) );
inv1 gate798( .a(N3765), .O(N3990) );
inv1 gate799( .a(N3766), .O(N3991) );
and3 gate800( .a(N3456), .b(N3119), .c(N3130), .O(N3998) );
or2 gate801( .a(N3723), .b(N2954), .O(N4008) );
or2 gate802( .a(N3680), .b(N2867), .O(N4011) );
inv1 gate803( .a(N3748), .O(N4021) );
nand2 gate804( .a(N1968), .b(N3822), .O(N4024) );
inv1 gate805( .a(N3705), .O(N4027) );
and2 gate806( .a(N3828), .b(N1583), .O(N4031) );
and3 gate807( .a(N24), .b(N2882), .c(N3691), .O(N4032) );
and3 gate808( .a(N25), .b(N1482), .c(N3691), .O(N4033) );
and3 gate809( .a(N26), .b(N2882), .c(N3691), .O(N4034) );
and3 gate810( .a(N81), .b(N1482), .c(N3691), .O(N4035) );
and2 gate811( .a(N3829), .b(N1583), .O(N4036) );
and3 gate812( .a(N79), .b(N2882), .c(N3691), .O(N4037) );
and3 gate813( .a(N23), .b(N1482), .c(N3691), .O(N4038) );
and3 gate814( .a(N82), .b(N2882), .c(N3691), .O(N4039) );
and3 gate815( .a(N80), .b(N1482), .c(N3691), .O(N4040) );
and2 gate816( .a(N3830), .b(N1583), .O(N4041) );
and2 gate817( .a(N3831), .b(N1583), .O(N4042) );
and2 gate818( .a(N3732), .b(N514), .O(N4067) );
and2 gate819( .a(N514), .b(N3732), .O(N4080) );
and2 gate820( .a(N3834), .b(N3668), .O(N4088) );
and2 gate821( .a(N3835), .b(N3669), .O(N4091) );
and2 gate822( .a(N3836), .b(N3670), .O(N4094) );
and2 gate823( .a(N3837), .b(N3671), .O(N4097) );
and2 gate824( .a(N3838), .b(N3676), .O(N4100) );
and2 gate825( .a(N3839), .b(N3677), .O(N4103) );
and2 gate826( .a(N3840), .b(N3678), .O(N4106) );
and2 gate827( .a(N3841), .b(N3679), .O(N4109) );
and2 gate828( .a(N3908), .b(N3703), .O(N4144) );
and2 gate829( .a(N3909), .b(N3704), .O(N4147) );
buf1 gate830( .a(N3705), .O(N4150) );
and2 gate831( .a(N3914), .b(N3711), .O(N4153) );
and2 gate832( .a(N3915), .b(N3712), .O(N4156) );
and2 gate833( .a(N3916), .b(N3713), .O(N4159) );
or2 gate834( .a(N3758), .b(N3980), .O(N4183) );
or2 gate835( .a(N3760), .b(N3981), .O(N4184) );
or3 gate836( .a(N3761), .b(N3982), .c(N446), .O(N4185) );
or3 gate837( .a(N3762), .b(N3983), .c(N446), .O(N4186) );
inv1 gate838( .a(N3771), .O(N4188) );
inv1 gate839( .a(N3775), .O(N4191) );
and3 gate840( .a(N3775), .b(N3771), .c(N3035), .O(N4196) );
and3 gate841( .a(N3987), .b(N3119), .c(N3130), .O(N4197) );
and2 gate842( .a(N3920), .b(N3722), .O(N4198) );
inv1 gate843( .a(N3816), .O(N4199) );
inv1 gate844( .a(N3789), .O(N4200) );
inv1 gate845( .a(N3793), .O(N4203) );
buf1 gate846( .a(N3797), .O(N4206) );
buf1 gate847( .a(N3797), .O(N4209) );
buf1 gate848( .a(N3732), .O(N4212) );
buf1 gate849( .a(N3732), .O(N4215) );
buf1 gate850( .a(N3732), .O(N4219) );
inv1 gate851( .a(N3810), .O(N4223) );
inv1 gate852( .a(N3813), .O(N4224) );
and2 gate853( .a(N3918), .b(N3720), .O(N4225) );
and2 gate854( .a(N3919), .b(N3721), .O(N4228) );
and2 gate855( .a(N3991), .b(N3770), .O(N4231) );
and2 gate856( .a(N3917), .b(N3719), .O(N4234) );
and2 gate857( .a(N3989), .b(N3768), .O(N4237) );
and2 gate858( .a(N3990), .b(N3769), .O(N4240) );
and2 gate859( .a(N3988), .b(N3767), .O(N4243) );
and2 gate860( .a(N3976), .b(N3746), .O(N4246) );
and2 gate861( .a(N3977), .b(N3747), .O(N4249) );
and2 gate862( .a(N3975), .b(N3745), .O(N4252) );
and2 gate863( .a(N3978), .b(N3751), .O(N4255) );
and2 gate864( .a(N3979), .b(N3752), .O(N4258) );
inv1 gate865( .a(N3819), .O(N4263) );

  xor2  gate2742(.a(N3823), .b(N4024), .O(gate866inter0));
  nand2 gate2743(.a(gate866inter0), .b(s_62), .O(gate866inter1));
  and2  gate2744(.a(N3823), .b(N4024), .O(gate866inter2));
  inv1  gate2745(.a(s_62), .O(gate866inter3));
  inv1  gate2746(.a(s_63), .O(gate866inter4));
  nand2 gate2747(.a(gate866inter4), .b(gate866inter3), .O(gate866inter5));
  nor2  gate2748(.a(gate866inter5), .b(gate866inter2), .O(gate866inter6));
  inv1  gate2749(.a(N4024), .O(gate866inter7));
  inv1  gate2750(.a(N3823), .O(gate866inter8));
  nand2 gate2751(.a(gate866inter8), .b(gate866inter7), .O(gate866inter9));
  nand2 gate2752(.a(s_63), .b(gate866inter3), .O(gate866inter10));
  nor2  gate2753(.a(gate866inter10), .b(gate866inter9), .O(gate866inter11));
  nor2  gate2754(.a(gate866inter11), .b(gate866inter6), .O(gate866inter12));
  nand2 gate2755(.a(gate866inter12), .b(gate866inter1), .O(N4264));
inv1 gate867( .a(N3824), .O(N4267) );
and2 gate868( .a(N446), .b(N3893), .O(N4268) );
inv1 gate869( .a(N3911), .O(N4269) );
inv1 gate870( .a(N3984), .O(N4270) );
and2 gate871( .a(N3893), .b(N446), .O(N4271) );
inv1 gate872( .a(N4031), .O(N4272) );
or4 gate873( .a(N4032), .b(N4033), .c(N3614), .d(N3615), .O(N4273) );
or4 gate874( .a(N4034), .b(N4035), .c(N3625), .d(N3626), .O(N4274) );
inv1 gate875( .a(N4036), .O(N4275) );
or4 gate876( .a(N4037), .b(N4038), .c(N3636), .d(N3637), .O(N4276) );
or4 gate877( .a(N4039), .b(N4040), .c(N3639), .d(N3640), .O(N4277) );
inv1 gate878( .a(N4041), .O(N4278) );
inv1 gate879( .a(N4042), .O(N4279) );
and2 gate880( .a(N3887), .b(N457), .O(N4280) );
and2 gate881( .a(N3881), .b(N468), .O(N4284) );
and2 gate882( .a(N422), .b(N3873), .O(N4290) );
and2 gate883( .a(N3867), .b(N435), .O(N4297) );
and2 gate884( .a(N3861), .b(N389), .O(N4298) );
and2 gate885( .a(N3855), .b(N400), .O(N4301) );
and2 gate886( .a(N3849), .b(N411), .O(N4305) );
and2 gate887( .a(N3842), .b(N374), .O(N4310) );
and2 gate888( .a(N457), .b(N3887), .O(N4316) );
and2 gate889( .a(N468), .b(N3881), .O(N4320) );
and2 gate890( .a(N422), .b(N3873), .O(N4325) );
and2 gate891( .a(N435), .b(N3867), .O(N4331) );
and2 gate892( .a(N389), .b(N3861), .O(N4332) );
and2 gate893( .a(N400), .b(N3855), .O(N4336) );
and2 gate894( .a(N411), .b(N3849), .O(N4342) );
and2 gate895( .a(N374), .b(N3842), .O(N4349) );
inv1 gate896( .a(N3968), .O(N4357) );
inv1 gate897( .a(N3962), .O(N4364) );
buf1 gate898( .a(N3962), .O(N4375) );
and2 gate899( .a(N3956), .b(N479), .O(N4379) );
and2 gate900( .a(N490), .b(N3948), .O(N4385) );
and2 gate901( .a(N3942), .b(N503), .O(N4392) );
and2 gate902( .a(N3933), .b(N523), .O(N4396) );
and2 gate903( .a(N3927), .b(N534), .O(N4400) );
inv1 gate904( .a(N3921), .O(N4405) );
buf1 gate905( .a(N3921), .O(N4412) );
inv1 gate906( .a(N3968), .O(N4418) );
inv1 gate907( .a(N3962), .O(N4425) );
buf1 gate908( .a(N3962), .O(N4436) );
and2 gate909( .a(N479), .b(N3956), .O(N4440) );
and2 gate910( .a(N490), .b(N3948), .O(N4445) );
and2 gate911( .a(N503), .b(N3942), .O(N4451) );
and2 gate912( .a(N523), .b(N3933), .O(N4456) );
and2 gate913( .a(N534), .b(N3927), .O(N4462) );
buf1 gate914( .a(N3921), .O(N4469) );
inv1 gate915( .a(N3921), .O(N4477) );
buf1 gate916( .a(N3968), .O(N4512) );
inv1 gate917( .a(N4183), .O(N4515) );
inv1 gate918( .a(N4184), .O(N4516) );
inv1 gate919( .a(N4008), .O(N4521) );
inv1 gate920( .a(N4011), .O(N4523) );
inv1 gate921( .a(N4198), .O(N4524) );
inv1 gate922( .a(N3984), .O(N4532) );
and3 gate923( .a(N3911), .b(N3169), .c(N3180), .O(N4547) );
buf1 gate924( .a(N3893), .O(N4548) );
buf1 gate925( .a(N3887), .O(N4551) );
buf1 gate926( .a(N3881), .O(N4554) );
buf1 gate927( .a(N3873), .O(N4557) );
buf1 gate928( .a(N3867), .O(N4560) );
buf1 gate929( .a(N3861), .O(N4563) );
buf1 gate930( .a(N3855), .O(N4566) );
buf1 gate931( .a(N3849), .O(N4569) );
buf1 gate932( .a(N3842), .O(N4572) );
nor2 gate933( .a(N422), .b(N3873), .O(N4575) );
buf1 gate934( .a(N3893), .O(N4578) );
buf1 gate935( .a(N3887), .O(N4581) );
buf1 gate936( .a(N3881), .O(N4584) );
buf1 gate937( .a(N3867), .O(N4587) );
buf1 gate938( .a(N3861), .O(N4590) );
buf1 gate939( .a(N3855), .O(N4593) );
buf1 gate940( .a(N3849), .O(N4596) );
buf1 gate941( .a(N3873), .O(N4599) );
buf1 gate942( .a(N3842), .O(N4602) );
nor2 gate943( .a(N422), .b(N3873), .O(N4605) );
nor2 gate944( .a(N374), .b(N3842), .O(N4608) );
buf1 gate945( .a(N3956), .O(N4611) );
buf1 gate946( .a(N3948), .O(N4614) );
buf1 gate947( .a(N3942), .O(N4617) );
buf1 gate948( .a(N3933), .O(N4621) );
buf1 gate949( .a(N3927), .O(N4624) );
nor2 gate950( .a(N490), .b(N3948), .O(N4627) );
buf1 gate951( .a(N3956), .O(N4630) );
buf1 gate952( .a(N3942), .O(N4633) );
buf1 gate953( .a(N3933), .O(N4637) );
buf1 gate954( .a(N3927), .O(N4640) );
buf1 gate955( .a(N3948), .O(N4643) );
nor2 gate956( .a(N490), .b(N3948), .O(N4646) );
buf1 gate957( .a(N3927), .O(N4649) );
buf1 gate958( .a(N3933), .O(N4652) );
buf1 gate959( .a(N3921), .O(N4655) );
buf1 gate960( .a(N3942), .O(N4658) );
buf1 gate961( .a(N3956), .O(N4662) );
buf1 gate962( .a(N3948), .O(N4665) );
buf1 gate963( .a(N3968), .O(N4668) );
buf1 gate964( .a(N3962), .O(N4671) );
buf1 gate965( .a(N3873), .O(N4674) );
buf1 gate966( .a(N3867), .O(N4677) );
buf1 gate967( .a(N3887), .O(N4680) );
buf1 gate968( .a(N3881), .O(N4683) );
buf1 gate969( .a(N3893), .O(N4686) );
buf1 gate970( .a(N3849), .O(N4689) );
buf1 gate971( .a(N3842), .O(N4692) );
buf1 gate972( .a(N3861), .O(N4695) );
buf1 gate973( .a(N3855), .O(N4698) );
nand2 gate974( .a(N3813), .b(N4223), .O(N4701) );

  xor2  gate3750(.a(N4224), .b(N3810), .O(gate975inter0));
  nand2 gate3751(.a(gate975inter0), .b(s_206), .O(gate975inter1));
  and2  gate3752(.a(N4224), .b(N3810), .O(gate975inter2));
  inv1  gate3753(.a(s_206), .O(gate975inter3));
  inv1  gate3754(.a(s_207), .O(gate975inter4));
  nand2 gate3755(.a(gate975inter4), .b(gate975inter3), .O(gate975inter5));
  nor2  gate3756(.a(gate975inter5), .b(gate975inter2), .O(gate975inter6));
  inv1  gate3757(.a(N3810), .O(gate975inter7));
  inv1  gate3758(.a(N4224), .O(gate975inter8));
  nand2 gate3759(.a(gate975inter8), .b(gate975inter7), .O(gate975inter9));
  nand2 gate3760(.a(s_207), .b(gate975inter3), .O(gate975inter10));
  nor2  gate3761(.a(gate975inter10), .b(gate975inter9), .O(gate975inter11));
  nor2  gate3762(.a(gate975inter11), .b(gate975inter6), .O(gate975inter12));
  nand2 gate3763(.a(gate975inter12), .b(gate975inter1), .O(N4702));
inv1 gate976( .a(N4021), .O(N4720) );

  xor2  gate2490(.a(N4263), .b(N4021), .O(gate977inter0));
  nand2 gate2491(.a(gate977inter0), .b(s_26), .O(gate977inter1));
  and2  gate2492(.a(N4263), .b(N4021), .O(gate977inter2));
  inv1  gate2493(.a(s_26), .O(gate977inter3));
  inv1  gate2494(.a(s_27), .O(gate977inter4));
  nand2 gate2495(.a(gate977inter4), .b(gate977inter3), .O(gate977inter5));
  nor2  gate2496(.a(gate977inter5), .b(gate977inter2), .O(gate977inter6));
  inv1  gate2497(.a(N4021), .O(gate977inter7));
  inv1  gate2498(.a(N4263), .O(gate977inter8));
  nand2 gate2499(.a(gate977inter8), .b(gate977inter7), .O(gate977inter9));
  nand2 gate2500(.a(s_27), .b(gate977inter3), .O(gate977inter10));
  nor2  gate2501(.a(gate977inter10), .b(gate977inter9), .O(gate977inter11));
  nor2  gate2502(.a(gate977inter11), .b(gate977inter6), .O(gate977inter12));
  nand2 gate2503(.a(gate977inter12), .b(gate977inter1), .O(N4721));
inv1 gate978( .a(N4147), .O(N4724) );
inv1 gate979( .a(N4144), .O(N4725) );
inv1 gate980( .a(N4159), .O(N4726) );
inv1 gate981( .a(N4156), .O(N4727) );
inv1 gate982( .a(N4153), .O(N4728) );
inv1 gate983( .a(N4097), .O(N4729) );
inv1 gate984( .a(N4094), .O(N4730) );
inv1 gate985( .a(N4091), .O(N4731) );
inv1 gate986( .a(N4088), .O(N4732) );
inv1 gate987( .a(N4109), .O(N4733) );
inv1 gate988( .a(N4106), .O(N4734) );
inv1 gate989( .a(N4103), .O(N4735) );
inv1 gate990( .a(N4100), .O(N4736) );
and2 gate991( .a(N4273), .b(N2877), .O(N4737) );
and2 gate992( .a(N4274), .b(N2877), .O(N4738) );
and2 gate993( .a(N4276), .b(N2877), .O(N4739) );
and2 gate994( .a(N4277), .b(N2877), .O(N4740) );
and3 gate995( .a(N4150), .b(N1758), .c(N1755), .O(N4741) );
inv1 gate996( .a(N4212), .O(N4855) );
nand2 gate997( .a(N4212), .b(N2712), .O(N4856) );
nand2 gate998( .a(N4215), .b(N2718), .O(N4908) );
inv1 gate999( .a(N4215), .O(N4909) );
and2 gate1000( .a(N4515), .b(N4185), .O(N4939) );
and2 gate1001( .a(N4516), .b(N4186), .O(N4942) );
inv1 gate1002( .a(N4219), .O(N4947) );
and3 gate1003( .a(N4188), .b(N3775), .c(N3779), .O(N4953) );
and3 gate1004( .a(N3771), .b(N4191), .c(N3780), .O(N4954) );
and3 gate1005( .a(N4191), .b(N4188), .c(N3038), .O(N4955) );
and3 gate1006( .a(N4109), .b(N3097), .c(N3108), .O(N4956) );
and3 gate1007( .a(N4106), .b(N3097), .c(N3108), .O(N4957) );
and3 gate1008( .a(N4103), .b(N3097), .c(N3108), .O(N4958) );
and3 gate1009( .a(N4100), .b(N3097), .c(N3108), .O(N4959) );
and3 gate1010( .a(N4159), .b(N3119), .c(N3130), .O(N4960) );
and3 gate1011( .a(N4156), .b(N3119), .c(N3130), .O(N4961) );
inv1 gate1012( .a(N4225), .O(N4965) );
inv1 gate1013( .a(N4228), .O(N4966) );
inv1 gate1014( .a(N4231), .O(N4967) );
inv1 gate1015( .a(N4234), .O(N4968) );
inv1 gate1016( .a(N4246), .O(N4972) );
inv1 gate1017( .a(N4249), .O(N4973) );
inv1 gate1018( .a(N4252), .O(N4974) );
nand2 gate1019( .a(N4252), .b(N4199), .O(N4975) );
inv1 gate1020( .a(N4206), .O(N4976) );
inv1 gate1021( .a(N4209), .O(N4977) );
and3 gate1022( .a(N3793), .b(N3789), .c(N4206), .O(N4978) );
and3 gate1023( .a(N4203), .b(N4200), .c(N4209), .O(N4979) );
and3 gate1024( .a(N4097), .b(N3147), .c(N3158), .O(N4980) );
and3 gate1025( .a(N4094), .b(N3147), .c(N3158), .O(N4981) );
and3 gate1026( .a(N4091), .b(N3147), .c(N3158), .O(N4982) );
and3 gate1027( .a(N4088), .b(N3147), .c(N3158), .O(N4983) );
and3 gate1028( .a(N4153), .b(N3169), .c(N3180), .O(N4984) );
and3 gate1029( .a(N4147), .b(N3169), .c(N3180), .O(N4985) );
and3 gate1030( .a(N4144), .b(N3169), .c(N3180), .O(N4986) );
and3 gate1031( .a(N4150), .b(N3169), .c(N3180), .O(N4987) );
nand2 gate1032( .a(N4701), .b(N4702), .O(N5049) );
inv1 gate1033( .a(N4237), .O(N5052) );
inv1 gate1034( .a(N4240), .O(N5053) );
inv1 gate1035( .a(N4243), .O(N5054) );
inv1 gate1036( .a(N4255), .O(N5055) );
inv1 gate1037( .a(N4258), .O(N5056) );

  xor2  gate3526(.a(N4720), .b(N3819), .O(gate1038inter0));
  nand2 gate3527(.a(gate1038inter0), .b(s_174), .O(gate1038inter1));
  and2  gate3528(.a(N4720), .b(N3819), .O(gate1038inter2));
  inv1  gate3529(.a(s_174), .O(gate1038inter3));
  inv1  gate3530(.a(s_175), .O(gate1038inter4));
  nand2 gate3531(.a(gate1038inter4), .b(gate1038inter3), .O(gate1038inter5));
  nor2  gate3532(.a(gate1038inter5), .b(gate1038inter2), .O(gate1038inter6));
  inv1  gate3533(.a(N3819), .O(gate1038inter7));
  inv1  gate3534(.a(N4720), .O(gate1038inter8));
  nand2 gate3535(.a(gate1038inter8), .b(gate1038inter7), .O(gate1038inter9));
  nand2 gate3536(.a(s_175), .b(gate1038inter3), .O(gate1038inter10));
  nor2  gate3537(.a(gate1038inter10), .b(gate1038inter9), .O(gate1038inter11));
  nor2  gate3538(.a(gate1038inter11), .b(gate1038inter6), .O(gate1038inter12));
  nand2 gate3539(.a(gate1038inter12), .b(gate1038inter1), .O(N5057));
inv1 gate1039( .a(N4264), .O(N5058) );
nand2 gate1040( .a(N4264), .b(N4267), .O(N5059) );
and4 gate1041( .a(N4724), .b(N4725), .c(N4269), .d(N4027), .O(N5060) );
and4 gate1042( .a(N4726), .b(N4727), .c(N3827), .d(N4728), .O(N5061) );
and4 gate1043( .a(N4729), .b(N4730), .c(N4731), .d(N4732), .O(N5062) );
and4 gate1044( .a(N4733), .b(N4734), .c(N4735), .d(N4736), .O(N5063) );
and2 gate1045( .a(N4357), .b(N4375), .O(N5065) );
and3 gate1046( .a(N4364), .b(N4357), .c(N4379), .O(N5066) );
and2 gate1047( .a(N4418), .b(N4436), .O(N5067) );
and3 gate1048( .a(N4425), .b(N4418), .c(N4440), .O(N5068) );
inv1 gate1049( .a(N4548), .O(N5069) );

  xor2  gate3736(.a(N2628), .b(N4548), .O(gate1050inter0));
  nand2 gate3737(.a(gate1050inter0), .b(s_204), .O(gate1050inter1));
  and2  gate3738(.a(N2628), .b(N4548), .O(gate1050inter2));
  inv1  gate3739(.a(s_204), .O(gate1050inter3));
  inv1  gate3740(.a(s_205), .O(gate1050inter4));
  nand2 gate3741(.a(gate1050inter4), .b(gate1050inter3), .O(gate1050inter5));
  nor2  gate3742(.a(gate1050inter5), .b(gate1050inter2), .O(gate1050inter6));
  inv1  gate3743(.a(N4548), .O(gate1050inter7));
  inv1  gate3744(.a(N2628), .O(gate1050inter8));
  nand2 gate3745(.a(gate1050inter8), .b(gate1050inter7), .O(gate1050inter9));
  nand2 gate3746(.a(s_205), .b(gate1050inter3), .O(gate1050inter10));
  nor2  gate3747(.a(gate1050inter10), .b(gate1050inter9), .O(gate1050inter11));
  nor2  gate3748(.a(gate1050inter11), .b(gate1050inter6), .O(gate1050inter12));
  nand2 gate3749(.a(gate1050inter12), .b(gate1050inter1), .O(N5070));
inv1 gate1051( .a(N4551), .O(N5071) );
nand2 gate1052( .a(N4551), .b(N2629), .O(N5072) );
inv1 gate1053( .a(N4554), .O(N5073) );
nand2 gate1054( .a(N4554), .b(N2630), .O(N5074) );
inv1 gate1055( .a(N4557), .O(N5075) );

  xor2  gate2644(.a(N2631), .b(N4557), .O(gate1056inter0));
  nand2 gate2645(.a(gate1056inter0), .b(s_48), .O(gate1056inter1));
  and2  gate2646(.a(N2631), .b(N4557), .O(gate1056inter2));
  inv1  gate2647(.a(s_48), .O(gate1056inter3));
  inv1  gate2648(.a(s_49), .O(gate1056inter4));
  nand2 gate2649(.a(gate1056inter4), .b(gate1056inter3), .O(gate1056inter5));
  nor2  gate2650(.a(gate1056inter5), .b(gate1056inter2), .O(gate1056inter6));
  inv1  gate2651(.a(N4557), .O(gate1056inter7));
  inv1  gate2652(.a(N2631), .O(gate1056inter8));
  nand2 gate2653(.a(gate1056inter8), .b(gate1056inter7), .O(gate1056inter9));
  nand2 gate2654(.a(s_49), .b(gate1056inter3), .O(gate1056inter10));
  nor2  gate2655(.a(gate1056inter10), .b(gate1056inter9), .O(gate1056inter11));
  nor2  gate2656(.a(gate1056inter11), .b(gate1056inter6), .O(gate1056inter12));
  nand2 gate2657(.a(gate1056inter12), .b(gate1056inter1), .O(N5076));
inv1 gate1057( .a(N4560), .O(N5077) );

  xor2  gate2938(.a(N2632), .b(N4560), .O(gate1058inter0));
  nand2 gate2939(.a(gate1058inter0), .b(s_90), .O(gate1058inter1));
  and2  gate2940(.a(N2632), .b(N4560), .O(gate1058inter2));
  inv1  gate2941(.a(s_90), .O(gate1058inter3));
  inv1  gate2942(.a(s_91), .O(gate1058inter4));
  nand2 gate2943(.a(gate1058inter4), .b(gate1058inter3), .O(gate1058inter5));
  nor2  gate2944(.a(gate1058inter5), .b(gate1058inter2), .O(gate1058inter6));
  inv1  gate2945(.a(N4560), .O(gate1058inter7));
  inv1  gate2946(.a(N2632), .O(gate1058inter8));
  nand2 gate2947(.a(gate1058inter8), .b(gate1058inter7), .O(gate1058inter9));
  nand2 gate2948(.a(s_91), .b(gate1058inter3), .O(gate1058inter10));
  nor2  gate2949(.a(gate1058inter10), .b(gate1058inter9), .O(gate1058inter11));
  nor2  gate2950(.a(gate1058inter11), .b(gate1058inter6), .O(gate1058inter12));
  nand2 gate2951(.a(gate1058inter12), .b(gate1058inter1), .O(N5078));
inv1 gate1059( .a(N4563), .O(N5079) );
nand2 gate1060( .a(N4563), .b(N2633), .O(N5080) );
inv1 gate1061( .a(N4566), .O(N5081) );

  xor2  gate3302(.a(N2634), .b(N4566), .O(gate1062inter0));
  nand2 gate3303(.a(gate1062inter0), .b(s_142), .O(gate1062inter1));
  and2  gate3304(.a(N2634), .b(N4566), .O(gate1062inter2));
  inv1  gate3305(.a(s_142), .O(gate1062inter3));
  inv1  gate3306(.a(s_143), .O(gate1062inter4));
  nand2 gate3307(.a(gate1062inter4), .b(gate1062inter3), .O(gate1062inter5));
  nor2  gate3308(.a(gate1062inter5), .b(gate1062inter2), .O(gate1062inter6));
  inv1  gate3309(.a(N4566), .O(gate1062inter7));
  inv1  gate3310(.a(N2634), .O(gate1062inter8));
  nand2 gate3311(.a(gate1062inter8), .b(gate1062inter7), .O(gate1062inter9));
  nand2 gate3312(.a(s_143), .b(gate1062inter3), .O(gate1062inter10));
  nor2  gate3313(.a(gate1062inter10), .b(gate1062inter9), .O(gate1062inter11));
  nor2  gate3314(.a(gate1062inter11), .b(gate1062inter6), .O(gate1062inter12));
  nand2 gate3315(.a(gate1062inter12), .b(gate1062inter1), .O(N5082));
inv1 gate1063( .a(N4569), .O(N5083) );
nand2 gate1064( .a(N4569), .b(N2635), .O(N5084) );
inv1 gate1065( .a(N4572), .O(N5085) );
nand2 gate1066( .a(N4572), .b(N2636), .O(N5086) );
inv1 gate1067( .a(N4575), .O(N5087) );

  xor2  gate3792(.a(N2638), .b(N4578), .O(gate1068inter0));
  nand2 gate3793(.a(gate1068inter0), .b(s_212), .O(gate1068inter1));
  and2  gate3794(.a(N2638), .b(N4578), .O(gate1068inter2));
  inv1  gate3795(.a(s_212), .O(gate1068inter3));
  inv1  gate3796(.a(s_213), .O(gate1068inter4));
  nand2 gate3797(.a(gate1068inter4), .b(gate1068inter3), .O(gate1068inter5));
  nor2  gate3798(.a(gate1068inter5), .b(gate1068inter2), .O(gate1068inter6));
  inv1  gate3799(.a(N4578), .O(gate1068inter7));
  inv1  gate3800(.a(N2638), .O(gate1068inter8));
  nand2 gate3801(.a(gate1068inter8), .b(gate1068inter7), .O(gate1068inter9));
  nand2 gate3802(.a(s_213), .b(gate1068inter3), .O(gate1068inter10));
  nor2  gate3803(.a(gate1068inter10), .b(gate1068inter9), .O(gate1068inter11));
  nor2  gate3804(.a(gate1068inter11), .b(gate1068inter6), .O(gate1068inter12));
  nand2 gate3805(.a(gate1068inter12), .b(gate1068inter1), .O(N5088));
inv1 gate1069( .a(N4578), .O(N5089) );
nand2 gate1070( .a(N4581), .b(N2639), .O(N5090) );
inv1 gate1071( .a(N4581), .O(N5091) );
nand2 gate1072( .a(N4584), .b(N2640), .O(N5092) );
inv1 gate1073( .a(N4584), .O(N5093) );
nand2 gate1074( .a(N4587), .b(N2641), .O(N5094) );
inv1 gate1075( .a(N4587), .O(N5095) );
nand2 gate1076( .a(N4590), .b(N2642), .O(N5096) );
inv1 gate1077( .a(N4590), .O(N5097) );

  xor2  gate2812(.a(N2643), .b(N4593), .O(gate1078inter0));
  nand2 gate2813(.a(gate1078inter0), .b(s_72), .O(gate1078inter1));
  and2  gate2814(.a(N2643), .b(N4593), .O(gate1078inter2));
  inv1  gate2815(.a(s_72), .O(gate1078inter3));
  inv1  gate2816(.a(s_73), .O(gate1078inter4));
  nand2 gate2817(.a(gate1078inter4), .b(gate1078inter3), .O(gate1078inter5));
  nor2  gate2818(.a(gate1078inter5), .b(gate1078inter2), .O(gate1078inter6));
  inv1  gate2819(.a(N4593), .O(gate1078inter7));
  inv1  gate2820(.a(N2643), .O(gate1078inter8));
  nand2 gate2821(.a(gate1078inter8), .b(gate1078inter7), .O(gate1078inter9));
  nand2 gate2822(.a(s_73), .b(gate1078inter3), .O(gate1078inter10));
  nor2  gate2823(.a(gate1078inter10), .b(gate1078inter9), .O(gate1078inter11));
  nor2  gate2824(.a(gate1078inter11), .b(gate1078inter6), .O(gate1078inter12));
  nand2 gate2825(.a(gate1078inter12), .b(gate1078inter1), .O(N5098));
inv1 gate1079( .a(N4593), .O(N5099) );
nand2 gate1080( .a(N4596), .b(N2644), .O(N5100) );
inv1 gate1081( .a(N4596), .O(N5101) );
nand2 gate1082( .a(N4599), .b(N2645), .O(N5102) );
inv1 gate1083( .a(N4599), .O(N5103) );
nand2 gate1084( .a(N4602), .b(N2646), .O(N5104) );
inv1 gate1085( .a(N4602), .O(N5105) );
inv1 gate1086( .a(N4611), .O(N5106) );

  xor2  gate2378(.a(N2709), .b(N4611), .O(gate1087inter0));
  nand2 gate2379(.a(gate1087inter0), .b(s_10), .O(gate1087inter1));
  and2  gate2380(.a(N2709), .b(N4611), .O(gate1087inter2));
  inv1  gate2381(.a(s_10), .O(gate1087inter3));
  inv1  gate2382(.a(s_11), .O(gate1087inter4));
  nand2 gate2383(.a(gate1087inter4), .b(gate1087inter3), .O(gate1087inter5));
  nor2  gate2384(.a(gate1087inter5), .b(gate1087inter2), .O(gate1087inter6));
  inv1  gate2385(.a(N4611), .O(gate1087inter7));
  inv1  gate2386(.a(N2709), .O(gate1087inter8));
  nand2 gate2387(.a(gate1087inter8), .b(gate1087inter7), .O(gate1087inter9));
  nand2 gate2388(.a(s_11), .b(gate1087inter3), .O(gate1087inter10));
  nor2  gate2389(.a(gate1087inter10), .b(gate1087inter9), .O(gate1087inter11));
  nor2  gate2390(.a(gate1087inter11), .b(gate1087inter6), .O(gate1087inter12));
  nand2 gate2391(.a(gate1087inter12), .b(gate1087inter1), .O(N5107));
inv1 gate1088( .a(N4614), .O(N5108) );

  xor2  gate3596(.a(N2710), .b(N4614), .O(gate1089inter0));
  nand2 gate3597(.a(gate1089inter0), .b(s_184), .O(gate1089inter1));
  and2  gate3598(.a(N2710), .b(N4614), .O(gate1089inter2));
  inv1  gate3599(.a(s_184), .O(gate1089inter3));
  inv1  gate3600(.a(s_185), .O(gate1089inter4));
  nand2 gate3601(.a(gate1089inter4), .b(gate1089inter3), .O(gate1089inter5));
  nor2  gate3602(.a(gate1089inter5), .b(gate1089inter2), .O(gate1089inter6));
  inv1  gate3603(.a(N4614), .O(gate1089inter7));
  inv1  gate3604(.a(N2710), .O(gate1089inter8));
  nand2 gate3605(.a(gate1089inter8), .b(gate1089inter7), .O(gate1089inter9));
  nand2 gate3606(.a(s_185), .b(gate1089inter3), .O(gate1089inter10));
  nor2  gate3607(.a(gate1089inter10), .b(gate1089inter9), .O(gate1089inter11));
  nor2  gate3608(.a(gate1089inter11), .b(gate1089inter6), .O(gate1089inter12));
  nand2 gate3609(.a(gate1089inter12), .b(gate1089inter1), .O(N5109));
inv1 gate1090( .a(N4617), .O(N5110) );

  xor2  gate3624(.a(N2711), .b(N4617), .O(gate1091inter0));
  nand2 gate3625(.a(gate1091inter0), .b(s_188), .O(gate1091inter1));
  and2  gate3626(.a(N2711), .b(N4617), .O(gate1091inter2));
  inv1  gate3627(.a(s_188), .O(gate1091inter3));
  inv1  gate3628(.a(s_189), .O(gate1091inter4));
  nand2 gate3629(.a(gate1091inter4), .b(gate1091inter3), .O(gate1091inter5));
  nor2  gate3630(.a(gate1091inter5), .b(gate1091inter2), .O(gate1091inter6));
  inv1  gate3631(.a(N4617), .O(gate1091inter7));
  inv1  gate3632(.a(N2711), .O(gate1091inter8));
  nand2 gate3633(.a(gate1091inter8), .b(gate1091inter7), .O(gate1091inter9));
  nand2 gate3634(.a(s_189), .b(gate1091inter3), .O(gate1091inter10));
  nor2  gate3635(.a(gate1091inter10), .b(gate1091inter9), .O(gate1091inter11));
  nor2  gate3636(.a(gate1091inter11), .b(gate1091inter6), .O(gate1091inter12));
  nand2 gate3637(.a(gate1091inter12), .b(gate1091inter1), .O(N5111));
nand2 gate1092( .a(N1890), .b(N4855), .O(N5112) );
inv1 gate1093( .a(N4621), .O(N5113) );
nand2 gate1094( .a(N4621), .b(N2713), .O(N5114) );
inv1 gate1095( .a(N4624), .O(N5115) );

  xor2  gate3176(.a(N2714), .b(N4624), .O(gate1096inter0));
  nand2 gate3177(.a(gate1096inter0), .b(s_124), .O(gate1096inter1));
  and2  gate3178(.a(N2714), .b(N4624), .O(gate1096inter2));
  inv1  gate3179(.a(s_124), .O(gate1096inter3));
  inv1  gate3180(.a(s_125), .O(gate1096inter4));
  nand2 gate3181(.a(gate1096inter4), .b(gate1096inter3), .O(gate1096inter5));
  nor2  gate3182(.a(gate1096inter5), .b(gate1096inter2), .O(gate1096inter6));
  inv1  gate3183(.a(N4624), .O(gate1096inter7));
  inv1  gate3184(.a(N2714), .O(gate1096inter8));
  nand2 gate3185(.a(gate1096inter8), .b(gate1096inter7), .O(gate1096inter9));
  nand2 gate3186(.a(s_125), .b(gate1096inter3), .O(gate1096inter10));
  nor2  gate3187(.a(gate1096inter10), .b(gate1096inter9), .O(gate1096inter11));
  nor2  gate3188(.a(gate1096inter11), .b(gate1096inter6), .O(gate1096inter12));
  nand2 gate3189(.a(gate1096inter12), .b(gate1096inter1), .O(N5116));
and2 gate1097( .a(N4364), .b(N4379), .O(N5117) );
and2 gate1098( .a(N4364), .b(N4379), .O(N5118) );
and2 gate1099( .a(N54), .b(N4405), .O(N5119) );
inv1 gate1100( .a(N4627), .O(N5120) );
nand2 gate1101( .a(N4630), .b(N2716), .O(N5121) );
inv1 gate1102( .a(N4630), .O(N5122) );
nand2 gate1103( .a(N4633), .b(N2717), .O(N5123) );
inv1 gate1104( .a(N4633), .O(N5124) );
nand2 gate1105( .a(N1908), .b(N4909), .O(N5125) );
nand2 gate1106( .a(N4637), .b(N2719), .O(N5126) );
inv1 gate1107( .a(N4637), .O(N5127) );

  xor2  gate3512(.a(N2720), .b(N4640), .O(gate1108inter0));
  nand2 gate3513(.a(gate1108inter0), .b(s_172), .O(gate1108inter1));
  and2  gate3514(.a(N2720), .b(N4640), .O(gate1108inter2));
  inv1  gate3515(.a(s_172), .O(gate1108inter3));
  inv1  gate3516(.a(s_173), .O(gate1108inter4));
  nand2 gate3517(.a(gate1108inter4), .b(gate1108inter3), .O(gate1108inter5));
  nor2  gate3518(.a(gate1108inter5), .b(gate1108inter2), .O(gate1108inter6));
  inv1  gate3519(.a(N4640), .O(gate1108inter7));
  inv1  gate3520(.a(N2720), .O(gate1108inter8));
  nand2 gate3521(.a(gate1108inter8), .b(gate1108inter7), .O(gate1108inter9));
  nand2 gate3522(.a(s_173), .b(gate1108inter3), .O(gate1108inter10));
  nor2  gate3523(.a(gate1108inter10), .b(gate1108inter9), .O(gate1108inter11));
  nor2  gate3524(.a(gate1108inter11), .b(gate1108inter6), .O(gate1108inter12));
  nand2 gate3525(.a(gate1108inter12), .b(gate1108inter1), .O(N5128));
inv1 gate1109( .a(N4640), .O(N5129) );
nand2 gate1110( .a(N4643), .b(N2721), .O(N5130) );
inv1 gate1111( .a(N4643), .O(N5131) );
and2 gate1112( .a(N4425), .b(N4440), .O(N5132) );
and2 gate1113( .a(N4425), .b(N4440), .O(N5133) );
inv1 gate1114( .a(N4649), .O(N5135) );
inv1 gate1115( .a(N4652), .O(N5136) );
nand2 gate1116( .a(N4655), .b(N4521), .O(N5137) );
inv1 gate1117( .a(N4655), .O(N5138) );
inv1 gate1118( .a(N4658), .O(N5139) );

  xor2  gate3470(.a(N4947), .b(N4658), .O(gate1119inter0));
  nand2 gate3471(.a(gate1119inter0), .b(s_166), .O(gate1119inter1));
  and2  gate3472(.a(N4947), .b(N4658), .O(gate1119inter2));
  inv1  gate3473(.a(s_166), .O(gate1119inter3));
  inv1  gate3474(.a(s_167), .O(gate1119inter4));
  nand2 gate3475(.a(gate1119inter4), .b(gate1119inter3), .O(gate1119inter5));
  nor2  gate3476(.a(gate1119inter5), .b(gate1119inter2), .O(gate1119inter6));
  inv1  gate3477(.a(N4658), .O(gate1119inter7));
  inv1  gate3478(.a(N4947), .O(gate1119inter8));
  nand2 gate3479(.a(gate1119inter8), .b(gate1119inter7), .O(gate1119inter9));
  nand2 gate3480(.a(s_167), .b(gate1119inter3), .O(gate1119inter10));
  nor2  gate3481(.a(gate1119inter10), .b(gate1119inter9), .O(gate1119inter11));
  nor2  gate3482(.a(gate1119inter11), .b(gate1119inter6), .O(gate1119inter12));
  nand2 gate3483(.a(gate1119inter12), .b(gate1119inter1), .O(N5140));
inv1 gate1120( .a(N4674), .O(N5141) );
inv1 gate1121( .a(N4677), .O(N5142) );
inv1 gate1122( .a(N4680), .O(N5143) );
inv1 gate1123( .a(N4683), .O(N5144) );
nand2 gate1124( .a(N4686), .b(N4523), .O(N5145) );
inv1 gate1125( .a(N4686), .O(N5146) );
nor2 gate1126( .a(N4953), .b(N4196), .O(N5147) );
nor2 gate1127( .a(N4954), .b(N4955), .O(N5148) );
inv1 gate1128( .a(N4524), .O(N5150) );
nand2 gate1129( .a(N4228), .b(N4965), .O(N5153) );

  xor2  gate2420(.a(N4966), .b(N4225), .O(gate1130inter0));
  nand2 gate2421(.a(gate1130inter0), .b(s_16), .O(gate1130inter1));
  and2  gate2422(.a(N4966), .b(N4225), .O(gate1130inter2));
  inv1  gate2423(.a(s_16), .O(gate1130inter3));
  inv1  gate2424(.a(s_17), .O(gate1130inter4));
  nand2 gate2425(.a(gate1130inter4), .b(gate1130inter3), .O(gate1130inter5));
  nor2  gate2426(.a(gate1130inter5), .b(gate1130inter2), .O(gate1130inter6));
  inv1  gate2427(.a(N4225), .O(gate1130inter7));
  inv1  gate2428(.a(N4966), .O(gate1130inter8));
  nand2 gate2429(.a(gate1130inter8), .b(gate1130inter7), .O(gate1130inter9));
  nand2 gate2430(.a(s_17), .b(gate1130inter3), .O(gate1130inter10));
  nor2  gate2431(.a(gate1130inter10), .b(gate1130inter9), .O(gate1130inter11));
  nor2  gate2432(.a(gate1130inter11), .b(gate1130inter6), .O(gate1130inter12));
  nand2 gate2433(.a(gate1130inter12), .b(gate1130inter1), .O(N5154));
nand2 gate1131( .a(N4234), .b(N4967), .O(N5155) );
nand2 gate1132( .a(N4231), .b(N4968), .O(N5156) );
inv1 gate1133( .a(N4532), .O(N5157) );
nand2 gate1134( .a(N4249), .b(N4972), .O(N5160) );
nand2 gate1135( .a(N4246), .b(N4973), .O(N5161) );
nand2 gate1136( .a(N3816), .b(N4974), .O(N5162) );
and3 gate1137( .a(N4200), .b(N3793), .c(N4976), .O(N5163) );
and3 gate1138( .a(N3789), .b(N4203), .c(N4977), .O(N5164) );
and3 gate1139( .a(N4942), .b(N3147), .c(N3158), .O(N5165) );
inv1 gate1140( .a(N4512), .O(N5166) );
buf1 gate1141( .a(N4290), .O(N5169) );
inv1 gate1142( .a(N4605), .O(N5172) );
buf1 gate1143( .a(N4325), .O(N5173) );
inv1 gate1144( .a(N4608), .O(N5176) );
buf1 gate1145( .a(N4349), .O(N5177) );
buf1 gate1146( .a(N4405), .O(N5180) );
buf1 gate1147( .a(N4357), .O(N5183) );
buf1 gate1148( .a(N4357), .O(N5186) );
buf1 gate1149( .a(N4364), .O(N5189) );
buf1 gate1150( .a(N4364), .O(N5192) );
buf1 gate1151( .a(N4385), .O(N5195) );
inv1 gate1152( .a(N4646), .O(N5198) );
buf1 gate1153( .a(N4418), .O(N5199) );
buf1 gate1154( .a(N4425), .O(N5202) );
buf1 gate1155( .a(N4445), .O(N5205) );
buf1 gate1156( .a(N4418), .O(N5208) );
buf1 gate1157( .a(N4425), .O(N5211) );
buf1 gate1158( .a(N4477), .O(N5214) );
buf1 gate1159( .a(N4469), .O(N5217) );
buf1 gate1160( .a(N4477), .O(N5220) );
inv1 gate1161( .a(N4662), .O(N5223) );
inv1 gate1162( .a(N4665), .O(N5224) );
inv1 gate1163( .a(N4668), .O(N5225) );
inv1 gate1164( .a(N4671), .O(N5226) );
inv1 gate1165( .a(N4689), .O(N5227) );
inv1 gate1166( .a(N4692), .O(N5228) );
inv1 gate1167( .a(N4695), .O(N5229) );
inv1 gate1168( .a(N4698), .O(N5230) );
nand2 gate1169( .a(N4240), .b(N5052), .O(N5232) );
nand2 gate1170( .a(N4237), .b(N5053), .O(N5233) );
nand2 gate1171( .a(N4258), .b(N5055), .O(N5234) );
nand2 gate1172( .a(N4255), .b(N5056), .O(N5235) );

  xor2  gate3862(.a(N5057), .b(N4721), .O(gate1173inter0));
  nand2 gate3863(.a(gate1173inter0), .b(s_222), .O(gate1173inter1));
  and2  gate3864(.a(N5057), .b(N4721), .O(gate1173inter2));
  inv1  gate3865(.a(s_222), .O(gate1173inter3));
  inv1  gate3866(.a(s_223), .O(gate1173inter4));
  nand2 gate3867(.a(gate1173inter4), .b(gate1173inter3), .O(gate1173inter5));
  nor2  gate3868(.a(gate1173inter5), .b(gate1173inter2), .O(gate1173inter6));
  inv1  gate3869(.a(N4721), .O(gate1173inter7));
  inv1  gate3870(.a(N5057), .O(gate1173inter8));
  nand2 gate3871(.a(gate1173inter8), .b(gate1173inter7), .O(gate1173inter9));
  nand2 gate3872(.a(s_223), .b(gate1173inter3), .O(gate1173inter10));
  nor2  gate3873(.a(gate1173inter10), .b(gate1173inter9), .O(gate1173inter11));
  nor2  gate3874(.a(gate1173inter11), .b(gate1173inter6), .O(gate1173inter12));
  nand2 gate3875(.a(gate1173inter12), .b(gate1173inter1), .O(N5236));
nand2 gate1174( .a(N3824), .b(N5058), .O(N5239) );
and3 gate1175( .a(N5060), .b(N5061), .c(N4270), .O(N5240) );
inv1 gate1176( .a(N4939), .O(N5241) );
nand2 gate1177( .a(N1824), .b(N5069), .O(N5242) );
nand2 gate1178( .a(N1827), .b(N5071), .O(N5243) );

  xor2  gate2560(.a(N5073), .b(N1830), .O(gate1179inter0));
  nand2 gate2561(.a(gate1179inter0), .b(s_36), .O(gate1179inter1));
  and2  gate2562(.a(N5073), .b(N1830), .O(gate1179inter2));
  inv1  gate2563(.a(s_36), .O(gate1179inter3));
  inv1  gate2564(.a(s_37), .O(gate1179inter4));
  nand2 gate2565(.a(gate1179inter4), .b(gate1179inter3), .O(gate1179inter5));
  nor2  gate2566(.a(gate1179inter5), .b(gate1179inter2), .O(gate1179inter6));
  inv1  gate2567(.a(N1830), .O(gate1179inter7));
  inv1  gate2568(.a(N5073), .O(gate1179inter8));
  nand2 gate2569(.a(gate1179inter8), .b(gate1179inter7), .O(gate1179inter9));
  nand2 gate2570(.a(s_37), .b(gate1179inter3), .O(gate1179inter10));
  nor2  gate2571(.a(gate1179inter10), .b(gate1179inter9), .O(gate1179inter11));
  nor2  gate2572(.a(gate1179inter11), .b(gate1179inter6), .O(gate1179inter12));
  nand2 gate2573(.a(gate1179inter12), .b(gate1179inter1), .O(N5244));
nand2 gate1180( .a(N1833), .b(N5075), .O(N5245) );
nand2 gate1181( .a(N1836), .b(N5077), .O(N5246) );

  xor2  gate3974(.a(N5079), .b(N1839), .O(gate1182inter0));
  nand2 gate3975(.a(gate1182inter0), .b(s_238), .O(gate1182inter1));
  and2  gate3976(.a(N5079), .b(N1839), .O(gate1182inter2));
  inv1  gate3977(.a(s_238), .O(gate1182inter3));
  inv1  gate3978(.a(s_239), .O(gate1182inter4));
  nand2 gate3979(.a(gate1182inter4), .b(gate1182inter3), .O(gate1182inter5));
  nor2  gate3980(.a(gate1182inter5), .b(gate1182inter2), .O(gate1182inter6));
  inv1  gate3981(.a(N1839), .O(gate1182inter7));
  inv1  gate3982(.a(N5079), .O(gate1182inter8));
  nand2 gate3983(.a(gate1182inter8), .b(gate1182inter7), .O(gate1182inter9));
  nand2 gate3984(.a(s_239), .b(gate1182inter3), .O(gate1182inter10));
  nor2  gate3985(.a(gate1182inter10), .b(gate1182inter9), .O(gate1182inter11));
  nor2  gate3986(.a(gate1182inter11), .b(gate1182inter6), .O(gate1182inter12));
  nand2 gate3987(.a(gate1182inter12), .b(gate1182inter1), .O(N5247));
nand2 gate1183( .a(N1842), .b(N5081), .O(N5248) );
nand2 gate1184( .a(N1845), .b(N5083), .O(N5249) );
nand2 gate1185( .a(N1848), .b(N5085), .O(N5250) );

  xor2  gate3960(.a(N5089), .b(N1854), .O(gate1186inter0));
  nand2 gate3961(.a(gate1186inter0), .b(s_236), .O(gate1186inter1));
  and2  gate3962(.a(N5089), .b(N1854), .O(gate1186inter2));
  inv1  gate3963(.a(s_236), .O(gate1186inter3));
  inv1  gate3964(.a(s_237), .O(gate1186inter4));
  nand2 gate3965(.a(gate1186inter4), .b(gate1186inter3), .O(gate1186inter5));
  nor2  gate3966(.a(gate1186inter5), .b(gate1186inter2), .O(gate1186inter6));
  inv1  gate3967(.a(N1854), .O(gate1186inter7));
  inv1  gate3968(.a(N5089), .O(gate1186inter8));
  nand2 gate3969(.a(gate1186inter8), .b(gate1186inter7), .O(gate1186inter9));
  nand2 gate3970(.a(s_237), .b(gate1186inter3), .O(gate1186inter10));
  nor2  gate3971(.a(gate1186inter10), .b(gate1186inter9), .O(gate1186inter11));
  nor2  gate3972(.a(gate1186inter11), .b(gate1186inter6), .O(gate1186inter12));
  nand2 gate3973(.a(gate1186inter12), .b(gate1186inter1), .O(N5252));
nand2 gate1187( .a(N1857), .b(N5091), .O(N5253) );
nand2 gate1188( .a(N1860), .b(N5093), .O(N5254) );

  xor2  gate3442(.a(N5095), .b(N1863), .O(gate1189inter0));
  nand2 gate3443(.a(gate1189inter0), .b(s_162), .O(gate1189inter1));
  and2  gate3444(.a(N5095), .b(N1863), .O(gate1189inter2));
  inv1  gate3445(.a(s_162), .O(gate1189inter3));
  inv1  gate3446(.a(s_163), .O(gate1189inter4));
  nand2 gate3447(.a(gate1189inter4), .b(gate1189inter3), .O(gate1189inter5));
  nor2  gate3448(.a(gate1189inter5), .b(gate1189inter2), .O(gate1189inter6));
  inv1  gate3449(.a(N1863), .O(gate1189inter7));
  inv1  gate3450(.a(N5095), .O(gate1189inter8));
  nand2 gate3451(.a(gate1189inter8), .b(gate1189inter7), .O(gate1189inter9));
  nand2 gate3452(.a(s_163), .b(gate1189inter3), .O(gate1189inter10));
  nor2  gate3453(.a(gate1189inter10), .b(gate1189inter9), .O(gate1189inter11));
  nor2  gate3454(.a(gate1189inter11), .b(gate1189inter6), .O(gate1189inter12));
  nand2 gate3455(.a(gate1189inter12), .b(gate1189inter1), .O(N5255));
nand2 gate1190( .a(N1866), .b(N5097), .O(N5256) );
nand2 gate1191( .a(N1869), .b(N5099), .O(N5257) );
nand2 gate1192( .a(N1872), .b(N5101), .O(N5258) );
nand2 gate1193( .a(N1875), .b(N5103), .O(N5259) );
nand2 gate1194( .a(N1878), .b(N5105), .O(N5260) );
nand2 gate1195( .a(N1881), .b(N5106), .O(N5261) );
nand2 gate1196( .a(N1884), .b(N5108), .O(N5262) );

  xor2  gate3022(.a(N5110), .b(N1887), .O(gate1197inter0));
  nand2 gate3023(.a(gate1197inter0), .b(s_102), .O(gate1197inter1));
  and2  gate3024(.a(N5110), .b(N1887), .O(gate1197inter2));
  inv1  gate3025(.a(s_102), .O(gate1197inter3));
  inv1  gate3026(.a(s_103), .O(gate1197inter4));
  nand2 gate3027(.a(gate1197inter4), .b(gate1197inter3), .O(gate1197inter5));
  nor2  gate3028(.a(gate1197inter5), .b(gate1197inter2), .O(gate1197inter6));
  inv1  gate3029(.a(N1887), .O(gate1197inter7));
  inv1  gate3030(.a(N5110), .O(gate1197inter8));
  nand2 gate3031(.a(gate1197inter8), .b(gate1197inter7), .O(gate1197inter9));
  nand2 gate3032(.a(s_103), .b(gate1197inter3), .O(gate1197inter10));
  nor2  gate3033(.a(gate1197inter10), .b(gate1197inter9), .O(gate1197inter11));
  nor2  gate3034(.a(gate1197inter11), .b(gate1197inter6), .O(gate1197inter12));
  nand2 gate3035(.a(gate1197inter12), .b(gate1197inter1), .O(N5263));
nand2 gate1198( .a(N5112), .b(N4856), .O(N5264) );
nand2 gate1199( .a(N1893), .b(N5113), .O(N5274) );
nand2 gate1200( .a(N1896), .b(N5115), .O(N5275) );
nand2 gate1201( .a(N1902), .b(N5122), .O(N5282) );
nand2 gate1202( .a(N1905), .b(N5124), .O(N5283) );
nand2 gate1203( .a(N4908), .b(N5125), .O(N5284) );
nand2 gate1204( .a(N1911), .b(N5127), .O(N5298) );
nand2 gate1205( .a(N1914), .b(N5129), .O(N5299) );
nand2 gate1206( .a(N1917), .b(N5131), .O(N5300) );
nand2 gate1207( .a(N4652), .b(N5135), .O(N5303) );
nand2 gate1208( .a(N4649), .b(N5136), .O(N5304) );
nand2 gate1209( .a(N4008), .b(N5138), .O(N5305) );
nand2 gate1210( .a(N4219), .b(N5139), .O(N5306) );
nand2 gate1211( .a(N4677), .b(N5141), .O(N5307) );
nand2 gate1212( .a(N4674), .b(N5142), .O(N5308) );

  xor2  gate2616(.a(N5143), .b(N4683), .O(gate1213inter0));
  nand2 gate2617(.a(gate1213inter0), .b(s_44), .O(gate1213inter1));
  and2  gate2618(.a(N5143), .b(N4683), .O(gate1213inter2));
  inv1  gate2619(.a(s_44), .O(gate1213inter3));
  inv1  gate2620(.a(s_45), .O(gate1213inter4));
  nand2 gate2621(.a(gate1213inter4), .b(gate1213inter3), .O(gate1213inter5));
  nor2  gate2622(.a(gate1213inter5), .b(gate1213inter2), .O(gate1213inter6));
  inv1  gate2623(.a(N4683), .O(gate1213inter7));
  inv1  gate2624(.a(N5143), .O(gate1213inter8));
  nand2 gate2625(.a(gate1213inter8), .b(gate1213inter7), .O(gate1213inter9));
  nand2 gate2626(.a(s_45), .b(gate1213inter3), .O(gate1213inter10));
  nor2  gate2627(.a(gate1213inter10), .b(gate1213inter9), .O(gate1213inter11));
  nor2  gate2628(.a(gate1213inter11), .b(gate1213inter6), .O(gate1213inter12));
  nand2 gate2629(.a(gate1213inter12), .b(gate1213inter1), .O(N5309));
nand2 gate1214( .a(N4680), .b(N5144), .O(N5310) );
nand2 gate1215( .a(N4011), .b(N5146), .O(N5311) );
inv1 gate1216( .a(N5049), .O(N5312) );
nand2 gate1217( .a(N5153), .b(N5154), .O(N5315) );
nand2 gate1218( .a(N5155), .b(N5156), .O(N5319) );

  xor2  gate2476(.a(N5161), .b(N5160), .O(gate1219inter0));
  nand2 gate2477(.a(gate1219inter0), .b(s_24), .O(gate1219inter1));
  and2  gate2478(.a(N5161), .b(N5160), .O(gate1219inter2));
  inv1  gate2479(.a(s_24), .O(gate1219inter3));
  inv1  gate2480(.a(s_25), .O(gate1219inter4));
  nand2 gate2481(.a(gate1219inter4), .b(gate1219inter3), .O(gate1219inter5));
  nor2  gate2482(.a(gate1219inter5), .b(gate1219inter2), .O(gate1219inter6));
  inv1  gate2483(.a(N5160), .O(gate1219inter7));
  inv1  gate2484(.a(N5161), .O(gate1219inter8));
  nand2 gate2485(.a(gate1219inter8), .b(gate1219inter7), .O(gate1219inter9));
  nand2 gate2486(.a(s_25), .b(gate1219inter3), .O(gate1219inter10));
  nor2  gate2487(.a(gate1219inter10), .b(gate1219inter9), .O(gate1219inter11));
  nor2  gate2488(.a(gate1219inter11), .b(gate1219inter6), .O(gate1219inter12));
  nand2 gate2489(.a(gate1219inter12), .b(gate1219inter1), .O(N5324));
nand2 gate1220( .a(N5162), .b(N4975), .O(N5328) );
nor2 gate1221( .a(N5163), .b(N4978), .O(N5331) );
nor2 gate1222( .a(N5164), .b(N4979), .O(N5332) );
or2 gate1223( .a(N4412), .b(N5119), .O(N5346) );
nand2 gate1224( .a(N4665), .b(N5223), .O(N5363) );
nand2 gate1225( .a(N4662), .b(N5224), .O(N5364) );

  xor2  gate3918(.a(N5225), .b(N4671), .O(gate1226inter0));
  nand2 gate3919(.a(gate1226inter0), .b(s_230), .O(gate1226inter1));
  and2  gate3920(.a(N5225), .b(N4671), .O(gate1226inter2));
  inv1  gate3921(.a(s_230), .O(gate1226inter3));
  inv1  gate3922(.a(s_231), .O(gate1226inter4));
  nand2 gate3923(.a(gate1226inter4), .b(gate1226inter3), .O(gate1226inter5));
  nor2  gate3924(.a(gate1226inter5), .b(gate1226inter2), .O(gate1226inter6));
  inv1  gate3925(.a(N4671), .O(gate1226inter7));
  inv1  gate3926(.a(N5225), .O(gate1226inter8));
  nand2 gate3927(.a(gate1226inter8), .b(gate1226inter7), .O(gate1226inter9));
  nand2 gate3928(.a(s_231), .b(gate1226inter3), .O(gate1226inter10));
  nor2  gate3929(.a(gate1226inter10), .b(gate1226inter9), .O(gate1226inter11));
  nor2  gate3930(.a(gate1226inter11), .b(gate1226inter6), .O(gate1226inter12));
  nand2 gate3931(.a(gate1226inter12), .b(gate1226inter1), .O(N5365));
nand2 gate1227( .a(N4668), .b(N5226), .O(N5366) );

  xor2  gate2910(.a(N5227), .b(N4692), .O(gate1228inter0));
  nand2 gate2911(.a(gate1228inter0), .b(s_86), .O(gate1228inter1));
  and2  gate2912(.a(N5227), .b(N4692), .O(gate1228inter2));
  inv1  gate2913(.a(s_86), .O(gate1228inter3));
  inv1  gate2914(.a(s_87), .O(gate1228inter4));
  nand2 gate2915(.a(gate1228inter4), .b(gate1228inter3), .O(gate1228inter5));
  nor2  gate2916(.a(gate1228inter5), .b(gate1228inter2), .O(gate1228inter6));
  inv1  gate2917(.a(N4692), .O(gate1228inter7));
  inv1  gate2918(.a(N5227), .O(gate1228inter8));
  nand2 gate2919(.a(gate1228inter8), .b(gate1228inter7), .O(gate1228inter9));
  nand2 gate2920(.a(s_87), .b(gate1228inter3), .O(gate1228inter10));
  nor2  gate2921(.a(gate1228inter10), .b(gate1228inter9), .O(gate1228inter11));
  nor2  gate2922(.a(gate1228inter11), .b(gate1228inter6), .O(gate1228inter12));
  nand2 gate2923(.a(gate1228inter12), .b(gate1228inter1), .O(N5367));
nand2 gate1229( .a(N4689), .b(N5228), .O(N5368) );
nand2 gate1230( .a(N4698), .b(N5229), .O(N5369) );
nand2 gate1231( .a(N4695), .b(N5230), .O(N5370) );

  xor2  gate2728(.a(N5147), .b(N5148), .O(gate1232inter0));
  nand2 gate2729(.a(gate1232inter0), .b(s_60), .O(gate1232inter1));
  and2  gate2730(.a(N5147), .b(N5148), .O(gate1232inter2));
  inv1  gate2731(.a(s_60), .O(gate1232inter3));
  inv1  gate2732(.a(s_61), .O(gate1232inter4));
  nand2 gate2733(.a(gate1232inter4), .b(gate1232inter3), .O(gate1232inter5));
  nor2  gate2734(.a(gate1232inter5), .b(gate1232inter2), .O(gate1232inter6));
  inv1  gate2735(.a(N5148), .O(gate1232inter7));
  inv1  gate2736(.a(N5147), .O(gate1232inter8));
  nand2 gate2737(.a(gate1232inter8), .b(gate1232inter7), .O(gate1232inter9));
  nand2 gate2738(.a(s_61), .b(gate1232inter3), .O(gate1232inter10));
  nor2  gate2739(.a(gate1232inter10), .b(gate1232inter9), .O(gate1232inter11));
  nor2  gate2740(.a(gate1232inter11), .b(gate1232inter6), .O(gate1232inter12));
  nand2 gate2741(.a(gate1232inter12), .b(gate1232inter1), .O(N5371));
buf1 gate1233( .a(N4939), .O(N5374) );
nand2 gate1234( .a(N5232), .b(N5233), .O(N5377) );
nand2 gate1235( .a(N5234), .b(N5235), .O(N5382) );
nand2 gate1236( .a(N5239), .b(N5059), .O(N5385) );
and3 gate1237( .a(N5062), .b(N5063), .c(N5241), .O(N5388) );
nand2 gate1238( .a(N5242), .b(N5070), .O(N5389) );
nand2 gate1239( .a(N5243), .b(N5072), .O(N5396) );
nand2 gate1240( .a(N5244), .b(N5074), .O(N5407) );
nand2 gate1241( .a(N5245), .b(N5076), .O(N5418) );
nand2 gate1242( .a(N5246), .b(N5078), .O(N5424) );
nand2 gate1243( .a(N5247), .b(N5080), .O(N5431) );

  xor2  gate3064(.a(N5082), .b(N5248), .O(gate1244inter0));
  nand2 gate3065(.a(gate1244inter0), .b(s_108), .O(gate1244inter1));
  and2  gate3066(.a(N5082), .b(N5248), .O(gate1244inter2));
  inv1  gate3067(.a(s_108), .O(gate1244inter3));
  inv1  gate3068(.a(s_109), .O(gate1244inter4));
  nand2 gate3069(.a(gate1244inter4), .b(gate1244inter3), .O(gate1244inter5));
  nor2  gate3070(.a(gate1244inter5), .b(gate1244inter2), .O(gate1244inter6));
  inv1  gate3071(.a(N5248), .O(gate1244inter7));
  inv1  gate3072(.a(N5082), .O(gate1244inter8));
  nand2 gate3073(.a(gate1244inter8), .b(gate1244inter7), .O(gate1244inter9));
  nand2 gate3074(.a(s_109), .b(gate1244inter3), .O(gate1244inter10));
  nor2  gate3075(.a(gate1244inter10), .b(gate1244inter9), .O(gate1244inter11));
  nor2  gate3076(.a(gate1244inter11), .b(gate1244inter6), .O(gate1244inter12));
  nand2 gate3077(.a(gate1244inter12), .b(gate1244inter1), .O(N5441));
nand2 gate1245( .a(N5249), .b(N5084), .O(N5452) );
nand2 gate1246( .a(N5250), .b(N5086), .O(N5462) );
inv1 gate1247( .a(N5169), .O(N5469) );
nand2 gate1248( .a(N5088), .b(N5252), .O(N5470) );
nand2 gate1249( .a(N5090), .b(N5253), .O(N5477) );
nand2 gate1250( .a(N5092), .b(N5254), .O(N5488) );
nand2 gate1251( .a(N5094), .b(N5255), .O(N5498) );

  xor2  gate2798(.a(N5256), .b(N5096), .O(gate1252inter0));
  nand2 gate2799(.a(gate1252inter0), .b(s_70), .O(gate1252inter1));
  and2  gate2800(.a(N5256), .b(N5096), .O(gate1252inter2));
  inv1  gate2801(.a(s_70), .O(gate1252inter3));
  inv1  gate2802(.a(s_71), .O(gate1252inter4));
  nand2 gate2803(.a(gate1252inter4), .b(gate1252inter3), .O(gate1252inter5));
  nor2  gate2804(.a(gate1252inter5), .b(gate1252inter2), .O(gate1252inter6));
  inv1  gate2805(.a(N5096), .O(gate1252inter7));
  inv1  gate2806(.a(N5256), .O(gate1252inter8));
  nand2 gate2807(.a(gate1252inter8), .b(gate1252inter7), .O(gate1252inter9));
  nand2 gate2808(.a(s_71), .b(gate1252inter3), .O(gate1252inter10));
  nor2  gate2809(.a(gate1252inter10), .b(gate1252inter9), .O(gate1252inter11));
  nor2  gate2810(.a(gate1252inter11), .b(gate1252inter6), .O(gate1252inter12));
  nand2 gate2811(.a(gate1252inter12), .b(gate1252inter1), .O(N5506));
nand2 gate1253( .a(N5098), .b(N5257), .O(N5520) );
nand2 gate1254( .a(N5100), .b(N5258), .O(N5536) );

  xor2  gate3162(.a(N5259), .b(N5102), .O(gate1255inter0));
  nand2 gate3163(.a(gate1255inter0), .b(s_122), .O(gate1255inter1));
  and2  gate3164(.a(N5259), .b(N5102), .O(gate1255inter2));
  inv1  gate3165(.a(s_122), .O(gate1255inter3));
  inv1  gate3166(.a(s_123), .O(gate1255inter4));
  nand2 gate3167(.a(gate1255inter4), .b(gate1255inter3), .O(gate1255inter5));
  nor2  gate3168(.a(gate1255inter5), .b(gate1255inter2), .O(gate1255inter6));
  inv1  gate3169(.a(N5102), .O(gate1255inter7));
  inv1  gate3170(.a(N5259), .O(gate1255inter8));
  nand2 gate3171(.a(gate1255inter8), .b(gate1255inter7), .O(gate1255inter9));
  nand2 gate3172(.a(s_123), .b(gate1255inter3), .O(gate1255inter10));
  nor2  gate3173(.a(gate1255inter10), .b(gate1255inter9), .O(gate1255inter11));
  nor2  gate3174(.a(gate1255inter11), .b(gate1255inter6), .O(gate1255inter12));
  nand2 gate3175(.a(gate1255inter12), .b(gate1255inter1), .O(N5549));
nand2 gate1256( .a(N5104), .b(N5260), .O(N5555) );
nand2 gate1257( .a(N5261), .b(N5107), .O(N5562) );
nand2 gate1258( .a(N5262), .b(N5109), .O(N5573) );
nand2 gate1259( .a(N5263), .b(N5111), .O(N5579) );
nand2 gate1260( .a(N5274), .b(N5114), .O(N5595) );
nand2 gate1261( .a(N5275), .b(N5116), .O(N5606) );
nand2 gate1262( .a(N5180), .b(N2715), .O(N5616) );
inv1 gate1263( .a(N5180), .O(N5617) );
inv1 gate1264( .a(N5183), .O(N5618) );
inv1 gate1265( .a(N5186), .O(N5619) );
inv1 gate1266( .a(N5189), .O(N5620) );
inv1 gate1267( .a(N5192), .O(N5621) );
inv1 gate1268( .a(N5195), .O(N5622) );

  xor2  gate3582(.a(N5282), .b(N5121), .O(gate1269inter0));
  nand2 gate3583(.a(gate1269inter0), .b(s_182), .O(gate1269inter1));
  and2  gate3584(.a(N5282), .b(N5121), .O(gate1269inter2));
  inv1  gate3585(.a(s_182), .O(gate1269inter3));
  inv1  gate3586(.a(s_183), .O(gate1269inter4));
  nand2 gate3587(.a(gate1269inter4), .b(gate1269inter3), .O(gate1269inter5));
  nor2  gate3588(.a(gate1269inter5), .b(gate1269inter2), .O(gate1269inter6));
  inv1  gate3589(.a(N5121), .O(gate1269inter7));
  inv1  gate3590(.a(N5282), .O(gate1269inter8));
  nand2 gate3591(.a(gate1269inter8), .b(gate1269inter7), .O(gate1269inter9));
  nand2 gate3592(.a(s_183), .b(gate1269inter3), .O(gate1269inter10));
  nor2  gate3593(.a(gate1269inter10), .b(gate1269inter9), .O(gate1269inter11));
  nor2  gate3594(.a(gate1269inter11), .b(gate1269inter6), .O(gate1269inter12));
  nand2 gate3595(.a(gate1269inter12), .b(gate1269inter1), .O(N5624));
nand2 gate1270( .a(N5123), .b(N5283), .O(N5634) );
nand2 gate1271( .a(N5126), .b(N5298), .O(N5655) );
nand2 gate1272( .a(N5128), .b(N5299), .O(N5671) );
nand2 gate1273( .a(N5130), .b(N5300), .O(N5684) );
inv1 gate1274( .a(N5202), .O(N5690) );
inv1 gate1275( .a(N5211), .O(N5691) );
nand2 gate1276( .a(N5303), .b(N5304), .O(N5692) );
nand2 gate1277( .a(N5137), .b(N5305), .O(N5696) );
nand2 gate1278( .a(N5306), .b(N5140), .O(N5700) );
nand2 gate1279( .a(N5307), .b(N5308), .O(N5703) );

  xor2  gate3946(.a(N5310), .b(N5309), .O(gate1280inter0));
  nand2 gate3947(.a(gate1280inter0), .b(s_234), .O(gate1280inter1));
  and2  gate3948(.a(N5310), .b(N5309), .O(gate1280inter2));
  inv1  gate3949(.a(s_234), .O(gate1280inter3));
  inv1  gate3950(.a(s_235), .O(gate1280inter4));
  nand2 gate3951(.a(gate1280inter4), .b(gate1280inter3), .O(gate1280inter5));
  nor2  gate3952(.a(gate1280inter5), .b(gate1280inter2), .O(gate1280inter6));
  inv1  gate3953(.a(N5309), .O(gate1280inter7));
  inv1  gate3954(.a(N5310), .O(gate1280inter8));
  nand2 gate3955(.a(gate1280inter8), .b(gate1280inter7), .O(gate1280inter9));
  nand2 gate3956(.a(s_235), .b(gate1280inter3), .O(gate1280inter10));
  nor2  gate3957(.a(gate1280inter10), .b(gate1280inter9), .O(gate1280inter11));
  nor2  gate3958(.a(gate1280inter11), .b(gate1280inter6), .O(gate1280inter12));
  nand2 gate3959(.a(gate1280inter12), .b(gate1280inter1), .O(N5707));
nand2 gate1281( .a(N5145), .b(N5311), .O(N5711) );
and2 gate1282( .a(N5166), .b(N4512), .O(N5726) );
inv1 gate1283( .a(N5173), .O(N5727) );
inv1 gate1284( .a(N5177), .O(N5728) );
inv1 gate1285( .a(N5199), .O(N5730) );
inv1 gate1286( .a(N5205), .O(N5731) );
inv1 gate1287( .a(N5208), .O(N5732) );
inv1 gate1288( .a(N5214), .O(N5733) );
inv1 gate1289( .a(N5217), .O(N5734) );
inv1 gate1290( .a(N5220), .O(N5735) );
nand2 gate1291( .a(N5365), .b(N5366), .O(N5736) );

  xor2  gate2980(.a(N5364), .b(N5363), .O(gate1292inter0));
  nand2 gate2981(.a(gate1292inter0), .b(s_96), .O(gate1292inter1));
  and2  gate2982(.a(N5364), .b(N5363), .O(gate1292inter2));
  inv1  gate2983(.a(s_96), .O(gate1292inter3));
  inv1  gate2984(.a(s_97), .O(gate1292inter4));
  nand2 gate2985(.a(gate1292inter4), .b(gate1292inter3), .O(gate1292inter5));
  nor2  gate2986(.a(gate1292inter5), .b(gate1292inter2), .O(gate1292inter6));
  inv1  gate2987(.a(N5363), .O(gate1292inter7));
  inv1  gate2988(.a(N5364), .O(gate1292inter8));
  nand2 gate2989(.a(gate1292inter8), .b(gate1292inter7), .O(gate1292inter9));
  nand2 gate2990(.a(s_97), .b(gate1292inter3), .O(gate1292inter10));
  nor2  gate2991(.a(gate1292inter10), .b(gate1292inter9), .O(gate1292inter11));
  nor2  gate2992(.a(gate1292inter11), .b(gate1292inter6), .O(gate1292inter12));
  nand2 gate2993(.a(gate1292inter12), .b(gate1292inter1), .O(N5739));

  xor2  gate3932(.a(N5370), .b(N5369), .O(gate1293inter0));
  nand2 gate3933(.a(gate1293inter0), .b(s_232), .O(gate1293inter1));
  and2  gate3934(.a(N5370), .b(N5369), .O(gate1293inter2));
  inv1  gate3935(.a(s_232), .O(gate1293inter3));
  inv1  gate3936(.a(s_233), .O(gate1293inter4));
  nand2 gate3937(.a(gate1293inter4), .b(gate1293inter3), .O(gate1293inter5));
  nor2  gate3938(.a(gate1293inter5), .b(gate1293inter2), .O(gate1293inter6));
  inv1  gate3939(.a(N5369), .O(gate1293inter7));
  inv1  gate3940(.a(N5370), .O(gate1293inter8));
  nand2 gate3941(.a(gate1293inter8), .b(gate1293inter7), .O(gate1293inter9));
  nand2 gate3942(.a(s_233), .b(gate1293inter3), .O(gate1293inter10));
  nor2  gate3943(.a(gate1293inter10), .b(gate1293inter9), .O(gate1293inter11));
  nor2  gate3944(.a(gate1293inter11), .b(gate1293inter6), .O(gate1293inter12));
  nand2 gate3945(.a(gate1293inter12), .b(gate1293inter1), .O(N5742));

  xor2  gate3260(.a(N5368), .b(N5367), .O(gate1294inter0));
  nand2 gate3261(.a(gate1294inter0), .b(s_136), .O(gate1294inter1));
  and2  gate3262(.a(N5368), .b(N5367), .O(gate1294inter2));
  inv1  gate3263(.a(s_136), .O(gate1294inter3));
  inv1  gate3264(.a(s_137), .O(gate1294inter4));
  nand2 gate3265(.a(gate1294inter4), .b(gate1294inter3), .O(gate1294inter5));
  nor2  gate3266(.a(gate1294inter5), .b(gate1294inter2), .O(gate1294inter6));
  inv1  gate3267(.a(N5367), .O(gate1294inter7));
  inv1  gate3268(.a(N5368), .O(gate1294inter8));
  nand2 gate3269(.a(gate1294inter8), .b(gate1294inter7), .O(gate1294inter9));
  nand2 gate3270(.a(s_137), .b(gate1294inter3), .O(gate1294inter10));
  nor2  gate3271(.a(gate1294inter10), .b(gate1294inter9), .O(gate1294inter11));
  nor2  gate3272(.a(gate1294inter11), .b(gate1294inter6), .O(gate1294inter12));
  nand2 gate3273(.a(gate1294inter12), .b(gate1294inter1), .O(N5745));
inv1 gate1295( .a(N5236), .O(N5755) );

  xor2  gate2518(.a(N5331), .b(N5332), .O(gate1296inter0));
  nand2 gate2519(.a(gate1296inter0), .b(s_30), .O(gate1296inter1));
  and2  gate2520(.a(N5331), .b(N5332), .O(gate1296inter2));
  inv1  gate2521(.a(s_30), .O(gate1296inter3));
  inv1  gate2522(.a(s_31), .O(gate1296inter4));
  nand2 gate2523(.a(gate1296inter4), .b(gate1296inter3), .O(gate1296inter5));
  nor2  gate2524(.a(gate1296inter5), .b(gate1296inter2), .O(gate1296inter6));
  inv1  gate2525(.a(N5332), .O(gate1296inter7));
  inv1  gate2526(.a(N5331), .O(gate1296inter8));
  nand2 gate2527(.a(gate1296inter8), .b(gate1296inter7), .O(gate1296inter9));
  nand2 gate2528(.a(s_31), .b(gate1296inter3), .O(gate1296inter10));
  nor2  gate2529(.a(gate1296inter10), .b(gate1296inter9), .O(gate1296inter11));
  nor2  gate2530(.a(gate1296inter11), .b(gate1296inter6), .O(gate1296inter12));
  nand2 gate2531(.a(gate1296inter12), .b(gate1296inter1), .O(N5756));
and2 gate1297( .a(N5264), .b(N4396), .O(N5954) );
nand2 gate1298( .a(N1899), .b(N5617), .O(N5955) );
inv1 gate1299( .a(N5346), .O(N5956) );
and2 gate1300( .a(N5284), .b(N4456), .O(N6005) );
and2 gate1301( .a(N5284), .b(N4456), .O(N6006) );
inv1 gate1302( .a(N5371), .O(N6023) );
nand2 gate1303( .a(N5371), .b(N5312), .O(N6024) );
inv1 gate1304( .a(N5315), .O(N6025) );
inv1 gate1305( .a(N5324), .O(N6028) );
buf1 gate1306( .a(N5319), .O(N6031) );
buf1 gate1307( .a(N5319), .O(N6034) );
buf1 gate1308( .a(N5328), .O(N6037) );
buf1 gate1309( .a(N5328), .O(N6040) );
inv1 gate1310( .a(N5385), .O(N6044) );
or2 gate1311( .a(N5166), .b(N5726), .O(N6045) );
buf1 gate1312( .a(N5264), .O(N6048) );
buf1 gate1313( .a(N5284), .O(N6051) );
buf1 gate1314( .a(N5284), .O(N6054) );
inv1 gate1315( .a(N5374), .O(N6065) );
nand2 gate1316( .a(N5374), .b(N5054), .O(N6066) );
inv1 gate1317( .a(N5377), .O(N6067) );
inv1 gate1318( .a(N5382), .O(N6068) );

  xor2  gate2658(.a(N5755), .b(N5382), .O(gate1319inter0));
  nand2 gate2659(.a(gate1319inter0), .b(s_50), .O(gate1319inter1));
  and2  gate2660(.a(N5755), .b(N5382), .O(gate1319inter2));
  inv1  gate2661(.a(s_50), .O(gate1319inter3));
  inv1  gate2662(.a(s_51), .O(gate1319inter4));
  nand2 gate2663(.a(gate1319inter4), .b(gate1319inter3), .O(gate1319inter5));
  nor2  gate2664(.a(gate1319inter5), .b(gate1319inter2), .O(gate1319inter6));
  inv1  gate2665(.a(N5382), .O(gate1319inter7));
  inv1  gate2666(.a(N5755), .O(gate1319inter8));
  nand2 gate2667(.a(gate1319inter8), .b(gate1319inter7), .O(gate1319inter9));
  nand2 gate2668(.a(s_51), .b(gate1319inter3), .O(gate1319inter10));
  nor2  gate2669(.a(gate1319inter10), .b(gate1319inter9), .O(gate1319inter11));
  nor2  gate2670(.a(gate1319inter11), .b(gate1319inter6), .O(gate1319inter12));
  nand2 gate2671(.a(gate1319inter12), .b(gate1319inter1), .O(N6069));
and2 gate1320( .a(N5470), .b(N4316), .O(N6071) );
and3 gate1321( .a(N5477), .b(N5470), .c(N4320), .O(N6072) );
and4 gate1322( .a(N5488), .b(N5470), .c(N4325), .d(N5477), .O(N6073) );
and4 gate1323( .a(N5562), .b(N4357), .c(N4385), .d(N4364), .O(N6074) );
and2 gate1324( .a(N5389), .b(N4280), .O(N6075) );
and3 gate1325( .a(N5396), .b(N5389), .c(N4284), .O(N6076) );
and4 gate1326( .a(N5407), .b(N5389), .c(N4290), .d(N5396), .O(N6077) );
and4 gate1327( .a(N5624), .b(N4418), .c(N4445), .d(N4425), .O(N6078) );
inv1 gate1328( .a(N5418), .O(N6079) );
and4 gate1329( .a(N5396), .b(N5418), .c(N5407), .d(N5389), .O(N6080) );
and2 gate1330( .a(N5396), .b(N4284), .O(N6083) );
and3 gate1331( .a(N5407), .b(N4290), .c(N5396), .O(N6084) );
and3 gate1332( .a(N5418), .b(N5407), .c(N5396), .O(N6085) );
and2 gate1333( .a(N5396), .b(N4284), .O(N6086) );
and3 gate1334( .a(N4290), .b(N5407), .c(N5396), .O(N6087) );
and2 gate1335( .a(N5407), .b(N4290), .O(N6088) );
and2 gate1336( .a(N5418), .b(N5407), .O(N6089) );
and2 gate1337( .a(N5407), .b(N4290), .O(N6090) );
and5 gate1338( .a(N5431), .b(N5462), .c(N5441), .d(N5424), .e(N5452), .O(N6091) );
and2 gate1339( .a(N5424), .b(N4298), .O(N6094) );
and3 gate1340( .a(N5431), .b(N5424), .c(N4301), .O(N6095) );
and4 gate1341( .a(N5441), .b(N5424), .c(N4305), .d(N5431), .O(N6096) );
and5 gate1342( .a(N5452), .b(N5441), .c(N5424), .d(N4310), .e(N5431), .O(N6097) );
and2 gate1343( .a(N5431), .b(N4301), .O(N6098) );
and3 gate1344( .a(N5441), .b(N4305), .c(N5431), .O(N6099) );
and4 gate1345( .a(N5452), .b(N5441), .c(N4310), .d(N5431), .O(N6100) );
and5 gate1346( .a(N4), .b(N5462), .c(N5441), .d(N5452), .e(N5431), .O(N6101) );
and2 gate1347( .a(N4305), .b(N5441), .O(N6102) );
and3 gate1348( .a(N5452), .b(N5441), .c(N4310), .O(N6103) );
and4 gate1349( .a(N4), .b(N5462), .c(N5441), .d(N5452), .O(N6104) );
and2 gate1350( .a(N5452), .b(N4310), .O(N6105) );
and3 gate1351( .a(N4), .b(N5462), .c(N5452), .O(N6106) );
and2 gate1352( .a(N4), .b(N5462), .O(N6107) );
and4 gate1353( .a(N5549), .b(N5488), .c(N5477), .d(N5470), .O(N6108) );
and2 gate1354( .a(N5477), .b(N4320), .O(N6111) );
and3 gate1355( .a(N5488), .b(N4325), .c(N5477), .O(N6112) );
and3 gate1356( .a(N5549), .b(N5488), .c(N5477), .O(N6113) );
and2 gate1357( .a(N5477), .b(N4320), .O(N6114) );
and3 gate1358( .a(N5488), .b(N4325), .c(N5477), .O(N6115) );
and2 gate1359( .a(N5488), .b(N4325), .O(N6116) );
and5 gate1360( .a(N5555), .b(N5536), .c(N5520), .d(N5506), .e(N5498), .O(N6117) );
and2 gate1361( .a(N5498), .b(N4332), .O(N6120) );
and3 gate1362( .a(N5506), .b(N5498), .c(N4336), .O(N6121) );
and4 gate1363( .a(N5520), .b(N5498), .c(N4342), .d(N5506), .O(N6122) );
and5 gate1364( .a(N5536), .b(N5520), .c(N5498), .d(N4349), .e(N5506), .O(N6123) );
and2 gate1365( .a(N5506), .b(N4336), .O(N6124) );
and3 gate1366( .a(N5520), .b(N4342), .c(N5506), .O(N6125) );
and4 gate1367( .a(N5536), .b(N5520), .c(N4349), .d(N5506), .O(N6126) );
and4 gate1368( .a(N5555), .b(N5520), .c(N5506), .d(N5536), .O(N6127) );
and2 gate1369( .a(N5506), .b(N4336), .O(N6128) );
and3 gate1370( .a(N5520), .b(N4342), .c(N5506), .O(N6129) );
and4 gate1371( .a(N5536), .b(N5520), .c(N4349), .d(N5506), .O(N6130) );
and2 gate1372( .a(N5520), .b(N4342), .O(N6131) );
and3 gate1373( .a(N5536), .b(N5520), .c(N4349), .O(N6132) );
and3 gate1374( .a(N5555), .b(N5520), .c(N5536), .O(N6133) );
and2 gate1375( .a(N5520), .b(N4342), .O(N6134) );
and3 gate1376( .a(N5536), .b(N5520), .c(N4349), .O(N6135) );
and2 gate1377( .a(N5536), .b(N4349), .O(N6136) );
and2 gate1378( .a(N5549), .b(N5488), .O(N6137) );
and2 gate1379( .a(N5555), .b(N5536), .O(N6138) );
inv1 gate1380( .a(N5573), .O(N6139) );
and4 gate1381( .a(N4364), .b(N5573), .c(N5562), .d(N4357), .O(N6140) );
and3 gate1382( .a(N5562), .b(N4385), .c(N4364), .O(N6143) );
and3 gate1383( .a(N5573), .b(N5562), .c(N4364), .O(N6144) );
and3 gate1384( .a(N4385), .b(N5562), .c(N4364), .O(N6145) );
and2 gate1385( .a(N5562), .b(N4385), .O(N6146) );
and2 gate1386( .a(N5573), .b(N5562), .O(N6147) );
and2 gate1387( .a(N5562), .b(N4385), .O(N6148) );
and5 gate1388( .a(N5264), .b(N4405), .c(N5595), .d(N5579), .e(N5606), .O(N6149) );
and2 gate1389( .a(N5579), .b(N4067), .O(N6152) );
and3 gate1390( .a(N5264), .b(N5579), .c(N4396), .O(N6153) );
and4 gate1391( .a(N5595), .b(N5579), .c(N4400), .d(N5264), .O(N6154) );
and5 gate1392( .a(N5606), .b(N5595), .c(N5579), .d(N4412), .e(N5264), .O(N6155) );
and3 gate1393( .a(N5595), .b(N4400), .c(N5264), .O(N6156) );
and4 gate1394( .a(N5606), .b(N5595), .c(N4412), .d(N5264), .O(N6157) );
and5 gate1395( .a(N54), .b(N4405), .c(N5595), .d(N5606), .e(N5264), .O(N6158) );
and2 gate1396( .a(N4400), .b(N5595), .O(N6159) );
and3 gate1397( .a(N5606), .b(N5595), .c(N4412), .O(N6160) );
and4 gate1398( .a(N54), .b(N4405), .c(N5595), .d(N5606), .O(N6161) );
and2 gate1399( .a(N5606), .b(N4412), .O(N6162) );
and3 gate1400( .a(N54), .b(N4405), .c(N5606), .O(N6163) );

  xor2  gate2308(.a(N5955), .b(N5616), .O(gate1401inter0));
  nand2 gate2309(.a(gate1401inter0), .b(s_0), .O(gate1401inter1));
  and2  gate2310(.a(N5955), .b(N5616), .O(gate1401inter2));
  inv1  gate2311(.a(s_0), .O(gate1401inter3));
  inv1  gate2312(.a(s_1), .O(gate1401inter4));
  nand2 gate2313(.a(gate1401inter4), .b(gate1401inter3), .O(gate1401inter5));
  nor2  gate2314(.a(gate1401inter5), .b(gate1401inter2), .O(gate1401inter6));
  inv1  gate2315(.a(N5616), .O(gate1401inter7));
  inv1  gate2316(.a(N5955), .O(gate1401inter8));
  nand2 gate2317(.a(gate1401inter8), .b(gate1401inter7), .O(gate1401inter9));
  nand2 gate2318(.a(s_1), .b(gate1401inter3), .O(gate1401inter10));
  nor2  gate2319(.a(gate1401inter10), .b(gate1401inter9), .O(gate1401inter11));
  nor2  gate2320(.a(gate1401inter11), .b(gate1401inter6), .O(gate1401inter12));
  nand2 gate2321(.a(gate1401inter12), .b(gate1401inter1), .O(N6164));
and4 gate1402( .a(N5684), .b(N5624), .c(N4425), .d(N4418), .O(N6168) );
and3 gate1403( .a(N5624), .b(N4445), .c(N4425), .O(N6171) );
and3 gate1404( .a(N5684), .b(N5624), .c(N4425), .O(N6172) );
and3 gate1405( .a(N5624), .b(N4445), .c(N4425), .O(N6173) );
and2 gate1406( .a(N5624), .b(N4445), .O(N6174) );
and5 gate1407( .a(N4477), .b(N5671), .c(N5655), .d(N5284), .e(N5634), .O(N6175) );
and2 gate1408( .a(N5634), .b(N4080), .O(N6178) );
and3 gate1409( .a(N5284), .b(N5634), .c(N4456), .O(N6179) );
and4 gate1410( .a(N5655), .b(N5634), .c(N4462), .d(N5284), .O(N6180) );
and5 gate1411( .a(N5671), .b(N5655), .c(N5634), .d(N4469), .e(N5284), .O(N6181) );
and3 gate1412( .a(N5655), .b(N4462), .c(N5284), .O(N6182) );
and4 gate1413( .a(N5671), .b(N5655), .c(N4469), .d(N5284), .O(N6183) );
and4 gate1414( .a(N4477), .b(N5655), .c(N5284), .d(N5671), .O(N6184) );
and3 gate1415( .a(N5655), .b(N4462), .c(N5284), .O(N6185) );
and4 gate1416( .a(N5671), .b(N5655), .c(N4469), .d(N5284), .O(N6186) );
and2 gate1417( .a(N5655), .b(N4462), .O(N6187) );
and3 gate1418( .a(N5671), .b(N5655), .c(N4469), .O(N6188) );
and3 gate1419( .a(N4477), .b(N5655), .c(N5671), .O(N6189) );
and2 gate1420( .a(N5655), .b(N4462), .O(N6190) );
and3 gate1421( .a(N5671), .b(N5655), .c(N4469), .O(N6191) );
and2 gate1422( .a(N5671), .b(N4469), .O(N6192) );
and2 gate1423( .a(N5684), .b(N5624), .O(N6193) );
and2 gate1424( .a(N4477), .b(N5671), .O(N6194) );
inv1 gate1425( .a(N5692), .O(N6197) );
inv1 gate1426( .a(N5696), .O(N6200) );
inv1 gate1427( .a(N5703), .O(N6203) );
inv1 gate1428( .a(N5707), .O(N6206) );
buf1 gate1429( .a(N5700), .O(N6209) );
buf1 gate1430( .a(N5700), .O(N6212) );
buf1 gate1431( .a(N5711), .O(N6215) );
buf1 gate1432( .a(N5711), .O(N6218) );
nand2 gate1433( .a(N5049), .b(N6023), .O(N6221) );
inv1 gate1434( .a(N5756), .O(N6234) );
nand2 gate1435( .a(N5756), .b(N6044), .O(N6235) );
buf1 gate1436( .a(N5462), .O(N6238) );
buf1 gate1437( .a(N5389), .O(N6241) );
buf1 gate1438( .a(N5389), .O(N6244) );
buf1 gate1439( .a(N5396), .O(N6247) );
buf1 gate1440( .a(N5396), .O(N6250) );
buf1 gate1441( .a(N5407), .O(N6253) );
buf1 gate1442( .a(N5407), .O(N6256) );
buf1 gate1443( .a(N5424), .O(N6259) );
buf1 gate1444( .a(N5431), .O(N6262) );
buf1 gate1445( .a(N5441), .O(N6265) );
buf1 gate1446( .a(N5452), .O(N6268) );
buf1 gate1447( .a(N5549), .O(N6271) );
buf1 gate1448( .a(N5488), .O(N6274) );
buf1 gate1449( .a(N5470), .O(N6277) );
buf1 gate1450( .a(N5477), .O(N6280) );
buf1 gate1451( .a(N5549), .O(N6283) );
buf1 gate1452( .a(N5488), .O(N6286) );
buf1 gate1453( .a(N5470), .O(N6289) );
buf1 gate1454( .a(N5477), .O(N6292) );
buf1 gate1455( .a(N5555), .O(N6295) );
buf1 gate1456( .a(N5536), .O(N6298) );
buf1 gate1457( .a(N5498), .O(N6301) );
buf1 gate1458( .a(N5520), .O(N6304) );
buf1 gate1459( .a(N5506), .O(N6307) );
buf1 gate1460( .a(N5506), .O(N6310) );
buf1 gate1461( .a(N5555), .O(N6313) );
buf1 gate1462( .a(N5536), .O(N6316) );
buf1 gate1463( .a(N5498), .O(N6319) );
buf1 gate1464( .a(N5520), .O(N6322) );
buf1 gate1465( .a(N5562), .O(N6325) );
buf1 gate1466( .a(N5562), .O(N6328) );
buf1 gate1467( .a(N5579), .O(N6331) );
buf1 gate1468( .a(N5595), .O(N6335) );
buf1 gate1469( .a(N5606), .O(N6338) );
buf1 gate1470( .a(N5684), .O(N6341) );
buf1 gate1471( .a(N5624), .O(N6344) );
buf1 gate1472( .a(N5684), .O(N6347) );
buf1 gate1473( .a(N5624), .O(N6350) );
buf1 gate1474( .a(N5671), .O(N6353) );
buf1 gate1475( .a(N5634), .O(N6356) );
buf1 gate1476( .a(N5655), .O(N6359) );
buf1 gate1477( .a(N5671), .O(N6364) );
buf1 gate1478( .a(N5634), .O(N6367) );
buf1 gate1479( .a(N5655), .O(N6370) );
inv1 gate1480( .a(N5736), .O(N6373) );
inv1 gate1481( .a(N5739), .O(N6374) );
inv1 gate1482( .a(N5742), .O(N6375) );
inv1 gate1483( .a(N5745), .O(N6376) );
nand2 gate1484( .a(N4243), .b(N6065), .O(N6377) );
nand2 gate1485( .a(N5236), .b(N6068), .O(N6378) );
or4 gate1486( .a(N4268), .b(N6071), .c(N6072), .d(N6073), .O(N6382) );
or4 gate1487( .a(N3968), .b(N5065), .c(N5066), .d(N6074), .O(N6386) );
or4 gate1488( .a(N4271), .b(N6075), .c(N6076), .d(N6077), .O(N6388) );
or4 gate1489( .a(N3968), .b(N5067), .c(N5068), .d(N6078), .O(N6392) );
or5 gate1490( .a(N4297), .b(N6094), .c(N6095), .d(N6096), .e(N6097), .O(N6397) );
or2 gate1491( .a(N4320), .b(N6116), .O(N6411) );
or5 gate1492( .a(N4331), .b(N6120), .c(N6121), .d(N6122), .e(N6123), .O(N6415) );
or2 gate1493( .a(N4342), .b(N6136), .O(N6419) );
or5 gate1494( .a(N4392), .b(N6152), .c(N6153), .d(N6154), .e(N6155), .O(N6427) );
inv1 gate1495( .a(N6048), .O(N6434) );
or2 gate1496( .a(N4440), .b(N6174), .O(N6437) );
or5 gate1497( .a(N4451), .b(N6178), .c(N6179), .d(N6180), .e(N6181), .O(N6441) );
or2 gate1498( .a(N4462), .b(N6192), .O(N6445) );
inv1 gate1499( .a(N6051), .O(N6448) );
inv1 gate1500( .a(N6054), .O(N6449) );
nand2 gate1501( .a(N6221), .b(N6024), .O(N6466) );
inv1 gate1502( .a(N6031), .O(N6469) );
inv1 gate1503( .a(N6034), .O(N6470) );
inv1 gate1504( .a(N6037), .O(N6471) );
inv1 gate1505( .a(N6040), .O(N6472) );
and3 gate1506( .a(N5315), .b(N4524), .c(N6031), .O(N6473) );
and3 gate1507( .a(N6025), .b(N5150), .c(N6034), .O(N6474) );
and3 gate1508( .a(N5324), .b(N4532), .c(N6037), .O(N6475) );
and3 gate1509( .a(N6028), .b(N5157), .c(N6040), .O(N6476) );
nand2 gate1510( .a(N5385), .b(N6234), .O(N6477) );
nand2 gate1511( .a(N6045), .b(N132), .O(N6478) );
or4 gate1512( .a(N4280), .b(N6083), .c(N6084), .d(N6085), .O(N6482) );
nor3 gate1513( .a(N4280), .b(N6086), .c(N6087), .O(N6486) );
or3 gate1514( .a(N4284), .b(N6088), .c(N6089), .O(N6490) );
nor2 gate1515( .a(N4284), .b(N6090), .O(N6494) );
or5 gate1516( .a(N4298), .b(N6098), .c(N6099), .d(N6100), .e(N6101), .O(N6500) );
or4 gate1517( .a(N4301), .b(N6102), .c(N6103), .d(N6104), .O(N6504) );
or3 gate1518( .a(N4305), .b(N6105), .c(N6106), .O(N6508) );
or2 gate1519( .a(N4310), .b(N6107), .O(N6512) );
or4 gate1520( .a(N4316), .b(N6111), .c(N6112), .d(N6113), .O(N6516) );
nor3 gate1521( .a(N4316), .b(N6114), .c(N6115), .O(N6526) );
or4 gate1522( .a(N4336), .b(N6131), .c(N6132), .d(N6133), .O(N6536) );
or5 gate1523( .a(N4332), .b(N6124), .c(N6125), .d(N6126), .e(N6127), .O(N6539) );
nor3 gate1524( .a(N4336), .b(N6134), .c(N6135), .O(N6553) );
nor4 gate1525( .a(N4332), .b(N6128), .c(N6129), .d(N6130), .O(N6556) );
or4 gate1526( .a(N4375), .b(N5117), .c(N6143), .d(N6144), .O(N6566) );
nor3 gate1527( .a(N4375), .b(N5118), .c(N6145), .O(N6569) );
or3 gate1528( .a(N4379), .b(N6146), .c(N6147), .O(N6572) );
nor2 gate1529( .a(N4379), .b(N6148), .O(N6575) );
or5 gate1530( .a(N4067), .b(N5954), .c(N6156), .d(N6157), .e(N6158), .O(N6580) );
or4 gate1531( .a(N4396), .b(N6159), .c(N6160), .d(N6161), .O(N6584) );
or3 gate1532( .a(N4400), .b(N6162), .c(N6163), .O(N6587) );
or4 gate1533( .a(N4436), .b(N5132), .c(N6171), .d(N6172), .O(N6592) );
nor3 gate1534( .a(N4436), .b(N5133), .c(N6173), .O(N6599) );
or4 gate1535( .a(N4456), .b(N6187), .c(N6188), .d(N6189), .O(N6606) );
or5 gate1536( .a(N4080), .b(N6005), .c(N6182), .d(N6183), .e(N6184), .O(N6609) );
nor3 gate1537( .a(N4456), .b(N6190), .c(N6191), .O(N6619) );
nor4 gate1538( .a(N4080), .b(N6006), .c(N6185), .d(N6186), .O(N6622) );
nand2 gate1539( .a(N5739), .b(N6373), .O(N6630) );
nand2 gate1540( .a(N5736), .b(N6374), .O(N6631) );
nand2 gate1541( .a(N5745), .b(N6375), .O(N6632) );
nand2 gate1542( .a(N5742), .b(N6376), .O(N6633) );
nand2 gate1543( .a(N6377), .b(N6066), .O(N6634) );
nand2 gate1544( .a(N6069), .b(N6378), .O(N6637) );
inv1 gate1545( .a(N6164), .O(N6640) );
and2 gate1546( .a(N6108), .b(N6117), .O(N6641) );
and2 gate1547( .a(N6140), .b(N6149), .O(N6643) );
and2 gate1548( .a(N6168), .b(N6175), .O(N6646) );
and2 gate1549( .a(N6080), .b(N6091), .O(N6648) );
nand2 gate1550( .a(N6238), .b(N2637), .O(N6650) );
inv1 gate1551( .a(N6238), .O(N6651) );
inv1 gate1552( .a(N6241), .O(N6653) );
inv1 gate1553( .a(N6244), .O(N6655) );
inv1 gate1554( .a(N6247), .O(N6657) );
inv1 gate1555( .a(N6250), .O(N6659) );
nand2 gate1556( .a(N6253), .b(N5087), .O(N6660) );
inv1 gate1557( .a(N6253), .O(N6661) );

  xor2  gate3722(.a(N5469), .b(N6256), .O(gate1558inter0));
  nand2 gate3723(.a(gate1558inter0), .b(s_202), .O(gate1558inter1));
  and2  gate3724(.a(N5469), .b(N6256), .O(gate1558inter2));
  inv1  gate3725(.a(s_202), .O(gate1558inter3));
  inv1  gate3726(.a(s_203), .O(gate1558inter4));
  nand2 gate3727(.a(gate1558inter4), .b(gate1558inter3), .O(gate1558inter5));
  nor2  gate3728(.a(gate1558inter5), .b(gate1558inter2), .O(gate1558inter6));
  inv1  gate3729(.a(N6256), .O(gate1558inter7));
  inv1  gate3730(.a(N5469), .O(gate1558inter8));
  nand2 gate3731(.a(gate1558inter8), .b(gate1558inter7), .O(gate1558inter9));
  nand2 gate3732(.a(s_203), .b(gate1558inter3), .O(gate1558inter10));
  nor2  gate3733(.a(gate1558inter10), .b(gate1558inter9), .O(gate1558inter11));
  nor2  gate3734(.a(gate1558inter11), .b(gate1558inter6), .O(gate1558inter12));
  nand2 gate3735(.a(gate1558inter12), .b(gate1558inter1), .O(N6662));
inv1 gate1559( .a(N6256), .O(N6663) );
and2 gate1560( .a(N6091), .b(N4), .O(N6664) );
inv1 gate1561( .a(N6259), .O(N6666) );
inv1 gate1562( .a(N6262), .O(N6668) );
inv1 gate1563( .a(N6265), .O(N6670) );
inv1 gate1564( .a(N6268), .O(N6672) );
inv1 gate1565( .a(N6117), .O(N6675) );
inv1 gate1566( .a(N6280), .O(N6680) );
inv1 gate1567( .a(N6292), .O(N6681) );
inv1 gate1568( .a(N6307), .O(N6682) );
inv1 gate1569( .a(N6310), .O(N6683) );
nand2 gate1570( .a(N6325), .b(N5120), .O(N6689) );
inv1 gate1571( .a(N6325), .O(N6690) );
nand2 gate1572( .a(N6328), .b(N5622), .O(N6691) );
inv1 gate1573( .a(N6328), .O(N6692) );
and2 gate1574( .a(N6149), .b(N54), .O(N6693) );
inv1 gate1575( .a(N6331), .O(N6695) );
inv1 gate1576( .a(N6335), .O(N6698) );
nand2 gate1577( .a(N6338), .b(N5956), .O(N6699) );
inv1 gate1578( .a(N6338), .O(N6700) );
inv1 gate1579( .a(N6175), .O(N6703) );
inv1 gate1580( .a(N6209), .O(N6708) );
inv1 gate1581( .a(N6212), .O(N6709) );
inv1 gate1582( .a(N6215), .O(N6710) );
inv1 gate1583( .a(N6218), .O(N6711) );
and3 gate1584( .a(N5696), .b(N5692), .c(N6209), .O(N6712) );
and3 gate1585( .a(N6200), .b(N6197), .c(N6212), .O(N6713) );
and3 gate1586( .a(N5707), .b(N5703), .c(N6215), .O(N6714) );
and3 gate1587( .a(N6206), .b(N6203), .c(N6218), .O(N6715) );
buf1 gate1588( .a(N6466), .O(N6716) );
and3 gate1589( .a(N6164), .b(N1777), .c(N3130), .O(N6718) );
and3 gate1590( .a(N5150), .b(N5315), .c(N6469), .O(N6719) );
and3 gate1591( .a(N4524), .b(N6025), .c(N6470), .O(N6720) );
and3 gate1592( .a(N5157), .b(N5324), .c(N6471), .O(N6721) );
and3 gate1593( .a(N4532), .b(N6028), .c(N6472), .O(N6722) );
nand2 gate1594( .a(N6477), .b(N6235), .O(N6724) );
inv1 gate1595( .a(N6271), .O(N6739) );
inv1 gate1596( .a(N6274), .O(N6740) );
inv1 gate1597( .a(N6277), .O(N6741) );
inv1 gate1598( .a(N6283), .O(N6744) );
inv1 gate1599( .a(N6286), .O(N6745) );
inv1 gate1600( .a(N6289), .O(N6746) );
inv1 gate1601( .a(N6295), .O(N6751) );
inv1 gate1602( .a(N6298), .O(N6752) );
inv1 gate1603( .a(N6301), .O(N6753) );
inv1 gate1604( .a(N6304), .O(N6754) );
inv1 gate1605( .a(N6322), .O(N6755) );
inv1 gate1606( .a(N6313), .O(N6760) );
inv1 gate1607( .a(N6316), .O(N6761) );
inv1 gate1608( .a(N6319), .O(N6762) );
inv1 gate1609( .a(N6341), .O(N6772) );
inv1 gate1610( .a(N6344), .O(N6773) );
inv1 gate1611( .a(N6347), .O(N6776) );
inv1 gate1612( .a(N6350), .O(N6777) );
inv1 gate1613( .a(N6353), .O(N6782) );
inv1 gate1614( .a(N6356), .O(N6783) );
inv1 gate1615( .a(N6359), .O(N6784) );
inv1 gate1616( .a(N6370), .O(N6785) );
inv1 gate1617( .a(N6364), .O(N6790) );
inv1 gate1618( .a(N6367), .O(N6791) );
nand2 gate1619( .a(N6630), .b(N6631), .O(N6792) );
nand2 gate1620( .a(N6632), .b(N6633), .O(N6795) );
and2 gate1621( .a(N6108), .b(N6415), .O(N6801) );
and2 gate1622( .a(N6427), .b(N6140), .O(N6802) );
and2 gate1623( .a(N6397), .b(N6080), .O(N6803) );
and2 gate1624( .a(N6168), .b(N6441), .O(N6804) );
inv1 gate1625( .a(N6466), .O(N6805) );
nand2 gate1626( .a(N1851), .b(N6651), .O(N6806) );
inv1 gate1627( .a(N6482), .O(N6807) );
nand2 gate1628( .a(N6482), .b(N6653), .O(N6808) );
inv1 gate1629( .a(N6486), .O(N6809) );
nand2 gate1630( .a(N6486), .b(N6655), .O(N6810) );
inv1 gate1631( .a(N6490), .O(N6811) );
nand2 gate1632( .a(N6490), .b(N6657), .O(N6812) );
inv1 gate1633( .a(N6494), .O(N6813) );
nand2 gate1634( .a(N6494), .b(N6659), .O(N6814) );

  xor2  gate2756(.a(N6661), .b(N4575), .O(gate1635inter0));
  nand2 gate2757(.a(gate1635inter0), .b(s_64), .O(gate1635inter1));
  and2  gate2758(.a(N6661), .b(N4575), .O(gate1635inter2));
  inv1  gate2759(.a(s_64), .O(gate1635inter3));
  inv1  gate2760(.a(s_65), .O(gate1635inter4));
  nand2 gate2761(.a(gate1635inter4), .b(gate1635inter3), .O(gate1635inter5));
  nor2  gate2762(.a(gate1635inter5), .b(gate1635inter2), .O(gate1635inter6));
  inv1  gate2763(.a(N4575), .O(gate1635inter7));
  inv1  gate2764(.a(N6661), .O(gate1635inter8));
  nand2 gate2765(.a(gate1635inter8), .b(gate1635inter7), .O(gate1635inter9));
  nand2 gate2766(.a(s_65), .b(gate1635inter3), .O(gate1635inter10));
  nor2  gate2767(.a(gate1635inter10), .b(gate1635inter9), .O(gate1635inter11));
  nor2  gate2768(.a(gate1635inter11), .b(gate1635inter6), .O(gate1635inter12));
  nand2 gate2769(.a(gate1635inter12), .b(gate1635inter1), .O(N6815));
nand2 gate1636( .a(N5169), .b(N6663), .O(N6816) );
or2 gate1637( .a(N6397), .b(N6664), .O(N6817) );
inv1 gate1638( .a(N6500), .O(N6823) );
nand2 gate1639( .a(N6500), .b(N6666), .O(N6824) );
inv1 gate1640( .a(N6504), .O(N6825) );
nand2 gate1641( .a(N6504), .b(N6668), .O(N6826) );
inv1 gate1642( .a(N6508), .O(N6827) );
nand2 gate1643( .a(N6508), .b(N6670), .O(N6828) );
inv1 gate1644( .a(N6512), .O(N6829) );
nand2 gate1645( .a(N6512), .b(N6672), .O(N6830) );
inv1 gate1646( .a(N6415), .O(N6831) );
inv1 gate1647( .a(N6566), .O(N6834) );
nand2 gate1648( .a(N6566), .b(N5618), .O(N6835) );
inv1 gate1649( .a(N6569), .O(N6836) );

  xor2  gate2350(.a(N5619), .b(N6569), .O(gate1650inter0));
  nand2 gate2351(.a(gate1650inter0), .b(s_6), .O(gate1650inter1));
  and2  gate2352(.a(N5619), .b(N6569), .O(gate1650inter2));
  inv1  gate2353(.a(s_6), .O(gate1650inter3));
  inv1  gate2354(.a(s_7), .O(gate1650inter4));
  nand2 gate2355(.a(gate1650inter4), .b(gate1650inter3), .O(gate1650inter5));
  nor2  gate2356(.a(gate1650inter5), .b(gate1650inter2), .O(gate1650inter6));
  inv1  gate2357(.a(N6569), .O(gate1650inter7));
  inv1  gate2358(.a(N5619), .O(gate1650inter8));
  nand2 gate2359(.a(gate1650inter8), .b(gate1650inter7), .O(gate1650inter9));
  nand2 gate2360(.a(s_7), .b(gate1650inter3), .O(gate1650inter10));
  nor2  gate2361(.a(gate1650inter10), .b(gate1650inter9), .O(gate1650inter11));
  nor2  gate2362(.a(gate1650inter11), .b(gate1650inter6), .O(gate1650inter12));
  nand2 gate2363(.a(gate1650inter12), .b(gate1650inter1), .O(N6837));
inv1 gate1651( .a(N6572), .O(N6838) );
nand2 gate1652( .a(N6572), .b(N5620), .O(N6839) );
inv1 gate1653( .a(N6575), .O(N6840) );
nand2 gate1654( .a(N6575), .b(N5621), .O(N6841) );
nand2 gate1655( .a(N4627), .b(N6690), .O(N6842) );
nand2 gate1656( .a(N5195), .b(N6692), .O(N6843) );
or2 gate1657( .a(N6427), .b(N6693), .O(N6844) );
inv1 gate1658( .a(N6580), .O(N6850) );
nand2 gate1659( .a(N6580), .b(N6695), .O(N6851) );
inv1 gate1660( .a(N6584), .O(N6852) );
nand2 gate1661( .a(N6584), .b(N6434), .O(N6853) );
inv1 gate1662( .a(N6587), .O(N6854) );
nand2 gate1663( .a(N6587), .b(N6698), .O(N6855) );
nand2 gate1664( .a(N5346), .b(N6700), .O(N6856) );
inv1 gate1665( .a(N6441), .O(N6857) );
and3 gate1666( .a(N6197), .b(N5696), .c(N6708), .O(N6860) );
and3 gate1667( .a(N5692), .b(N6200), .c(N6709), .O(N6861) );
and3 gate1668( .a(N6203), .b(N5707), .c(N6710), .O(N6862) );
and3 gate1669( .a(N5703), .b(N6206), .c(N6711), .O(N6863) );
or3 gate1670( .a(N4197), .b(N6718), .c(N3785), .O(N6866) );

  xor2  gate3540(.a(N6473), .b(N6719), .O(gate1671inter0));
  nand2 gate3541(.a(gate1671inter0), .b(s_176), .O(gate1671inter1));
  and2  gate3542(.a(N6473), .b(N6719), .O(gate1671inter2));
  inv1  gate3543(.a(s_176), .O(gate1671inter3));
  inv1  gate3544(.a(s_177), .O(gate1671inter4));
  nand2 gate3545(.a(gate1671inter4), .b(gate1671inter3), .O(gate1671inter5));
  nor2  gate3546(.a(gate1671inter5), .b(gate1671inter2), .O(gate1671inter6));
  inv1  gate3547(.a(N6719), .O(gate1671inter7));
  inv1  gate3548(.a(N6473), .O(gate1671inter8));
  nand2 gate3549(.a(gate1671inter8), .b(gate1671inter7), .O(gate1671inter9));
  nand2 gate3550(.a(s_177), .b(gate1671inter3), .O(gate1671inter10));
  nor2  gate3551(.a(gate1671inter10), .b(gate1671inter9), .O(gate1671inter11));
  nor2  gate3552(.a(gate1671inter11), .b(gate1671inter6), .O(gate1671inter12));
  nand2 gate3553(.a(gate1671inter12), .b(gate1671inter1), .O(N6872));
nor2 gate1672( .a(N6720), .b(N6474), .O(N6873) );
nor2 gate1673( .a(N6721), .b(N6475), .O(N6874) );

  xor2  gate2994(.a(N6476), .b(N6722), .O(gate1674inter0));
  nand2 gate2995(.a(gate1674inter0), .b(s_98), .O(gate1674inter1));
  and2  gate2996(.a(N6476), .b(N6722), .O(gate1674inter2));
  inv1  gate2997(.a(s_98), .O(gate1674inter3));
  inv1  gate2998(.a(s_99), .O(gate1674inter4));
  nand2 gate2999(.a(gate1674inter4), .b(gate1674inter3), .O(gate1674inter5));
  nor2  gate3000(.a(gate1674inter5), .b(gate1674inter2), .O(gate1674inter6));
  inv1  gate3001(.a(N6722), .O(gate1674inter7));
  inv1  gate3002(.a(N6476), .O(gate1674inter8));
  nand2 gate3003(.a(gate1674inter8), .b(gate1674inter7), .O(gate1674inter9));
  nand2 gate3004(.a(s_99), .b(gate1674inter3), .O(gate1674inter10));
  nor2  gate3005(.a(gate1674inter10), .b(gate1674inter9), .O(gate1674inter11));
  nor2  gate3006(.a(gate1674inter11), .b(gate1674inter6), .O(gate1674inter12));
  nand2 gate3007(.a(gate1674inter12), .b(gate1674inter1), .O(N6875));
inv1 gate1675( .a(N6637), .O(N6876) );
buf1 gate1676( .a(N6724), .O(N6877) );
and2 gate1677( .a(N6045), .b(N6478), .O(N6879) );
and2 gate1678( .a(N6478), .b(N132), .O(N6880) );
or2 gate1679( .a(N6411), .b(N6137), .O(N6881) );
inv1 gate1680( .a(N6516), .O(N6884) );
inv1 gate1681( .a(N6411), .O(N6885) );
inv1 gate1682( .a(N6526), .O(N6888) );
inv1 gate1683( .a(N6536), .O(N6889) );
nand2 gate1684( .a(N6536), .b(N5176), .O(N6890) );
or2 gate1685( .a(N6419), .b(N6138), .O(N6891) );
inv1 gate1686( .a(N6539), .O(N6894) );
inv1 gate1687( .a(N6553), .O(N6895) );
nand2 gate1688( .a(N6553), .b(N5728), .O(N6896) );
inv1 gate1689( .a(N6419), .O(N6897) );
inv1 gate1690( .a(N6556), .O(N6900) );
or2 gate1691( .a(N6437), .b(N6193), .O(N6901) );
inv1 gate1692( .a(N6592), .O(N6904) );
inv1 gate1693( .a(N6437), .O(N6905) );
inv1 gate1694( .a(N6599), .O(N6908) );
or2 gate1695( .a(N6445), .b(N6194), .O(N6909) );
inv1 gate1696( .a(N6606), .O(N6912) );
inv1 gate1697( .a(N6609), .O(N6913) );
inv1 gate1698( .a(N6619), .O(N6914) );
nand2 gate1699( .a(N6619), .b(N5734), .O(N6915) );
inv1 gate1700( .a(N6445), .O(N6916) );
inv1 gate1701( .a(N6622), .O(N6919) );
inv1 gate1702( .a(N6634), .O(N6922) );
nand2 gate1703( .a(N6634), .b(N6067), .O(N6923) );
or2 gate1704( .a(N6382), .b(N6801), .O(N6924) );
or2 gate1705( .a(N6386), .b(N6802), .O(N6925) );
or2 gate1706( .a(N6388), .b(N6803), .O(N6926) );
or2 gate1707( .a(N6392), .b(N6804), .O(N6927) );
inv1 gate1708( .a(N6724), .O(N6930) );
nand2 gate1709( .a(N6650), .b(N6806), .O(N6932) );
nand2 gate1710( .a(N6241), .b(N6807), .O(N6935) );
nand2 gate1711( .a(N6244), .b(N6809), .O(N6936) );
nand2 gate1712( .a(N6247), .b(N6811), .O(N6937) );
nand2 gate1713( .a(N6250), .b(N6813), .O(N6938) );
nand2 gate1714( .a(N6660), .b(N6815), .O(N6939) );
nand2 gate1715( .a(N6662), .b(N6816), .O(N6940) );

  xor2  gate2504(.a(N6823), .b(N6259), .O(gate1716inter0));
  nand2 gate2505(.a(gate1716inter0), .b(s_28), .O(gate1716inter1));
  and2  gate2506(.a(N6823), .b(N6259), .O(gate1716inter2));
  inv1  gate2507(.a(s_28), .O(gate1716inter3));
  inv1  gate2508(.a(s_29), .O(gate1716inter4));
  nand2 gate2509(.a(gate1716inter4), .b(gate1716inter3), .O(gate1716inter5));
  nor2  gate2510(.a(gate1716inter5), .b(gate1716inter2), .O(gate1716inter6));
  inv1  gate2511(.a(N6259), .O(gate1716inter7));
  inv1  gate2512(.a(N6823), .O(gate1716inter8));
  nand2 gate2513(.a(gate1716inter8), .b(gate1716inter7), .O(gate1716inter9));
  nand2 gate2514(.a(s_29), .b(gate1716inter3), .O(gate1716inter10));
  nor2  gate2515(.a(gate1716inter10), .b(gate1716inter9), .O(gate1716inter11));
  nor2  gate2516(.a(gate1716inter11), .b(gate1716inter6), .O(gate1716inter12));
  nand2 gate2517(.a(gate1716inter12), .b(gate1716inter1), .O(N6946));
nand2 gate1717( .a(N6262), .b(N6825), .O(N6947) );
nand2 gate1718( .a(N6265), .b(N6827), .O(N6948) );
nand2 gate1719( .a(N6268), .b(N6829), .O(N6949) );

  xor2  gate2392(.a(N6834), .b(N5183), .O(gate1720inter0));
  nand2 gate2393(.a(gate1720inter0), .b(s_12), .O(gate1720inter1));
  and2  gate2394(.a(N6834), .b(N5183), .O(gate1720inter2));
  inv1  gate2395(.a(s_12), .O(gate1720inter3));
  inv1  gate2396(.a(s_13), .O(gate1720inter4));
  nand2 gate2397(.a(gate1720inter4), .b(gate1720inter3), .O(gate1720inter5));
  nor2  gate2398(.a(gate1720inter5), .b(gate1720inter2), .O(gate1720inter6));
  inv1  gate2399(.a(N5183), .O(gate1720inter7));
  inv1  gate2400(.a(N6834), .O(gate1720inter8));
  nand2 gate2401(.a(gate1720inter8), .b(gate1720inter7), .O(gate1720inter9));
  nand2 gate2402(.a(s_13), .b(gate1720inter3), .O(gate1720inter10));
  nor2  gate2403(.a(gate1720inter10), .b(gate1720inter9), .O(gate1720inter11));
  nor2  gate2404(.a(gate1720inter11), .b(gate1720inter6), .O(gate1720inter12));
  nand2 gate2405(.a(gate1720inter12), .b(gate1720inter1), .O(N6953));

  xor2  gate2546(.a(N6836), .b(N5186), .O(gate1721inter0));
  nand2 gate2547(.a(gate1721inter0), .b(s_34), .O(gate1721inter1));
  and2  gate2548(.a(N6836), .b(N5186), .O(gate1721inter2));
  inv1  gate2549(.a(s_34), .O(gate1721inter3));
  inv1  gate2550(.a(s_35), .O(gate1721inter4));
  nand2 gate2551(.a(gate1721inter4), .b(gate1721inter3), .O(gate1721inter5));
  nor2  gate2552(.a(gate1721inter5), .b(gate1721inter2), .O(gate1721inter6));
  inv1  gate2553(.a(N5186), .O(gate1721inter7));
  inv1  gate2554(.a(N6836), .O(gate1721inter8));
  nand2 gate2555(.a(gate1721inter8), .b(gate1721inter7), .O(gate1721inter9));
  nand2 gate2556(.a(s_35), .b(gate1721inter3), .O(gate1721inter10));
  nor2  gate2557(.a(gate1721inter10), .b(gate1721inter9), .O(gate1721inter11));
  nor2  gate2558(.a(gate1721inter11), .b(gate1721inter6), .O(gate1721inter12));
  nand2 gate2559(.a(gate1721inter12), .b(gate1721inter1), .O(N6954));
nand2 gate1722( .a(N5189), .b(N6838), .O(N6955) );
nand2 gate1723( .a(N5192), .b(N6840), .O(N6956) );
nand2 gate1724( .a(N6689), .b(N6842), .O(N6957) );
nand2 gate1725( .a(N6691), .b(N6843), .O(N6958) );
nand2 gate1726( .a(N6331), .b(N6850), .O(N6964) );
nand2 gate1727( .a(N6048), .b(N6852), .O(N6965) );
nand2 gate1728( .a(N6335), .b(N6854), .O(N6966) );
nand2 gate1729( .a(N6699), .b(N6856), .O(N6967) );
nor2 gate1730( .a(N6860), .b(N6712), .O(N6973) );
nor2 gate1731( .a(N6861), .b(N6713), .O(N6974) );

  xor2  gate3652(.a(N6714), .b(N6862), .O(gate1732inter0));
  nand2 gate3653(.a(gate1732inter0), .b(s_192), .O(gate1732inter1));
  and2  gate3654(.a(N6714), .b(N6862), .O(gate1732inter2));
  inv1  gate3655(.a(s_192), .O(gate1732inter3));
  inv1  gate3656(.a(s_193), .O(gate1732inter4));
  nand2 gate3657(.a(gate1732inter4), .b(gate1732inter3), .O(gate1732inter5));
  nor2  gate3658(.a(gate1732inter5), .b(gate1732inter2), .O(gate1732inter6));
  inv1  gate3659(.a(N6862), .O(gate1732inter7));
  inv1  gate3660(.a(N6714), .O(gate1732inter8));
  nand2 gate3661(.a(gate1732inter8), .b(gate1732inter7), .O(gate1732inter9));
  nand2 gate3662(.a(s_193), .b(gate1732inter3), .O(gate1732inter10));
  nor2  gate3663(.a(gate1732inter10), .b(gate1732inter9), .O(gate1732inter11));
  nor2  gate3664(.a(gate1732inter11), .b(gate1732inter6), .O(gate1732inter12));
  nand2 gate3665(.a(gate1732inter12), .b(gate1732inter1), .O(N6975));
nor2 gate1733( .a(N6863), .b(N6715), .O(N6976) );
inv1 gate1734( .a(N6792), .O(N6977) );
inv1 gate1735( .a(N6795), .O(N6978) );
or2 gate1736( .a(N6879), .b(N6880), .O(N6979) );
nand2 gate1737( .a(N4608), .b(N6889), .O(N6987) );
nand2 gate1738( .a(N5177), .b(N6895), .O(N6990) );
nand2 gate1739( .a(N5217), .b(N6914), .O(N6999) );
nand2 gate1740( .a(N5377), .b(N6922), .O(N7002) );

  xor2  gate3568(.a(N6872), .b(N6873), .O(gate1741inter0));
  nand2 gate3569(.a(gate1741inter0), .b(s_180), .O(gate1741inter1));
  and2  gate3570(.a(N6872), .b(N6873), .O(gate1741inter2));
  inv1  gate3571(.a(s_180), .O(gate1741inter3));
  inv1  gate3572(.a(s_181), .O(gate1741inter4));
  nand2 gate3573(.a(gate1741inter4), .b(gate1741inter3), .O(gate1741inter5));
  nor2  gate3574(.a(gate1741inter5), .b(gate1741inter2), .O(gate1741inter6));
  inv1  gate3575(.a(N6873), .O(gate1741inter7));
  inv1  gate3576(.a(N6872), .O(gate1741inter8));
  nand2 gate3577(.a(gate1741inter8), .b(gate1741inter7), .O(gate1741inter9));
  nand2 gate3578(.a(s_181), .b(gate1741inter3), .O(gate1741inter10));
  nor2  gate3579(.a(gate1741inter10), .b(gate1741inter9), .O(gate1741inter11));
  nor2  gate3580(.a(gate1741inter11), .b(gate1741inter6), .O(gate1741inter12));
  nand2 gate3581(.a(gate1741inter12), .b(gate1741inter1), .O(N7003));
nand2 gate1742( .a(N6875), .b(N6874), .O(N7006) );
and3 gate1743( .a(N6866), .b(N2681), .c(N2692), .O(N7011) );
and3 gate1744( .a(N6866), .b(N2756), .c(N2767), .O(N7012) );
and3 gate1745( .a(N6866), .b(N2779), .c(N2790), .O(N7013) );
inv1 gate1746( .a(N6866), .O(N7015) );
and3 gate1747( .a(N6866), .b(N2801), .c(N2812), .O(N7016) );
nand2 gate1748( .a(N6935), .b(N6808), .O(N7018) );
nand2 gate1749( .a(N6936), .b(N6810), .O(N7019) );
nand2 gate1750( .a(N6937), .b(N6812), .O(N7020) );
nand2 gate1751( .a(N6938), .b(N6814), .O(N7021) );
inv1 gate1752( .a(N6939), .O(N7022) );
inv1 gate1753( .a(N6817), .O(N7023) );
nand2 gate1754( .a(N6946), .b(N6824), .O(N7028) );
nand2 gate1755( .a(N6947), .b(N6826), .O(N7031) );
nand2 gate1756( .a(N6948), .b(N6828), .O(N7034) );

  xor2  gate2602(.a(N6830), .b(N6949), .O(gate1757inter0));
  nand2 gate2603(.a(gate1757inter0), .b(s_42), .O(gate1757inter1));
  and2  gate2604(.a(N6830), .b(N6949), .O(gate1757inter2));
  inv1  gate2605(.a(s_42), .O(gate1757inter3));
  inv1  gate2606(.a(s_43), .O(gate1757inter4));
  nand2 gate2607(.a(gate1757inter4), .b(gate1757inter3), .O(gate1757inter5));
  nor2  gate2608(.a(gate1757inter5), .b(gate1757inter2), .O(gate1757inter6));
  inv1  gate2609(.a(N6949), .O(gate1757inter7));
  inv1  gate2610(.a(N6830), .O(gate1757inter8));
  nand2 gate2611(.a(gate1757inter8), .b(gate1757inter7), .O(gate1757inter9));
  nand2 gate2612(.a(s_43), .b(gate1757inter3), .O(gate1757inter10));
  nor2  gate2613(.a(gate1757inter10), .b(gate1757inter9), .O(gate1757inter11));
  nor2  gate2614(.a(gate1757inter11), .b(gate1757inter6), .O(gate1757inter12));
  nand2 gate2615(.a(gate1757inter12), .b(gate1757inter1), .O(N7037));
and2 gate1758( .a(N6817), .b(N6079), .O(N7040) );
and2 gate1759( .a(N6831), .b(N6675), .O(N7041) );
nand2 gate1760( .a(N6953), .b(N6835), .O(N7044) );
nand2 gate1761( .a(N6954), .b(N6837), .O(N7045) );
nand2 gate1762( .a(N6955), .b(N6839), .O(N7046) );
nand2 gate1763( .a(N6956), .b(N6841), .O(N7047) );
inv1 gate1764( .a(N6957), .O(N7048) );
inv1 gate1765( .a(N6844), .O(N7049) );
nand2 gate1766( .a(N6964), .b(N6851), .O(N7054) );
nand2 gate1767( .a(N6965), .b(N6853), .O(N7057) );
nand2 gate1768( .a(N6966), .b(N6855), .O(N7060) );
and2 gate1769( .a(N6844), .b(N6139), .O(N7064) );
and2 gate1770( .a(N6857), .b(N6703), .O(N7065) );
inv1 gate1771( .a(N6881), .O(N7072) );

  xor2  gate3288(.a(N5172), .b(N6881), .O(gate1772inter0));
  nand2 gate3289(.a(gate1772inter0), .b(s_140), .O(gate1772inter1));
  and2  gate3290(.a(N5172), .b(N6881), .O(gate1772inter2));
  inv1  gate3291(.a(s_140), .O(gate1772inter3));
  inv1  gate3292(.a(s_141), .O(gate1772inter4));
  nand2 gate3293(.a(gate1772inter4), .b(gate1772inter3), .O(gate1772inter5));
  nor2  gate3294(.a(gate1772inter5), .b(gate1772inter2), .O(gate1772inter6));
  inv1  gate3295(.a(N6881), .O(gate1772inter7));
  inv1  gate3296(.a(N5172), .O(gate1772inter8));
  nand2 gate3297(.a(gate1772inter8), .b(gate1772inter7), .O(gate1772inter9));
  nand2 gate3298(.a(s_141), .b(gate1772inter3), .O(gate1772inter10));
  nor2  gate3299(.a(gate1772inter10), .b(gate1772inter9), .O(gate1772inter11));
  nor2  gate3300(.a(gate1772inter11), .b(gate1772inter6), .O(gate1772inter12));
  nand2 gate3301(.a(gate1772inter12), .b(gate1772inter1), .O(N7073));
inv1 gate1773( .a(N6885), .O(N7074) );

  xor2  gate2924(.a(N5727), .b(N6885), .O(gate1774inter0));
  nand2 gate2925(.a(gate1774inter0), .b(s_88), .O(gate1774inter1));
  and2  gate2926(.a(N5727), .b(N6885), .O(gate1774inter2));
  inv1  gate2927(.a(s_88), .O(gate1774inter3));
  inv1  gate2928(.a(s_89), .O(gate1774inter4));
  nand2 gate2929(.a(gate1774inter4), .b(gate1774inter3), .O(gate1774inter5));
  nor2  gate2930(.a(gate1774inter5), .b(gate1774inter2), .O(gate1774inter6));
  inv1  gate2931(.a(N6885), .O(gate1774inter7));
  inv1  gate2932(.a(N5727), .O(gate1774inter8));
  nand2 gate2933(.a(gate1774inter8), .b(gate1774inter7), .O(gate1774inter9));
  nand2 gate2934(.a(s_89), .b(gate1774inter3), .O(gate1774inter10));
  nor2  gate2935(.a(gate1774inter10), .b(gate1774inter9), .O(gate1774inter11));
  nor2  gate2936(.a(gate1774inter11), .b(gate1774inter6), .O(gate1774inter12));
  nand2 gate2937(.a(gate1774inter12), .b(gate1774inter1), .O(N7075));

  xor2  gate3372(.a(N6987), .b(N6890), .O(gate1775inter0));
  nand2 gate3373(.a(gate1775inter0), .b(s_152), .O(gate1775inter1));
  and2  gate3374(.a(N6987), .b(N6890), .O(gate1775inter2));
  inv1  gate3375(.a(s_152), .O(gate1775inter3));
  inv1  gate3376(.a(s_153), .O(gate1775inter4));
  nand2 gate3377(.a(gate1775inter4), .b(gate1775inter3), .O(gate1775inter5));
  nor2  gate3378(.a(gate1775inter5), .b(gate1775inter2), .O(gate1775inter6));
  inv1  gate3379(.a(N6890), .O(gate1775inter7));
  inv1  gate3380(.a(N6987), .O(gate1775inter8));
  nand2 gate3381(.a(gate1775inter8), .b(gate1775inter7), .O(gate1775inter9));
  nand2 gate3382(.a(s_153), .b(gate1775inter3), .O(gate1775inter10));
  nor2  gate3383(.a(gate1775inter10), .b(gate1775inter9), .O(gate1775inter11));
  nor2  gate3384(.a(gate1775inter11), .b(gate1775inter6), .O(gate1775inter12));
  nand2 gate3385(.a(gate1775inter12), .b(gate1775inter1), .O(N7076));
inv1 gate1776( .a(N6891), .O(N7079) );
nand2 gate1777( .a(N6896), .b(N6990), .O(N7080) );
inv1 gate1778( .a(N6897), .O(N7083) );
inv1 gate1779( .a(N6901), .O(N7084) );
nand2 gate1780( .a(N6901), .b(N5198), .O(N7085) );
inv1 gate1781( .a(N6905), .O(N7086) );
nand2 gate1782( .a(N6905), .b(N5731), .O(N7087) );
inv1 gate1783( .a(N6909), .O(N7088) );

  xor2  gate3764(.a(N6912), .b(N6909), .O(gate1784inter0));
  nand2 gate3765(.a(gate1784inter0), .b(s_208), .O(gate1784inter1));
  and2  gate3766(.a(N6912), .b(N6909), .O(gate1784inter2));
  inv1  gate3767(.a(s_208), .O(gate1784inter3));
  inv1  gate3768(.a(s_209), .O(gate1784inter4));
  nand2 gate3769(.a(gate1784inter4), .b(gate1784inter3), .O(gate1784inter5));
  nor2  gate3770(.a(gate1784inter5), .b(gate1784inter2), .O(gate1784inter6));
  inv1  gate3771(.a(N6909), .O(gate1784inter7));
  inv1  gate3772(.a(N6912), .O(gate1784inter8));
  nand2 gate3773(.a(gate1784inter8), .b(gate1784inter7), .O(gate1784inter9));
  nand2 gate3774(.a(s_209), .b(gate1784inter3), .O(gate1784inter10));
  nor2  gate3775(.a(gate1784inter10), .b(gate1784inter9), .O(gate1784inter11));
  nor2  gate3776(.a(gate1784inter11), .b(gate1784inter6), .O(gate1784inter12));
  nand2 gate3777(.a(gate1784inter12), .b(gate1784inter1), .O(N7089));
nand2 gate1785( .a(N6915), .b(N6999), .O(N7090) );
inv1 gate1786( .a(N6916), .O(N7093) );
nand2 gate1787( .a(N6974), .b(N6973), .O(N7094) );

  xor2  gate2686(.a(N6975), .b(N6976), .O(gate1788inter0));
  nand2 gate2687(.a(gate1788inter0), .b(s_54), .O(gate1788inter1));
  and2  gate2688(.a(N6975), .b(N6976), .O(gate1788inter2));
  inv1  gate2689(.a(s_54), .O(gate1788inter3));
  inv1  gate2690(.a(s_55), .O(gate1788inter4));
  nand2 gate2691(.a(gate1788inter4), .b(gate1788inter3), .O(gate1788inter5));
  nor2  gate2692(.a(gate1788inter5), .b(gate1788inter2), .O(gate1788inter6));
  inv1  gate2693(.a(N6976), .O(gate1788inter7));
  inv1  gate2694(.a(N6975), .O(gate1788inter8));
  nand2 gate2695(.a(gate1788inter8), .b(gate1788inter7), .O(gate1788inter9));
  nand2 gate2696(.a(s_55), .b(gate1788inter3), .O(gate1788inter10));
  nor2  gate2697(.a(gate1788inter10), .b(gate1788inter9), .O(gate1788inter11));
  nor2  gate2698(.a(gate1788inter11), .b(gate1788inter6), .O(gate1788inter12));
  nand2 gate2699(.a(gate1788inter12), .b(gate1788inter1), .O(N7097));
nand2 gate1789( .a(N7002), .b(N6923), .O(N7101) );
inv1 gate1790( .a(N6932), .O(N7105) );
inv1 gate1791( .a(N6967), .O(N7110) );
and3 gate1792( .a(N6979), .b(N603), .c(N1755), .O(N7114) );
inv1 gate1793( .a(N7019), .O(N7115) );
inv1 gate1794( .a(N7021), .O(N7116) );
and2 gate1795( .a(N6817), .b(N7018), .O(N7125) );
and2 gate1796( .a(N6817), .b(N7020), .O(N7126) );
and2 gate1797( .a(N6817), .b(N7022), .O(N7127) );
inv1 gate1798( .a(N7045), .O(N7130) );
inv1 gate1799( .a(N7047), .O(N7131) );
and2 gate1800( .a(N6844), .b(N7044), .O(N7139) );
and2 gate1801( .a(N6844), .b(N7046), .O(N7140) );
and2 gate1802( .a(N6844), .b(N7048), .O(N7141) );
and3 gate1803( .a(N6932), .b(N1761), .c(N3108), .O(N7146) );
and3 gate1804( .a(N6967), .b(N1777), .c(N3130), .O(N7147) );
inv1 gate1805( .a(N7003), .O(N7149) );
inv1 gate1806( .a(N7006), .O(N7150) );
nand2 gate1807( .a(N7006), .b(N6876), .O(N7151) );
nand2 gate1808( .a(N4605), .b(N7072), .O(N7152) );
nand2 gate1809( .a(N5173), .b(N7074), .O(N7153) );

  xor2  gate2854(.a(N7084), .b(N4646), .O(gate1810inter0));
  nand2 gate2855(.a(gate1810inter0), .b(s_78), .O(gate1810inter1));
  and2  gate2856(.a(N7084), .b(N4646), .O(gate1810inter2));
  inv1  gate2857(.a(s_78), .O(gate1810inter3));
  inv1  gate2858(.a(s_79), .O(gate1810inter4));
  nand2 gate2859(.a(gate1810inter4), .b(gate1810inter3), .O(gate1810inter5));
  nor2  gate2860(.a(gate1810inter5), .b(gate1810inter2), .O(gate1810inter6));
  inv1  gate2861(.a(N4646), .O(gate1810inter7));
  inv1  gate2862(.a(N7084), .O(gate1810inter8));
  nand2 gate2863(.a(gate1810inter8), .b(gate1810inter7), .O(gate1810inter9));
  nand2 gate2864(.a(s_79), .b(gate1810inter3), .O(gate1810inter10));
  nor2  gate2865(.a(gate1810inter10), .b(gate1810inter9), .O(gate1810inter11));
  nor2  gate2866(.a(gate1810inter11), .b(gate1810inter6), .O(gate1810inter12));
  nand2 gate2867(.a(gate1810inter12), .b(gate1810inter1), .O(N7158));
nand2 gate1811( .a(N5205), .b(N7086), .O(N7159) );
nand2 gate1812( .a(N6606), .b(N7088), .O(N7160) );
inv1 gate1813( .a(N7037), .O(N7166) );
inv1 gate1814( .a(N7034), .O(N7167) );
inv1 gate1815( .a(N7031), .O(N7168) );
inv1 gate1816( .a(N7028), .O(N7169) );
inv1 gate1817( .a(N7060), .O(N7170) );
inv1 gate1818( .a(N7057), .O(N7171) );
inv1 gate1819( .a(N7054), .O(N7172) );
and2 gate1820( .a(N7115), .b(N7023), .O(N7173) );
and2 gate1821( .a(N7116), .b(N7023), .O(N7174) );
and2 gate1822( .a(N6940), .b(N7023), .O(N7175) );
and2 gate1823( .a(N5418), .b(N7023), .O(N7176) );
inv1 gate1824( .a(N7041), .O(N7177) );
and2 gate1825( .a(N7130), .b(N7049), .O(N7178) );
and2 gate1826( .a(N7131), .b(N7049), .O(N7179) );
and2 gate1827( .a(N6958), .b(N7049), .O(N7180) );
and2 gate1828( .a(N5573), .b(N7049), .O(N7181) );
inv1 gate1829( .a(N7065), .O(N7182) );
inv1 gate1830( .a(N7094), .O(N7183) );
nand2 gate1831( .a(N7094), .b(N6977), .O(N7184) );
inv1 gate1832( .a(N7097), .O(N7185) );
nand2 gate1833( .a(N7097), .b(N6978), .O(N7186) );
and3 gate1834( .a(N7037), .b(N1761), .c(N3108), .O(N7187) );
and3 gate1835( .a(N7034), .b(N1761), .c(N3108), .O(N7188) );
and3 gate1836( .a(N7031), .b(N1761), .c(N3108), .O(N7189) );
or3 gate1837( .a(N4956), .b(N7146), .c(N3781), .O(N7190) );
and3 gate1838( .a(N7060), .b(N1777), .c(N3130), .O(N7196) );
and3 gate1839( .a(N7057), .b(N1777), .c(N3130), .O(N7197) );
or3 gate1840( .a(N4960), .b(N7147), .c(N3786), .O(N7198) );
nand2 gate1841( .a(N7101), .b(N7149), .O(N7204) );
inv1 gate1842( .a(N7101), .O(N7205) );
nand2 gate1843( .a(N6637), .b(N7150), .O(N7206) );
and3 gate1844( .a(N7028), .b(N1793), .c(N3158), .O(N7207) );
and3 gate1845( .a(N7054), .b(N1807), .c(N3180), .O(N7208) );
nand2 gate1846( .a(N7073), .b(N7152), .O(N7209) );
nand2 gate1847( .a(N7075), .b(N7153), .O(N7212) );
inv1 gate1848( .a(N7076), .O(N7215) );

  xor2  gate2952(.a(N7079), .b(N7076), .O(gate1849inter0));
  nand2 gate2953(.a(gate1849inter0), .b(s_92), .O(gate1849inter1));
  and2  gate2954(.a(N7079), .b(N7076), .O(gate1849inter2));
  inv1  gate2955(.a(s_92), .O(gate1849inter3));
  inv1  gate2956(.a(s_93), .O(gate1849inter4));
  nand2 gate2957(.a(gate1849inter4), .b(gate1849inter3), .O(gate1849inter5));
  nor2  gate2958(.a(gate1849inter5), .b(gate1849inter2), .O(gate1849inter6));
  inv1  gate2959(.a(N7076), .O(gate1849inter7));
  inv1  gate2960(.a(N7079), .O(gate1849inter8));
  nand2 gate2961(.a(gate1849inter8), .b(gate1849inter7), .O(gate1849inter9));
  nand2 gate2962(.a(s_93), .b(gate1849inter3), .O(gate1849inter10));
  nor2  gate2963(.a(gate1849inter10), .b(gate1849inter9), .O(gate1849inter11));
  nor2  gate2964(.a(gate1849inter11), .b(gate1849inter6), .O(gate1849inter12));
  nand2 gate2965(.a(gate1849inter12), .b(gate1849inter1), .O(N7216));
inv1 gate1850( .a(N7080), .O(N7217) );
nand2 gate1851( .a(N7080), .b(N7083), .O(N7218) );
nand2 gate1852( .a(N7085), .b(N7158), .O(N7219) );
nand2 gate1853( .a(N7087), .b(N7159), .O(N7222) );

  xor2  gate3904(.a(N7160), .b(N7089), .O(gate1854inter0));
  nand2 gate3905(.a(gate1854inter0), .b(s_228), .O(gate1854inter1));
  and2  gate3906(.a(N7160), .b(N7089), .O(gate1854inter2));
  inv1  gate3907(.a(s_228), .O(gate1854inter3));
  inv1  gate3908(.a(s_229), .O(gate1854inter4));
  nand2 gate3909(.a(gate1854inter4), .b(gate1854inter3), .O(gate1854inter5));
  nor2  gate3910(.a(gate1854inter5), .b(gate1854inter2), .O(gate1854inter6));
  inv1  gate3911(.a(N7089), .O(gate1854inter7));
  inv1  gate3912(.a(N7160), .O(gate1854inter8));
  nand2 gate3913(.a(gate1854inter8), .b(gate1854inter7), .O(gate1854inter9));
  nand2 gate3914(.a(s_229), .b(gate1854inter3), .O(gate1854inter10));
  nor2  gate3915(.a(gate1854inter10), .b(gate1854inter9), .O(gate1854inter11));
  nor2  gate3916(.a(gate1854inter11), .b(gate1854inter6), .O(gate1854inter12));
  nand2 gate3917(.a(gate1854inter12), .b(gate1854inter1), .O(N7225));
inv1 gate1855( .a(N7090), .O(N7228) );

  xor2  gate3274(.a(N7093), .b(N7090), .O(gate1856inter0));
  nand2 gate3275(.a(gate1856inter0), .b(s_138), .O(gate1856inter1));
  and2  gate3276(.a(N7093), .b(N7090), .O(gate1856inter2));
  inv1  gate3277(.a(s_138), .O(gate1856inter3));
  inv1  gate3278(.a(s_139), .O(gate1856inter4));
  nand2 gate3279(.a(gate1856inter4), .b(gate1856inter3), .O(gate1856inter5));
  nor2  gate3280(.a(gate1856inter5), .b(gate1856inter2), .O(gate1856inter6));
  inv1  gate3281(.a(N7090), .O(gate1856inter7));
  inv1  gate3282(.a(N7093), .O(gate1856inter8));
  nand2 gate3283(.a(gate1856inter8), .b(gate1856inter7), .O(gate1856inter9));
  nand2 gate3284(.a(s_139), .b(gate1856inter3), .O(gate1856inter10));
  nor2  gate3285(.a(gate1856inter10), .b(gate1856inter9), .O(gate1856inter11));
  nor2  gate3286(.a(gate1856inter11), .b(gate1856inter6), .O(gate1856inter12));
  nand2 gate3287(.a(gate1856inter12), .b(gate1856inter1), .O(N7229));
or2 gate1857( .a(N7173), .b(N7125), .O(N7236) );
or2 gate1858( .a(N7174), .b(N7126), .O(N7239) );
or2 gate1859( .a(N7175), .b(N7127), .O(N7242) );
or2 gate1860( .a(N7176), .b(N7040), .O(N7245) );
or2 gate1861( .a(N7178), .b(N7139), .O(N7250) );
or2 gate1862( .a(N7179), .b(N7140), .O(N7257) );
or2 gate1863( .a(N7180), .b(N7141), .O(N7260) );
or2 gate1864( .a(N7181), .b(N7064), .O(N7263) );

  xor2  gate3834(.a(N7183), .b(N6792), .O(gate1865inter0));
  nand2 gate3835(.a(gate1865inter0), .b(s_218), .O(gate1865inter1));
  and2  gate3836(.a(N7183), .b(N6792), .O(gate1865inter2));
  inv1  gate3837(.a(s_218), .O(gate1865inter3));
  inv1  gate3838(.a(s_219), .O(gate1865inter4));
  nand2 gate3839(.a(gate1865inter4), .b(gate1865inter3), .O(gate1865inter5));
  nor2  gate3840(.a(gate1865inter5), .b(gate1865inter2), .O(gate1865inter6));
  inv1  gate3841(.a(N6792), .O(gate1865inter7));
  inv1  gate3842(.a(N7183), .O(gate1865inter8));
  nand2 gate3843(.a(gate1865inter8), .b(gate1865inter7), .O(gate1865inter9));
  nand2 gate3844(.a(s_219), .b(gate1865inter3), .O(gate1865inter10));
  nor2  gate3845(.a(gate1865inter10), .b(gate1865inter9), .O(gate1865inter11));
  nor2  gate3846(.a(gate1865inter11), .b(gate1865inter6), .O(gate1865inter12));
  nand2 gate3847(.a(gate1865inter12), .b(gate1865inter1), .O(N7268));

  xor2  gate2966(.a(N7185), .b(N6795), .O(gate1866inter0));
  nand2 gate2967(.a(gate1866inter0), .b(s_94), .O(gate1866inter1));
  and2  gate2968(.a(N7185), .b(N6795), .O(gate1866inter2));
  inv1  gate2969(.a(s_94), .O(gate1866inter3));
  inv1  gate2970(.a(s_95), .O(gate1866inter4));
  nand2 gate2971(.a(gate1866inter4), .b(gate1866inter3), .O(gate1866inter5));
  nor2  gate2972(.a(gate1866inter5), .b(gate1866inter2), .O(gate1866inter6));
  inv1  gate2973(.a(N6795), .O(gate1866inter7));
  inv1  gate2974(.a(N7185), .O(gate1866inter8));
  nand2 gate2975(.a(gate1866inter8), .b(gate1866inter7), .O(gate1866inter9));
  nand2 gate2976(.a(s_95), .b(gate1866inter3), .O(gate1866inter10));
  nor2  gate2977(.a(gate1866inter10), .b(gate1866inter9), .O(gate1866inter11));
  nor2  gate2978(.a(gate1866inter11), .b(gate1866inter6), .O(gate1866inter12));
  nand2 gate2979(.a(gate1866inter12), .b(gate1866inter1), .O(N7269));
or3 gate1867( .a(N4957), .b(N7187), .c(N3782), .O(N7270) );
or3 gate1868( .a(N4958), .b(N7188), .c(N3783), .O(N7276) );
or3 gate1869( .a(N4959), .b(N7189), .c(N3784), .O(N7282) );
or3 gate1870( .a(N4961), .b(N7196), .c(N3787), .O(N7288) );
or3 gate1871( .a(N3998), .b(N7197), .c(N3788), .O(N7294) );

  xor2  gate2588(.a(N7205), .b(N7003), .O(gate1872inter0));
  nand2 gate2589(.a(gate1872inter0), .b(s_40), .O(gate1872inter1));
  and2  gate2590(.a(N7205), .b(N7003), .O(gate1872inter2));
  inv1  gate2591(.a(s_40), .O(gate1872inter3));
  inv1  gate2592(.a(s_41), .O(gate1872inter4));
  nand2 gate2593(.a(gate1872inter4), .b(gate1872inter3), .O(gate1872inter5));
  nor2  gate2594(.a(gate1872inter5), .b(gate1872inter2), .O(gate1872inter6));
  inv1  gate2595(.a(N7003), .O(gate1872inter7));
  inv1  gate2596(.a(N7205), .O(gate1872inter8));
  nand2 gate2597(.a(gate1872inter8), .b(gate1872inter7), .O(gate1872inter9));
  nand2 gate2598(.a(s_41), .b(gate1872inter3), .O(gate1872inter10));
  nor2  gate2599(.a(gate1872inter10), .b(gate1872inter9), .O(gate1872inter11));
  nor2  gate2600(.a(gate1872inter11), .b(gate1872inter6), .O(gate1872inter12));
  nand2 gate2601(.a(gate1872inter12), .b(gate1872inter1), .O(N7300));
nand2 gate1873( .a(N7206), .b(N7151), .O(N7301) );
or3 gate1874( .a(N4980), .b(N7207), .c(N3800), .O(N7304) );
or3 gate1875( .a(N4984), .b(N7208), .c(N3805), .O(N7310) );
nand2 gate1876( .a(N6891), .b(N7215), .O(N7320) );
nand2 gate1877( .a(N6897), .b(N7217), .O(N7321) );
nand2 gate1878( .a(N6916), .b(N7228), .O(N7328) );
and3 gate1879( .a(N7190), .b(N1185), .c(N2692), .O(N7338) );
and3 gate1880( .a(N7198), .b(N2681), .c(N2692), .O(N7339) );
and3 gate1881( .a(N7190), .b(N1247), .c(N2767), .O(N7340) );
and3 gate1882( .a(N7198), .b(N2756), .c(N2767), .O(N7341) );
and3 gate1883( .a(N7190), .b(N1327), .c(N2790), .O(N7342) );
and3 gate1884( .a(N7198), .b(N2779), .c(N2790), .O(N7349) );
and3 gate1885( .a(N7198), .b(N2801), .c(N2812), .O(N7357) );
inv1 gate1886( .a(N7198), .O(N7363) );
and3 gate1887( .a(N7190), .b(N1351), .c(N2812), .O(N7364) );
inv1 gate1888( .a(N7190), .O(N7365) );

  xor2  gate3232(.a(N7184), .b(N7268), .O(gate1889inter0));
  nand2 gate3233(.a(gate1889inter0), .b(s_132), .O(gate1889inter1));
  and2  gate3234(.a(N7184), .b(N7268), .O(gate1889inter2));
  inv1  gate3235(.a(s_132), .O(gate1889inter3));
  inv1  gate3236(.a(s_133), .O(gate1889inter4));
  nand2 gate3237(.a(gate1889inter4), .b(gate1889inter3), .O(gate1889inter5));
  nor2  gate3238(.a(gate1889inter5), .b(gate1889inter2), .O(gate1889inter6));
  inv1  gate3239(.a(N7268), .O(gate1889inter7));
  inv1  gate3240(.a(N7184), .O(gate1889inter8));
  nand2 gate3241(.a(gate1889inter8), .b(gate1889inter7), .O(gate1889inter9));
  nand2 gate3242(.a(s_133), .b(gate1889inter3), .O(gate1889inter10));
  nor2  gate3243(.a(gate1889inter10), .b(gate1889inter9), .O(gate1889inter11));
  nor2  gate3244(.a(gate1889inter11), .b(gate1889inter6), .O(gate1889inter12));
  nand2 gate3245(.a(gate1889inter12), .b(gate1889inter1), .O(N7394));
nand2 gate1890( .a(N7269), .b(N7186), .O(N7397) );
nand2 gate1891( .a(N7204), .b(N7300), .O(N7402) );
inv1 gate1892( .a(N7209), .O(N7405) );
nand2 gate1893( .a(N7209), .b(N6884), .O(N7406) );
inv1 gate1894( .a(N7212), .O(N7407) );
nand2 gate1895( .a(N7212), .b(N6888), .O(N7408) );
nand2 gate1896( .a(N7320), .b(N7216), .O(N7409) );
nand2 gate1897( .a(N7321), .b(N7218), .O(N7412) );
inv1 gate1898( .a(N7219), .O(N7415) );
nand2 gate1899( .a(N7219), .b(N6904), .O(N7416) );
inv1 gate1900( .a(N7222), .O(N7417) );
nand2 gate1901( .a(N7222), .b(N6908), .O(N7418) );
inv1 gate1902( .a(N7225), .O(N7419) );
nand2 gate1903( .a(N7225), .b(N6913), .O(N7420) );

  xor2  gate3316(.a(N7229), .b(N7328), .O(gate1904inter0));
  nand2 gate3317(.a(gate1904inter0), .b(s_144), .O(gate1904inter1));
  and2  gate3318(.a(N7229), .b(N7328), .O(gate1904inter2));
  inv1  gate3319(.a(s_144), .O(gate1904inter3));
  inv1  gate3320(.a(s_145), .O(gate1904inter4));
  nand2 gate3321(.a(gate1904inter4), .b(gate1904inter3), .O(gate1904inter5));
  nor2  gate3322(.a(gate1904inter5), .b(gate1904inter2), .O(gate1904inter6));
  inv1  gate3323(.a(N7328), .O(gate1904inter7));
  inv1  gate3324(.a(N7229), .O(gate1904inter8));
  nand2 gate3325(.a(gate1904inter8), .b(gate1904inter7), .O(gate1904inter9));
  nand2 gate3326(.a(s_145), .b(gate1904inter3), .O(gate1904inter10));
  nor2  gate3327(.a(gate1904inter10), .b(gate1904inter9), .O(gate1904inter11));
  nor2  gate3328(.a(gate1904inter11), .b(gate1904inter6), .O(gate1904inter12));
  nand2 gate3329(.a(gate1904inter12), .b(gate1904inter1), .O(N7421));
inv1 gate1905( .a(N7245), .O(N7424) );
inv1 gate1906( .a(N7242), .O(N7425) );
inv1 gate1907( .a(N7239), .O(N7426) );
inv1 gate1908( .a(N7236), .O(N7427) );
inv1 gate1909( .a(N7263), .O(N7428) );
inv1 gate1910( .a(N7260), .O(N7429) );
inv1 gate1911( .a(N7257), .O(N7430) );
inv1 gate1912( .a(N7250), .O(N7431) );
inv1 gate1913( .a(N7250), .O(N7432) );
and3 gate1914( .a(N7310), .b(N2653), .c(N2664), .O(N7433) );
and3 gate1915( .a(N7304), .b(N1161), .c(N2664), .O(N7434) );
or4 gate1916( .a(N7011), .b(N7338), .c(N3621), .d(N2591), .O(N7435) );
and3 gate1917( .a(N7270), .b(N1185), .c(N2692), .O(N7436) );
and3 gate1918( .a(N7288), .b(N2681), .c(N2692), .O(N7437) );
and3 gate1919( .a(N7276), .b(N1185), .c(N2692), .O(N7438) );
and3 gate1920( .a(N7294), .b(N2681), .c(N2692), .O(N7439) );
and3 gate1921( .a(N7282), .b(N1185), .c(N2692), .O(N7440) );
and3 gate1922( .a(N7310), .b(N2728), .c(N2739), .O(N7441) );
and3 gate1923( .a(N7304), .b(N1223), .c(N2739), .O(N7442) );
or4 gate1924( .a(N7012), .b(N7340), .c(N3632), .d(N2600), .O(N7443) );
and3 gate1925( .a(N7270), .b(N1247), .c(N2767), .O(N7444) );
and3 gate1926( .a(N7288), .b(N2756), .c(N2767), .O(N7445) );
and3 gate1927( .a(N7276), .b(N1247), .c(N2767), .O(N7446) );
and3 gate1928( .a(N7294), .b(N2756), .c(N2767), .O(N7447) );
and3 gate1929( .a(N7282), .b(N1247), .c(N2767), .O(N7448) );
or4 gate1930( .a(N7013), .b(N7342), .c(N3641), .d(N2605), .O(N7449) );
and3 gate1931( .a(N7310), .b(N3041), .c(N3052), .O(N7450) );
and3 gate1932( .a(N7304), .b(N1697), .c(N3052), .O(N7451) );
and3 gate1933( .a(N7294), .b(N2779), .c(N2790), .O(N7452) );
and3 gate1934( .a(N7282), .b(N1327), .c(N2790), .O(N7453) );
and3 gate1935( .a(N7288), .b(N2779), .c(N2790), .O(N7454) );
and3 gate1936( .a(N7276), .b(N1327), .c(N2790), .O(N7455) );
and3 gate1937( .a(N7270), .b(N1327), .c(N2790), .O(N7456) );
and3 gate1938( .a(N7310), .b(N3075), .c(N3086), .O(N7457) );
and3 gate1939( .a(N7304), .b(N1731), .c(N3086), .O(N7458) );
and3 gate1940( .a(N7294), .b(N2801), .c(N2812), .O(N7459) );
and3 gate1941( .a(N7282), .b(N1351), .c(N2812), .O(N7460) );
and3 gate1942( .a(N7288), .b(N2801), .c(N2812), .O(N7461) );
and3 gate1943( .a(N7276), .b(N1351), .c(N2812), .O(N7462) );
and3 gate1944( .a(N7270), .b(N1351), .c(N2812), .O(N7463) );
and3 gate1945( .a(N7250), .b(N603), .c(N599), .O(N7464) );
inv1 gate1946( .a(N7310), .O(N7465) );
inv1 gate1947( .a(N7294), .O(N7466) );
inv1 gate1948( .a(N7288), .O(N7467) );
inv1 gate1949( .a(N7301), .O(N7468) );
or4 gate1950( .a(N7016), .b(N7364), .c(N3660), .d(N2626), .O(N7469) );
inv1 gate1951( .a(N7304), .O(N7470) );
inv1 gate1952( .a(N7282), .O(N7471) );
inv1 gate1953( .a(N7276), .O(N7472) );
inv1 gate1954( .a(N7270), .O(N7473) );
buf1 gate1955( .a(N7394), .O(N7474) );
buf1 gate1956( .a(N7397), .O(N7476) );
and2 gate1957( .a(N7301), .b(N3068), .O(N7479) );
and3 gate1958( .a(N7245), .b(N1793), .c(N3158), .O(N7481) );
and3 gate1959( .a(N7242), .b(N1793), .c(N3158), .O(N7482) );
and3 gate1960( .a(N7239), .b(N1793), .c(N3158), .O(N7483) );
and3 gate1961( .a(N7236), .b(N1793), .c(N3158), .O(N7484) );
and3 gate1962( .a(N7263), .b(N1807), .c(N3180), .O(N7485) );
and3 gate1963( .a(N7260), .b(N1807), .c(N3180), .O(N7486) );
and3 gate1964( .a(N7257), .b(N1807), .c(N3180), .O(N7487) );
and3 gate1965( .a(N7250), .b(N1807), .c(N3180), .O(N7488) );
nand2 gate1966( .a(N6979), .b(N7250), .O(N7489) );
nand2 gate1967( .a(N6516), .b(N7405), .O(N7492) );

  xor2  gate2462(.a(N7407), .b(N6526), .O(gate1968inter0));
  nand2 gate2463(.a(gate1968inter0), .b(s_22), .O(gate1968inter1));
  and2  gate2464(.a(N7407), .b(N6526), .O(gate1968inter2));
  inv1  gate2465(.a(s_22), .O(gate1968inter3));
  inv1  gate2466(.a(s_23), .O(gate1968inter4));
  nand2 gate2467(.a(gate1968inter4), .b(gate1968inter3), .O(gate1968inter5));
  nor2  gate2468(.a(gate1968inter5), .b(gate1968inter2), .O(gate1968inter6));
  inv1  gate2469(.a(N6526), .O(gate1968inter7));
  inv1  gate2470(.a(N7407), .O(gate1968inter8));
  nand2 gate2471(.a(gate1968inter8), .b(gate1968inter7), .O(gate1968inter9));
  nand2 gate2472(.a(s_23), .b(gate1968inter3), .O(gate1968inter10));
  nor2  gate2473(.a(gate1968inter10), .b(gate1968inter9), .O(gate1968inter11));
  nor2  gate2474(.a(gate1968inter11), .b(gate1968inter6), .O(gate1968inter12));
  nand2 gate2475(.a(gate1968inter12), .b(gate1968inter1), .O(N7493));
nand2 gate1969( .a(N6592), .b(N7415), .O(N7498) );

  xor2  gate2714(.a(N7417), .b(N6599), .O(gate1970inter0));
  nand2 gate2715(.a(gate1970inter0), .b(s_58), .O(gate1970inter1));
  and2  gate2716(.a(N7417), .b(N6599), .O(gate1970inter2));
  inv1  gate2717(.a(s_58), .O(gate1970inter3));
  inv1  gate2718(.a(s_59), .O(gate1970inter4));
  nand2 gate2719(.a(gate1970inter4), .b(gate1970inter3), .O(gate1970inter5));
  nor2  gate2720(.a(gate1970inter5), .b(gate1970inter2), .O(gate1970inter6));
  inv1  gate2721(.a(N6599), .O(gate1970inter7));
  inv1  gate2722(.a(N7417), .O(gate1970inter8));
  nand2 gate2723(.a(gate1970inter8), .b(gate1970inter7), .O(gate1970inter9));
  nand2 gate2724(.a(s_59), .b(gate1970inter3), .O(gate1970inter10));
  nor2  gate2725(.a(gate1970inter10), .b(gate1970inter9), .O(gate1970inter11));
  nor2  gate2726(.a(gate1970inter11), .b(gate1970inter6), .O(gate1970inter12));
  nand2 gate2727(.a(gate1970inter12), .b(gate1970inter1), .O(N7499));

  xor2  gate3204(.a(N7419), .b(N6609), .O(gate1971inter0));
  nand2 gate3205(.a(gate1971inter0), .b(s_128), .O(gate1971inter1));
  and2  gate3206(.a(N7419), .b(N6609), .O(gate1971inter2));
  inv1  gate3207(.a(s_128), .O(gate1971inter3));
  inv1  gate3208(.a(s_129), .O(gate1971inter4));
  nand2 gate3209(.a(gate1971inter4), .b(gate1971inter3), .O(gate1971inter5));
  nor2  gate3210(.a(gate1971inter5), .b(gate1971inter2), .O(gate1971inter6));
  inv1  gate3211(.a(N6609), .O(gate1971inter7));
  inv1  gate3212(.a(N7419), .O(gate1971inter8));
  nand2 gate3213(.a(gate1971inter8), .b(gate1971inter7), .O(gate1971inter9));
  nand2 gate3214(.a(s_129), .b(gate1971inter3), .O(gate1971inter10));
  nor2  gate3215(.a(gate1971inter10), .b(gate1971inter9), .O(gate1971inter11));
  nor2  gate3216(.a(gate1971inter11), .b(gate1971inter6), .O(gate1971inter12));
  nand2 gate3217(.a(gate1971inter12), .b(gate1971inter1), .O(N7500));
and9 gate1972( .a(N7105), .b(N7166), .c(N7167), .d(N7168), .e(N7169), .f(N7424), .g(N7425), .h(N7426), .i(N7427), .O(N7503) );
and9 gate1973( .a(N6640), .b(N7110), .c(N7170), .d(N7171), .e(N7172), .f(N7428), .g(N7429), .h(N7430), .i(N7431), .O(N7504) );
or4 gate1974( .a(N7433), .b(N7434), .c(N3616), .d(N2585), .O(N7505) );
and2 gate1975( .a(N7435), .b(N2675), .O(N7506) );
or4 gate1976( .a(N7339), .b(N7436), .c(N3622), .d(N2592), .O(N7507) );
or4 gate1977( .a(N7437), .b(N7438), .c(N3623), .d(N2593), .O(N7508) );
or4 gate1978( .a(N7439), .b(N7440), .c(N3624), .d(N2594), .O(N7509) );
or4 gate1979( .a(N7441), .b(N7442), .c(N3627), .d(N2595), .O(N7510) );
and2 gate1980( .a(N7443), .b(N2750), .O(N7511) );
or4 gate1981( .a(N7341), .b(N7444), .c(N3633), .d(N2601), .O(N7512) );
or4 gate1982( .a(N7445), .b(N7446), .c(N3634), .d(N2602), .O(N7513) );
or4 gate1983( .a(N7447), .b(N7448), .c(N3635), .d(N2603), .O(N7514) );
or4 gate1984( .a(N7450), .b(N7451), .c(N3646), .d(N2610), .O(N7515) );
or4 gate1985( .a(N7452), .b(N7453), .c(N3647), .d(N2611), .O(N7516) );
or4 gate1986( .a(N7454), .b(N7455), .c(N3648), .d(N2612), .O(N7517) );
or4 gate1987( .a(N7349), .b(N7456), .c(N3649), .d(N2613), .O(N7518) );
or4 gate1988( .a(N7457), .b(N7458), .c(N3654), .d(N2618), .O(N7519) );
or4 gate1989( .a(N7459), .b(N7460), .c(N3655), .d(N2619), .O(N7520) );
or4 gate1990( .a(N7461), .b(N7462), .c(N3656), .d(N2620), .O(N7521) );
or4 gate1991( .a(N7357), .b(N7463), .c(N3657), .d(N2621), .O(N7522) );
or4 gate1992( .a(N4741), .b(N7114), .c(N2624), .d(N7464), .O(N7525) );
and3 gate1993( .a(N7468), .b(N3119), .c(N3130), .O(N7526) );
inv1 gate1994( .a(N7394), .O(N7527) );
inv1 gate1995( .a(N7397), .O(N7528) );
inv1 gate1996( .a(N7402), .O(N7529) );
and2 gate1997( .a(N7402), .b(N3068), .O(N7530) );
or3 gate1998( .a(N4981), .b(N7481), .c(N3801), .O(N7531) );
or3 gate1999( .a(N4982), .b(N7482), .c(N3802), .O(N7537) );
or3 gate2000( .a(N4983), .b(N7483), .c(N3803), .O(N7543) );
or3 gate2001( .a(N5165), .b(N7484), .c(N3804), .O(N7549) );
or3 gate2002( .a(N4985), .b(N7485), .c(N3806), .O(N7555) );
or3 gate2003( .a(N4986), .b(N7486), .c(N3807), .O(N7561) );
or3 gate2004( .a(N4547), .b(N7487), .c(N3808), .O(N7567) );
or3 gate2005( .a(N4987), .b(N7488), .c(N3809), .O(N7573) );

  xor2  gate3820(.a(N7406), .b(N7492), .O(gate2006inter0));
  nand2 gate3821(.a(gate2006inter0), .b(s_216), .O(gate2006inter1));
  and2  gate3822(.a(N7406), .b(N7492), .O(gate2006inter2));
  inv1  gate3823(.a(s_216), .O(gate2006inter3));
  inv1  gate3824(.a(s_217), .O(gate2006inter4));
  nand2 gate3825(.a(gate2006inter4), .b(gate2006inter3), .O(gate2006inter5));
  nor2  gate3826(.a(gate2006inter5), .b(gate2006inter2), .O(gate2006inter6));
  inv1  gate3827(.a(N7492), .O(gate2006inter7));
  inv1  gate3828(.a(N7406), .O(gate2006inter8));
  nand2 gate3829(.a(gate2006inter8), .b(gate2006inter7), .O(gate2006inter9));
  nand2 gate3830(.a(s_217), .b(gate2006inter3), .O(gate2006inter10));
  nor2  gate3831(.a(gate2006inter10), .b(gate2006inter9), .O(gate2006inter11));
  nor2  gate3832(.a(gate2006inter11), .b(gate2006inter6), .O(gate2006inter12));
  nand2 gate3833(.a(gate2006inter12), .b(gate2006inter1), .O(N7579));

  xor2  gate3848(.a(N7408), .b(N7493), .O(gate2007inter0));
  nand2 gate3849(.a(gate2007inter0), .b(s_220), .O(gate2007inter1));
  and2  gate3850(.a(N7408), .b(N7493), .O(gate2007inter2));
  inv1  gate3851(.a(s_220), .O(gate2007inter3));
  inv1  gate3852(.a(s_221), .O(gate2007inter4));
  nand2 gate3853(.a(gate2007inter4), .b(gate2007inter3), .O(gate2007inter5));
  nor2  gate3854(.a(gate2007inter5), .b(gate2007inter2), .O(gate2007inter6));
  inv1  gate3855(.a(N7493), .O(gate2007inter7));
  inv1  gate3856(.a(N7408), .O(gate2007inter8));
  nand2 gate3857(.a(gate2007inter8), .b(gate2007inter7), .O(gate2007inter9));
  nand2 gate3858(.a(s_221), .b(gate2007inter3), .O(gate2007inter10));
  nor2  gate3859(.a(gate2007inter10), .b(gate2007inter9), .O(gate2007inter11));
  nor2  gate3860(.a(gate2007inter11), .b(gate2007inter6), .O(gate2007inter12));
  nand2 gate3861(.a(gate2007inter12), .b(gate2007inter1), .O(N7582));
inv1 gate2008( .a(N7409), .O(N7585) );
nand2 gate2009( .a(N7409), .b(N6894), .O(N7586) );
inv1 gate2010( .a(N7412), .O(N7587) );
nand2 gate2011( .a(N7412), .b(N6900), .O(N7588) );

  xor2  gate3680(.a(N7416), .b(N7498), .O(gate2012inter0));
  nand2 gate3681(.a(gate2012inter0), .b(s_196), .O(gate2012inter1));
  and2  gate3682(.a(N7416), .b(N7498), .O(gate2012inter2));
  inv1  gate3683(.a(s_196), .O(gate2012inter3));
  inv1  gate3684(.a(s_197), .O(gate2012inter4));
  nand2 gate3685(.a(gate2012inter4), .b(gate2012inter3), .O(gate2012inter5));
  nor2  gate3686(.a(gate2012inter5), .b(gate2012inter2), .O(gate2012inter6));
  inv1  gate3687(.a(N7498), .O(gate2012inter7));
  inv1  gate3688(.a(N7416), .O(gate2012inter8));
  nand2 gate3689(.a(gate2012inter8), .b(gate2012inter7), .O(gate2012inter9));
  nand2 gate3690(.a(s_197), .b(gate2012inter3), .O(gate2012inter10));
  nor2  gate3691(.a(gate2012inter10), .b(gate2012inter9), .O(gate2012inter11));
  nor2  gate3692(.a(gate2012inter11), .b(gate2012inter6), .O(gate2012inter12));
  nand2 gate3693(.a(gate2012inter12), .b(gate2012inter1), .O(N7589));

  xor2  gate3386(.a(N7418), .b(N7499), .O(gate2013inter0));
  nand2 gate3387(.a(gate2013inter0), .b(s_154), .O(gate2013inter1));
  and2  gate3388(.a(N7418), .b(N7499), .O(gate2013inter2));
  inv1  gate3389(.a(s_154), .O(gate2013inter3));
  inv1  gate3390(.a(s_155), .O(gate2013inter4));
  nand2 gate3391(.a(gate2013inter4), .b(gate2013inter3), .O(gate2013inter5));
  nor2  gate3392(.a(gate2013inter5), .b(gate2013inter2), .O(gate2013inter6));
  inv1  gate3393(.a(N7499), .O(gate2013inter7));
  inv1  gate3394(.a(N7418), .O(gate2013inter8));
  nand2 gate3395(.a(gate2013inter8), .b(gate2013inter7), .O(gate2013inter9));
  nand2 gate3396(.a(s_155), .b(gate2013inter3), .O(gate2013inter10));
  nor2  gate3397(.a(gate2013inter10), .b(gate2013inter9), .O(gate2013inter11));
  nor2  gate3398(.a(gate2013inter11), .b(gate2013inter6), .O(gate2013inter12));
  nand2 gate3399(.a(gate2013inter12), .b(gate2013inter1), .O(N7592));

  xor2  gate3694(.a(N7420), .b(N7500), .O(gate2014inter0));
  nand2 gate3695(.a(gate2014inter0), .b(s_198), .O(gate2014inter1));
  and2  gate3696(.a(N7420), .b(N7500), .O(gate2014inter2));
  inv1  gate3697(.a(s_198), .O(gate2014inter3));
  inv1  gate3698(.a(s_199), .O(gate2014inter4));
  nand2 gate3699(.a(gate2014inter4), .b(gate2014inter3), .O(gate2014inter5));
  nor2  gate3700(.a(gate2014inter5), .b(gate2014inter2), .O(gate2014inter6));
  inv1  gate3701(.a(N7500), .O(gate2014inter7));
  inv1  gate3702(.a(N7420), .O(gate2014inter8));
  nand2 gate3703(.a(gate2014inter8), .b(gate2014inter7), .O(gate2014inter9));
  nand2 gate3704(.a(s_199), .b(gate2014inter3), .O(gate2014inter10));
  nor2  gate3705(.a(gate2014inter10), .b(gate2014inter9), .O(gate2014inter11));
  nor2  gate3706(.a(gate2014inter11), .b(gate2014inter6), .O(gate2014inter12));
  nand2 gate3707(.a(gate2014inter12), .b(gate2014inter1), .O(N7595));
inv1 gate2015( .a(N7421), .O(N7598) );

  xor2  gate3400(.a(N6919), .b(N7421), .O(gate2016inter0));
  nand2 gate3401(.a(gate2016inter0), .b(s_156), .O(gate2016inter1));
  and2  gate3402(.a(N6919), .b(N7421), .O(gate2016inter2));
  inv1  gate3403(.a(s_156), .O(gate2016inter3));
  inv1  gate3404(.a(s_157), .O(gate2016inter4));
  nand2 gate3405(.a(gate2016inter4), .b(gate2016inter3), .O(gate2016inter5));
  nor2  gate3406(.a(gate2016inter5), .b(gate2016inter2), .O(gate2016inter6));
  inv1  gate3407(.a(N7421), .O(gate2016inter7));
  inv1  gate3408(.a(N6919), .O(gate2016inter8));
  nand2 gate3409(.a(gate2016inter8), .b(gate2016inter7), .O(gate2016inter9));
  nand2 gate3410(.a(s_157), .b(gate2016inter3), .O(gate2016inter10));
  nor2  gate3411(.a(gate2016inter10), .b(gate2016inter9), .O(gate2016inter11));
  nor2  gate3412(.a(gate2016inter11), .b(gate2016inter6), .O(gate2016inter12));
  nand2 gate3413(.a(gate2016inter12), .b(gate2016inter1), .O(N7599));
and2 gate2017( .a(N7505), .b(N2647), .O(N7600) );
and2 gate2018( .a(N7507), .b(N2675), .O(N7601) );
and2 gate2019( .a(N7508), .b(N2675), .O(N7602) );
and2 gate2020( .a(N7509), .b(N2675), .O(N7603) );
and2 gate2021( .a(N7510), .b(N2722), .O(N7604) );
and2 gate2022( .a(N7512), .b(N2750), .O(N7605) );
and2 gate2023( .a(N7513), .b(N2750), .O(N7606) );
and2 gate2024( .a(N7514), .b(N2750), .O(N7607) );
and2 gate2025( .a(N6979), .b(N7489), .O(N7624) );
and2 gate2026( .a(N7489), .b(N7250), .O(N7625) );
and2 gate2027( .a(N1149), .b(N7525), .O(N7626) );
and5 gate2028( .a(N562), .b(N7527), .c(N7528), .d(N6805), .e(N6930), .O(N7631) );
and3 gate2029( .a(N7529), .b(N3097), .c(N3108), .O(N7636) );
nand2 gate2030( .a(N6539), .b(N7585), .O(N7657) );

  xor2  gate2882(.a(N7587), .b(N6556), .O(gate2031inter0));
  nand2 gate2883(.a(gate2031inter0), .b(s_82), .O(gate2031inter1));
  and2  gate2884(.a(N7587), .b(N6556), .O(gate2031inter2));
  inv1  gate2885(.a(s_82), .O(gate2031inter3));
  inv1  gate2886(.a(s_83), .O(gate2031inter4));
  nand2 gate2887(.a(gate2031inter4), .b(gate2031inter3), .O(gate2031inter5));
  nor2  gate2888(.a(gate2031inter5), .b(gate2031inter2), .O(gate2031inter6));
  inv1  gate2889(.a(N6556), .O(gate2031inter7));
  inv1  gate2890(.a(N7587), .O(gate2031inter8));
  nand2 gate2891(.a(gate2031inter8), .b(gate2031inter7), .O(gate2031inter9));
  nand2 gate2892(.a(s_83), .b(gate2031inter3), .O(gate2031inter10));
  nor2  gate2893(.a(gate2031inter10), .b(gate2031inter9), .O(gate2031inter11));
  nor2  gate2894(.a(gate2031inter11), .b(gate2031inter6), .O(gate2031inter12));
  nand2 gate2895(.a(gate2031inter12), .b(gate2031inter1), .O(N7658));

  xor2  gate2434(.a(N7598), .b(N6622), .O(gate2032inter0));
  nand2 gate2435(.a(gate2032inter0), .b(s_18), .O(gate2032inter1));
  and2  gate2436(.a(N7598), .b(N6622), .O(gate2032inter2));
  inv1  gate2437(.a(s_18), .O(gate2032inter3));
  inv1  gate2438(.a(s_19), .O(gate2032inter4));
  nand2 gate2439(.a(gate2032inter4), .b(gate2032inter3), .O(gate2032inter5));
  nor2  gate2440(.a(gate2032inter5), .b(gate2032inter2), .O(gate2032inter6));
  inv1  gate2441(.a(N6622), .O(gate2032inter7));
  inv1  gate2442(.a(N7598), .O(gate2032inter8));
  nand2 gate2443(.a(gate2032inter8), .b(gate2032inter7), .O(gate2032inter9));
  nand2 gate2444(.a(s_19), .b(gate2032inter3), .O(gate2032inter10));
  nor2  gate2445(.a(gate2032inter10), .b(gate2032inter9), .O(gate2032inter11));
  nor2  gate2446(.a(gate2032inter11), .b(gate2032inter6), .O(gate2032inter12));
  nand2 gate2447(.a(gate2032inter12), .b(gate2032inter1), .O(N7665));
and3 gate2033( .a(N7555), .b(N2653), .c(N2664), .O(N7666) );
and3 gate2034( .a(N7531), .b(N1161), .c(N2664), .O(N7667) );
and3 gate2035( .a(N7561), .b(N2653), .c(N2664), .O(N7668) );
and3 gate2036( .a(N7537), .b(N1161), .c(N2664), .O(N7669) );
and3 gate2037( .a(N7567), .b(N2653), .c(N2664), .O(N7670) );
and3 gate2038( .a(N7543), .b(N1161), .c(N2664), .O(N7671) );
and3 gate2039( .a(N7573), .b(N2653), .c(N2664), .O(N7672) );
and3 gate2040( .a(N7549), .b(N1161), .c(N2664), .O(N7673) );
and3 gate2041( .a(N7555), .b(N2728), .c(N2739), .O(N7674) );
and3 gate2042( .a(N7531), .b(N1223), .c(N2739), .O(N7675) );
and3 gate2043( .a(N7561), .b(N2728), .c(N2739), .O(N7676) );
and3 gate2044( .a(N7537), .b(N1223), .c(N2739), .O(N7677) );
and3 gate2045( .a(N7567), .b(N2728), .c(N2739), .O(N7678) );
and3 gate2046( .a(N7543), .b(N1223), .c(N2739), .O(N7679) );
and3 gate2047( .a(N7573), .b(N2728), .c(N2739), .O(N7680) );
and3 gate2048( .a(N7549), .b(N1223), .c(N2739), .O(N7681) );
and3 gate2049( .a(N7573), .b(N3075), .c(N3086), .O(N7682) );
and3 gate2050( .a(N7549), .b(N1731), .c(N3086), .O(N7683) );
and3 gate2051( .a(N7573), .b(N3041), .c(N3052), .O(N7684) );
and3 gate2052( .a(N7549), .b(N1697), .c(N3052), .O(N7685) );
and3 gate2053( .a(N7567), .b(N3041), .c(N3052), .O(N7686) );
and3 gate2054( .a(N7543), .b(N1697), .c(N3052), .O(N7687) );
and3 gate2055( .a(N7561), .b(N3041), .c(N3052), .O(N7688) );
and3 gate2056( .a(N7537), .b(N1697), .c(N3052), .O(N7689) );
and3 gate2057( .a(N7555), .b(N3041), .c(N3052), .O(N7690) );
and3 gate2058( .a(N7531), .b(N1697), .c(N3052), .O(N7691) );
and3 gate2059( .a(N7567), .b(N3075), .c(N3086), .O(N7692) );
and3 gate2060( .a(N7543), .b(N1731), .c(N3086), .O(N7693) );
and3 gate2061( .a(N7561), .b(N3075), .c(N3086), .O(N7694) );
and3 gate2062( .a(N7537), .b(N1731), .c(N3086), .O(N7695) );
and3 gate2063( .a(N7555), .b(N3075), .c(N3086), .O(N7696) );
and3 gate2064( .a(N7531), .b(N1731), .c(N3086), .O(N7697) );
or2 gate2065( .a(N7624), .b(N7625), .O(N7698) );
inv1 gate2066( .a(N7573), .O(N7699) );
inv1 gate2067( .a(N7567), .O(N7700) );
inv1 gate2068( .a(N7561), .O(N7701) );
inv1 gate2069( .a(N7555), .O(N7702) );
and3 gate2070( .a(N1156), .b(N7631), .c(N245), .O(N7703) );
inv1 gate2071( .a(N7549), .O(N7704) );
inv1 gate2072( .a(N7543), .O(N7705) );
inv1 gate2073( .a(N7537), .O(N7706) );
inv1 gate2074( .a(N7531), .O(N7707) );
inv1 gate2075( .a(N7579), .O(N7708) );
nand2 gate2076( .a(N7579), .b(N6739), .O(N7709) );
inv1 gate2077( .a(N7582), .O(N7710) );
nand2 gate2078( .a(N7582), .b(N6744), .O(N7711) );

  xor2  gate3036(.a(N7586), .b(N7657), .O(gate2079inter0));
  nand2 gate3037(.a(gate2079inter0), .b(s_104), .O(gate2079inter1));
  and2  gate3038(.a(N7586), .b(N7657), .O(gate2079inter2));
  inv1  gate3039(.a(s_104), .O(gate2079inter3));
  inv1  gate3040(.a(s_105), .O(gate2079inter4));
  nand2 gate3041(.a(gate2079inter4), .b(gate2079inter3), .O(gate2079inter5));
  nor2  gate3042(.a(gate2079inter5), .b(gate2079inter2), .O(gate2079inter6));
  inv1  gate3043(.a(N7657), .O(gate2079inter7));
  inv1  gate3044(.a(N7586), .O(gate2079inter8));
  nand2 gate3045(.a(gate2079inter8), .b(gate2079inter7), .O(gate2079inter9));
  nand2 gate3046(.a(s_105), .b(gate2079inter3), .O(gate2079inter10));
  nor2  gate3047(.a(gate2079inter10), .b(gate2079inter9), .O(gate2079inter11));
  nor2  gate3048(.a(gate2079inter11), .b(gate2079inter6), .O(gate2079inter12));
  nand2 gate3049(.a(gate2079inter12), .b(gate2079inter1), .O(N7712));
nand2 gate2080( .a(N7658), .b(N7588), .O(N7715) );
inv1 gate2081( .a(N7589), .O(N7718) );
nand2 gate2082( .a(N7589), .b(N6772), .O(N7719) );
inv1 gate2083( .a(N7592), .O(N7720) );
nand2 gate2084( .a(N7592), .b(N6776), .O(N7721) );
inv1 gate2085( .a(N7595), .O(N7722) );
nand2 gate2086( .a(N7595), .b(N5733), .O(N7723) );
nand2 gate2087( .a(N7665), .b(N7599), .O(N7724) );
or4 gate2088( .a(N7666), .b(N7667), .c(N3617), .d(N2586), .O(N7727) );
or4 gate2089( .a(N7668), .b(N7669), .c(N3618), .d(N2587), .O(N7728) );
or4 gate2090( .a(N7670), .b(N7671), .c(N3619), .d(N2588), .O(N7729) );
or4 gate2091( .a(N7672), .b(N7673), .c(N3620), .d(N2589), .O(N7730) );
or4 gate2092( .a(N7674), .b(N7675), .c(N3628), .d(N2596), .O(N7731) );
or4 gate2093( .a(N7676), .b(N7677), .c(N3629), .d(N2597), .O(N7732) );
or4 gate2094( .a(N7678), .b(N7679), .c(N3630), .d(N2598), .O(N7733) );
or4 gate2095( .a(N7680), .b(N7681), .c(N3631), .d(N2599), .O(N7734) );
or4 gate2096( .a(N7682), .b(N7683), .c(N3638), .d(N2604), .O(N7735) );
or4 gate2097( .a(N7684), .b(N7685), .c(N3642), .d(N2606), .O(N7736) );
or4 gate2098( .a(N7686), .b(N7687), .c(N3643), .d(N2607), .O(N7737) );
or4 gate2099( .a(N7688), .b(N7689), .c(N3644), .d(N2608), .O(N7738) );
or4 gate2100( .a(N7690), .b(N7691), .c(N3645), .d(N2609), .O(N7739) );
or4 gate2101( .a(N7692), .b(N7693), .c(N3651), .d(N2615), .O(N7740) );
or4 gate2102( .a(N7694), .b(N7695), .c(N3652), .d(N2616), .O(N7741) );
or4 gate2103( .a(N7696), .b(N7697), .c(N3653), .d(N2617), .O(N7742) );
nand2 gate2104( .a(N6271), .b(N7708), .O(N7743) );
nand2 gate2105( .a(N6283), .b(N7710), .O(N7744) );

  xor2  gate3456(.a(N7718), .b(N6341), .O(gate2106inter0));
  nand2 gate3457(.a(gate2106inter0), .b(s_164), .O(gate2106inter1));
  and2  gate3458(.a(N7718), .b(N6341), .O(gate2106inter2));
  inv1  gate3459(.a(s_164), .O(gate2106inter3));
  inv1  gate3460(.a(s_165), .O(gate2106inter4));
  nand2 gate3461(.a(gate2106inter4), .b(gate2106inter3), .O(gate2106inter5));
  nor2  gate3462(.a(gate2106inter5), .b(gate2106inter2), .O(gate2106inter6));
  inv1  gate3463(.a(N6341), .O(gate2106inter7));
  inv1  gate3464(.a(N7718), .O(gate2106inter8));
  nand2 gate3465(.a(gate2106inter8), .b(gate2106inter7), .O(gate2106inter9));
  nand2 gate3466(.a(s_165), .b(gate2106inter3), .O(gate2106inter10));
  nor2  gate3467(.a(gate2106inter10), .b(gate2106inter9), .O(gate2106inter11));
  nor2  gate3468(.a(gate2106inter11), .b(gate2106inter6), .O(gate2106inter12));
  nand2 gate3469(.a(gate2106inter12), .b(gate2106inter1), .O(N7749));

  xor2  gate3988(.a(N7720), .b(N6347), .O(gate2107inter0));
  nand2 gate3989(.a(gate2107inter0), .b(s_240), .O(gate2107inter1));
  and2  gate3990(.a(N7720), .b(N6347), .O(gate2107inter2));
  inv1  gate3991(.a(s_240), .O(gate2107inter3));
  inv1  gate3992(.a(s_241), .O(gate2107inter4));
  nand2 gate3993(.a(gate2107inter4), .b(gate2107inter3), .O(gate2107inter5));
  nor2  gate3994(.a(gate2107inter5), .b(gate2107inter2), .O(gate2107inter6));
  inv1  gate3995(.a(N6347), .O(gate2107inter7));
  inv1  gate3996(.a(N7720), .O(gate2107inter8));
  nand2 gate3997(.a(gate2107inter8), .b(gate2107inter7), .O(gate2107inter9));
  nand2 gate3998(.a(s_241), .b(gate2107inter3), .O(gate2107inter10));
  nor2  gate3999(.a(gate2107inter10), .b(gate2107inter9), .O(gate2107inter11));
  nor2  gate4000(.a(gate2107inter11), .b(gate2107inter6), .O(gate2107inter12));
  nand2 gate4001(.a(gate2107inter12), .b(gate2107inter1), .O(N7750));

  xor2  gate3876(.a(N7722), .b(N5214), .O(gate2108inter0));
  nand2 gate3877(.a(gate2108inter0), .b(s_224), .O(gate2108inter1));
  and2  gate3878(.a(N7722), .b(N5214), .O(gate2108inter2));
  inv1  gate3879(.a(s_224), .O(gate2108inter3));
  inv1  gate3880(.a(s_225), .O(gate2108inter4));
  nand2 gate3881(.a(gate2108inter4), .b(gate2108inter3), .O(gate2108inter5));
  nor2  gate3882(.a(gate2108inter5), .b(gate2108inter2), .O(gate2108inter6));
  inv1  gate3883(.a(N5214), .O(gate2108inter7));
  inv1  gate3884(.a(N7722), .O(gate2108inter8));
  nand2 gate3885(.a(gate2108inter8), .b(gate2108inter7), .O(gate2108inter9));
  nand2 gate3886(.a(s_225), .b(gate2108inter3), .O(gate2108inter10));
  nor2  gate3887(.a(gate2108inter10), .b(gate2108inter9), .O(gate2108inter11));
  nor2  gate3888(.a(gate2108inter11), .b(gate2108inter6), .O(gate2108inter12));
  nand2 gate3889(.a(gate2108inter12), .b(gate2108inter1), .O(N7751));
and2 gate2109( .a(N7727), .b(N2647), .O(N7754) );
and2 gate2110( .a(N7728), .b(N2647), .O(N7755) );
and2 gate2111( .a(N7729), .b(N2647), .O(N7756) );
and2 gate2112( .a(N7730), .b(N2647), .O(N7757) );
and2 gate2113( .a(N7731), .b(N2722), .O(N7758) );
and2 gate2114( .a(N7732), .b(N2722), .O(N7759) );
and2 gate2115( .a(N7733), .b(N2722), .O(N7760) );
and2 gate2116( .a(N7734), .b(N2722), .O(N7761) );
nand2 gate2117( .a(N7743), .b(N7709), .O(N7762) );
nand2 gate2118( .a(N7744), .b(N7711), .O(N7765) );
inv1 gate2119( .a(N7712), .O(N7768) );
nand2 gate2120( .a(N7712), .b(N6751), .O(N7769) );
inv1 gate2121( .a(N7715), .O(N7770) );
nand2 gate2122( .a(N7715), .b(N6760), .O(N7771) );

  xor2  gate2896(.a(N7719), .b(N7749), .O(gate2123inter0));
  nand2 gate2897(.a(gate2123inter0), .b(s_84), .O(gate2123inter1));
  and2  gate2898(.a(N7719), .b(N7749), .O(gate2123inter2));
  inv1  gate2899(.a(s_84), .O(gate2123inter3));
  inv1  gate2900(.a(s_85), .O(gate2123inter4));
  nand2 gate2901(.a(gate2123inter4), .b(gate2123inter3), .O(gate2123inter5));
  nor2  gate2902(.a(gate2123inter5), .b(gate2123inter2), .O(gate2123inter6));
  inv1  gate2903(.a(N7749), .O(gate2123inter7));
  inv1  gate2904(.a(N7719), .O(gate2123inter8));
  nand2 gate2905(.a(gate2123inter8), .b(gate2123inter7), .O(gate2123inter9));
  nand2 gate2906(.a(s_85), .b(gate2123inter3), .O(gate2123inter10));
  nor2  gate2907(.a(gate2123inter10), .b(gate2123inter9), .O(gate2123inter11));
  nor2  gate2908(.a(gate2123inter11), .b(gate2123inter6), .O(gate2123inter12));
  nand2 gate2909(.a(gate2123inter12), .b(gate2123inter1), .O(N7772));

  xor2  gate3638(.a(N7721), .b(N7750), .O(gate2124inter0));
  nand2 gate3639(.a(gate2124inter0), .b(s_190), .O(gate2124inter1));
  and2  gate3640(.a(N7721), .b(N7750), .O(gate2124inter2));
  inv1  gate3641(.a(s_190), .O(gate2124inter3));
  inv1  gate3642(.a(s_191), .O(gate2124inter4));
  nand2 gate3643(.a(gate2124inter4), .b(gate2124inter3), .O(gate2124inter5));
  nor2  gate3644(.a(gate2124inter5), .b(gate2124inter2), .O(gate2124inter6));
  inv1  gate3645(.a(N7750), .O(gate2124inter7));
  inv1  gate3646(.a(N7721), .O(gate2124inter8));
  nand2 gate3647(.a(gate2124inter8), .b(gate2124inter7), .O(gate2124inter9));
  nand2 gate3648(.a(s_191), .b(gate2124inter3), .O(gate2124inter10));
  nor2  gate3649(.a(gate2124inter10), .b(gate2124inter9), .O(gate2124inter11));
  nor2  gate3650(.a(gate2124inter11), .b(gate2124inter6), .O(gate2124inter12));
  nand2 gate3651(.a(gate2124inter12), .b(gate2124inter1), .O(N7775));
nand2 gate2125( .a(N7751), .b(N7723), .O(N7778) );
inv1 gate2126( .a(N7724), .O(N7781) );
nand2 gate2127( .a(N7724), .b(N5735), .O(N7782) );
nand2 gate2128( .a(N6295), .b(N7768), .O(N7787) );
nand2 gate2129( .a(N6313), .b(N7770), .O(N7788) );
nand2 gate2130( .a(N5220), .b(N7781), .O(N7795) );
inv1 gate2131( .a(N7762), .O(N7796) );
nand2 gate2132( .a(N7762), .b(N6740), .O(N7797) );
inv1 gate2133( .a(N7765), .O(N7798) );

  xor2  gate3806(.a(N6745), .b(N7765), .O(gate2134inter0));
  nand2 gate3807(.a(gate2134inter0), .b(s_214), .O(gate2134inter1));
  and2  gate3808(.a(N6745), .b(N7765), .O(gate2134inter2));
  inv1  gate3809(.a(s_214), .O(gate2134inter3));
  inv1  gate3810(.a(s_215), .O(gate2134inter4));
  nand2 gate3811(.a(gate2134inter4), .b(gate2134inter3), .O(gate2134inter5));
  nor2  gate3812(.a(gate2134inter5), .b(gate2134inter2), .O(gate2134inter6));
  inv1  gate3813(.a(N7765), .O(gate2134inter7));
  inv1  gate3814(.a(N6745), .O(gate2134inter8));
  nand2 gate3815(.a(gate2134inter8), .b(gate2134inter7), .O(gate2134inter9));
  nand2 gate3816(.a(s_215), .b(gate2134inter3), .O(gate2134inter10));
  nor2  gate3817(.a(gate2134inter10), .b(gate2134inter9), .O(gate2134inter11));
  nor2  gate3818(.a(gate2134inter11), .b(gate2134inter6), .O(gate2134inter12));
  nand2 gate3819(.a(gate2134inter12), .b(gate2134inter1), .O(N7799));
nand2 gate2135( .a(N7787), .b(N7769), .O(N7800) );
nand2 gate2136( .a(N7788), .b(N7771), .O(N7803) );
inv1 gate2137( .a(N7772), .O(N7806) );

  xor2  gate3106(.a(N6773), .b(N7772), .O(gate2138inter0));
  nand2 gate3107(.a(gate2138inter0), .b(s_114), .O(gate2138inter1));
  and2  gate3108(.a(N6773), .b(N7772), .O(gate2138inter2));
  inv1  gate3109(.a(s_114), .O(gate2138inter3));
  inv1  gate3110(.a(s_115), .O(gate2138inter4));
  nand2 gate3111(.a(gate2138inter4), .b(gate2138inter3), .O(gate2138inter5));
  nor2  gate3112(.a(gate2138inter5), .b(gate2138inter2), .O(gate2138inter6));
  inv1  gate3113(.a(N7772), .O(gate2138inter7));
  inv1  gate3114(.a(N6773), .O(gate2138inter8));
  nand2 gate3115(.a(gate2138inter8), .b(gate2138inter7), .O(gate2138inter9));
  nand2 gate3116(.a(s_115), .b(gate2138inter3), .O(gate2138inter10));
  nor2  gate3117(.a(gate2138inter10), .b(gate2138inter9), .O(gate2138inter11));
  nor2  gate3118(.a(gate2138inter11), .b(gate2138inter6), .O(gate2138inter12));
  nand2 gate3119(.a(gate2138inter12), .b(gate2138inter1), .O(N7807));
inv1 gate2139( .a(N7775), .O(N7808) );

  xor2  gate2532(.a(N6777), .b(N7775), .O(gate2140inter0));
  nand2 gate2533(.a(gate2140inter0), .b(s_32), .O(gate2140inter1));
  and2  gate2534(.a(N6777), .b(N7775), .O(gate2140inter2));
  inv1  gate2535(.a(s_32), .O(gate2140inter3));
  inv1  gate2536(.a(s_33), .O(gate2140inter4));
  nand2 gate2537(.a(gate2140inter4), .b(gate2140inter3), .O(gate2140inter5));
  nor2  gate2538(.a(gate2140inter5), .b(gate2140inter2), .O(gate2140inter6));
  inv1  gate2539(.a(N7775), .O(gate2140inter7));
  inv1  gate2540(.a(N6777), .O(gate2140inter8));
  nand2 gate2541(.a(gate2140inter8), .b(gate2140inter7), .O(gate2140inter9));
  nand2 gate2542(.a(s_33), .b(gate2140inter3), .O(gate2140inter10));
  nor2  gate2543(.a(gate2140inter10), .b(gate2140inter9), .O(gate2140inter11));
  nor2  gate2544(.a(gate2140inter11), .b(gate2140inter6), .O(gate2140inter12));
  nand2 gate2545(.a(gate2140inter12), .b(gate2140inter1), .O(N7809));
inv1 gate2141( .a(N7778), .O(N7810) );
nand2 gate2142( .a(N7778), .b(N6782), .O(N7811) );

  xor2  gate3008(.a(N7782), .b(N7795), .O(gate2143inter0));
  nand2 gate3009(.a(gate2143inter0), .b(s_100), .O(gate2143inter1));
  and2  gate3010(.a(N7782), .b(N7795), .O(gate2143inter2));
  inv1  gate3011(.a(s_100), .O(gate2143inter3));
  inv1  gate3012(.a(s_101), .O(gate2143inter4));
  nand2 gate3013(.a(gate2143inter4), .b(gate2143inter3), .O(gate2143inter5));
  nor2  gate3014(.a(gate2143inter5), .b(gate2143inter2), .O(gate2143inter6));
  inv1  gate3015(.a(N7795), .O(gate2143inter7));
  inv1  gate3016(.a(N7782), .O(gate2143inter8));
  nand2 gate3017(.a(gate2143inter8), .b(gate2143inter7), .O(gate2143inter9));
  nand2 gate3018(.a(s_101), .b(gate2143inter3), .O(gate2143inter10));
  nor2  gate3019(.a(gate2143inter10), .b(gate2143inter9), .O(gate2143inter11));
  nor2  gate3020(.a(gate2143inter11), .b(gate2143inter6), .O(gate2143inter12));
  nand2 gate3021(.a(gate2143inter12), .b(gate2143inter1), .O(N7812));
nand2 gate2144( .a(N6274), .b(N7796), .O(N7815) );
nand2 gate2145( .a(N6286), .b(N7798), .O(N7816) );
nand2 gate2146( .a(N6344), .b(N7806), .O(N7821) );
nand2 gate2147( .a(N6350), .b(N7808), .O(N7822) );
nand2 gate2148( .a(N6353), .b(N7810), .O(N7823) );
nand2 gate2149( .a(N7815), .b(N7797), .O(N7826) );
nand2 gate2150( .a(N7816), .b(N7799), .O(N7829) );
inv1 gate2151( .a(N7800), .O(N7832) );
nand2 gate2152( .a(N7800), .b(N6752), .O(N7833) );
inv1 gate2153( .a(N7803), .O(N7834) );
nand2 gate2154( .a(N7803), .b(N6761), .O(N7835) );

  xor2  gate3414(.a(N7807), .b(N7821), .O(gate2155inter0));
  nand2 gate3415(.a(gate2155inter0), .b(s_158), .O(gate2155inter1));
  and2  gate3416(.a(N7807), .b(N7821), .O(gate2155inter2));
  inv1  gate3417(.a(s_158), .O(gate2155inter3));
  inv1  gate3418(.a(s_159), .O(gate2155inter4));
  nand2 gate3419(.a(gate2155inter4), .b(gate2155inter3), .O(gate2155inter5));
  nor2  gate3420(.a(gate2155inter5), .b(gate2155inter2), .O(gate2155inter6));
  inv1  gate3421(.a(N7821), .O(gate2155inter7));
  inv1  gate3422(.a(N7807), .O(gate2155inter8));
  nand2 gate3423(.a(gate2155inter8), .b(gate2155inter7), .O(gate2155inter9));
  nand2 gate3424(.a(s_159), .b(gate2155inter3), .O(gate2155inter10));
  nor2  gate3425(.a(gate2155inter10), .b(gate2155inter9), .O(gate2155inter11));
  nor2  gate3426(.a(gate2155inter11), .b(gate2155inter6), .O(gate2155inter12));
  nand2 gate3427(.a(gate2155inter12), .b(gate2155inter1), .O(N7836));
nand2 gate2156( .a(N7822), .b(N7809), .O(N7839) );

  xor2  gate2630(.a(N7811), .b(N7823), .O(gate2157inter0));
  nand2 gate2631(.a(gate2157inter0), .b(s_46), .O(gate2157inter1));
  and2  gate2632(.a(N7811), .b(N7823), .O(gate2157inter2));
  inv1  gate2633(.a(s_46), .O(gate2157inter3));
  inv1  gate2634(.a(s_47), .O(gate2157inter4));
  nand2 gate2635(.a(gate2157inter4), .b(gate2157inter3), .O(gate2157inter5));
  nor2  gate2636(.a(gate2157inter5), .b(gate2157inter2), .O(gate2157inter6));
  inv1  gate2637(.a(N7823), .O(gate2157inter7));
  inv1  gate2638(.a(N7811), .O(gate2157inter8));
  nand2 gate2639(.a(gate2157inter8), .b(gate2157inter7), .O(gate2157inter9));
  nand2 gate2640(.a(s_47), .b(gate2157inter3), .O(gate2157inter10));
  nor2  gate2641(.a(gate2157inter10), .b(gate2157inter9), .O(gate2157inter11));
  nor2  gate2642(.a(gate2157inter11), .b(gate2157inter6), .O(gate2157inter12));
  nand2 gate2643(.a(gate2157inter12), .b(gate2157inter1), .O(N7842));
inv1 gate2158( .a(N7812), .O(N7845) );

  xor2  gate3498(.a(N6790), .b(N7812), .O(gate2159inter0));
  nand2 gate3499(.a(gate2159inter0), .b(s_170), .O(gate2159inter1));
  and2  gate3500(.a(N6790), .b(N7812), .O(gate2159inter2));
  inv1  gate3501(.a(s_170), .O(gate2159inter3));
  inv1  gate3502(.a(s_171), .O(gate2159inter4));
  nand2 gate3503(.a(gate2159inter4), .b(gate2159inter3), .O(gate2159inter5));
  nor2  gate3504(.a(gate2159inter5), .b(gate2159inter2), .O(gate2159inter6));
  inv1  gate3505(.a(N7812), .O(gate2159inter7));
  inv1  gate3506(.a(N6790), .O(gate2159inter8));
  nand2 gate3507(.a(gate2159inter8), .b(gate2159inter7), .O(gate2159inter9));
  nand2 gate3508(.a(s_171), .b(gate2159inter3), .O(gate2159inter10));
  nor2  gate3509(.a(gate2159inter10), .b(gate2159inter9), .O(gate2159inter11));
  nor2  gate3510(.a(gate2159inter11), .b(gate2159inter6), .O(gate2159inter12));
  nand2 gate3511(.a(gate2159inter12), .b(gate2159inter1), .O(N7846));
nand2 gate2160( .a(N6298), .b(N7832), .O(N7851) );

  xor2  gate2784(.a(N7834), .b(N6316), .O(gate2161inter0));
  nand2 gate2785(.a(gate2161inter0), .b(s_68), .O(gate2161inter1));
  and2  gate2786(.a(N7834), .b(N6316), .O(gate2161inter2));
  inv1  gate2787(.a(s_68), .O(gate2161inter3));
  inv1  gate2788(.a(s_69), .O(gate2161inter4));
  nand2 gate2789(.a(gate2161inter4), .b(gate2161inter3), .O(gate2161inter5));
  nor2  gate2790(.a(gate2161inter5), .b(gate2161inter2), .O(gate2161inter6));
  inv1  gate2791(.a(N6316), .O(gate2161inter7));
  inv1  gate2792(.a(N7834), .O(gate2161inter8));
  nand2 gate2793(.a(gate2161inter8), .b(gate2161inter7), .O(gate2161inter9));
  nand2 gate2794(.a(s_69), .b(gate2161inter3), .O(gate2161inter10));
  nor2  gate2795(.a(gate2161inter10), .b(gate2161inter9), .O(gate2161inter11));
  nor2  gate2796(.a(gate2161inter11), .b(gate2161inter6), .O(gate2161inter12));
  nand2 gate2797(.a(gate2161inter12), .b(gate2161inter1), .O(N7852));
nand2 gate2162( .a(N6364), .b(N7845), .O(N7859) );
inv1 gate2163( .a(N7826), .O(N7860) );
nand2 gate2164( .a(N7826), .b(N6741), .O(N7861) );
inv1 gate2165( .a(N7829), .O(N7862) );
nand2 gate2166( .a(N7829), .b(N6746), .O(N7863) );

  xor2  gate3092(.a(N7833), .b(N7851), .O(gate2167inter0));
  nand2 gate3093(.a(gate2167inter0), .b(s_112), .O(gate2167inter1));
  and2  gate3094(.a(N7833), .b(N7851), .O(gate2167inter2));
  inv1  gate3095(.a(s_112), .O(gate2167inter3));
  inv1  gate3096(.a(s_113), .O(gate2167inter4));
  nand2 gate3097(.a(gate2167inter4), .b(gate2167inter3), .O(gate2167inter5));
  nor2  gate3098(.a(gate2167inter5), .b(gate2167inter2), .O(gate2167inter6));
  inv1  gate3099(.a(N7851), .O(gate2167inter7));
  inv1  gate3100(.a(N7833), .O(gate2167inter8));
  nand2 gate3101(.a(gate2167inter8), .b(gate2167inter7), .O(gate2167inter9));
  nand2 gate3102(.a(s_113), .b(gate2167inter3), .O(gate2167inter10));
  nor2  gate3103(.a(gate2167inter10), .b(gate2167inter9), .O(gate2167inter11));
  nor2  gate3104(.a(gate2167inter11), .b(gate2167inter6), .O(gate2167inter12));
  nand2 gate3105(.a(gate2167inter12), .b(gate2167inter1), .O(N7864));
nand2 gate2168( .a(N7852), .b(N7835), .O(N7867) );
inv1 gate2169( .a(N7836), .O(N7870) );

  xor2  gate3134(.a(N5730), .b(N7836), .O(gate2170inter0));
  nand2 gate3135(.a(gate2170inter0), .b(s_118), .O(gate2170inter1));
  and2  gate3136(.a(N5730), .b(N7836), .O(gate2170inter2));
  inv1  gate3137(.a(s_118), .O(gate2170inter3));
  inv1  gate3138(.a(s_119), .O(gate2170inter4));
  nand2 gate3139(.a(gate2170inter4), .b(gate2170inter3), .O(gate2170inter5));
  nor2  gate3140(.a(gate2170inter5), .b(gate2170inter2), .O(gate2170inter6));
  inv1  gate3141(.a(N7836), .O(gate2170inter7));
  inv1  gate3142(.a(N5730), .O(gate2170inter8));
  nand2 gate3143(.a(gate2170inter8), .b(gate2170inter7), .O(gate2170inter9));
  nand2 gate3144(.a(s_119), .b(gate2170inter3), .O(gate2170inter10));
  nor2  gate3145(.a(gate2170inter10), .b(gate2170inter9), .O(gate2170inter11));
  nor2  gate3146(.a(gate2170inter11), .b(gate2170inter6), .O(gate2170inter12));
  nand2 gate3147(.a(gate2170inter12), .b(gate2170inter1), .O(N7871));
inv1 gate2171( .a(N7839), .O(N7872) );

  xor2  gate3120(.a(N5732), .b(N7839), .O(gate2172inter0));
  nand2 gate3121(.a(gate2172inter0), .b(s_116), .O(gate2172inter1));
  and2  gate3122(.a(N5732), .b(N7839), .O(gate2172inter2));
  inv1  gate3123(.a(s_116), .O(gate2172inter3));
  inv1  gate3124(.a(s_117), .O(gate2172inter4));
  nand2 gate3125(.a(gate2172inter4), .b(gate2172inter3), .O(gate2172inter5));
  nor2  gate3126(.a(gate2172inter5), .b(gate2172inter2), .O(gate2172inter6));
  inv1  gate3127(.a(N7839), .O(gate2172inter7));
  inv1  gate3128(.a(N5732), .O(gate2172inter8));
  nand2 gate3129(.a(gate2172inter8), .b(gate2172inter7), .O(gate2172inter9));
  nand2 gate3130(.a(s_117), .b(gate2172inter3), .O(gate2172inter10));
  nor2  gate3131(.a(gate2172inter10), .b(gate2172inter9), .O(gate2172inter11));
  nor2  gate3132(.a(gate2172inter11), .b(gate2172inter6), .O(gate2172inter12));
  nand2 gate3133(.a(gate2172inter12), .b(gate2172inter1), .O(N7873));
inv1 gate2173( .a(N7842), .O(N7874) );
nand2 gate2174( .a(N7842), .b(N6783), .O(N7875) );
nand2 gate2175( .a(N7859), .b(N7846), .O(N7876) );

  xor2  gate2700(.a(N7860), .b(N6277), .O(gate2176inter0));
  nand2 gate2701(.a(gate2176inter0), .b(s_56), .O(gate2176inter1));
  and2  gate2702(.a(N7860), .b(N6277), .O(gate2176inter2));
  inv1  gate2703(.a(s_56), .O(gate2176inter3));
  inv1  gate2704(.a(s_57), .O(gate2176inter4));
  nand2 gate2705(.a(gate2176inter4), .b(gate2176inter3), .O(gate2176inter5));
  nor2  gate2706(.a(gate2176inter5), .b(gate2176inter2), .O(gate2176inter6));
  inv1  gate2707(.a(N6277), .O(gate2176inter7));
  inv1  gate2708(.a(N7860), .O(gate2176inter8));
  nand2 gate2709(.a(gate2176inter8), .b(gate2176inter7), .O(gate2176inter9));
  nand2 gate2710(.a(s_57), .b(gate2176inter3), .O(gate2176inter10));
  nor2  gate2711(.a(gate2176inter10), .b(gate2176inter9), .O(gate2176inter11));
  nor2  gate2712(.a(gate2176inter11), .b(gate2176inter6), .O(gate2176inter12));
  nand2 gate2713(.a(gate2176inter12), .b(gate2176inter1), .O(N7879));
nand2 gate2177( .a(N6289), .b(N7862), .O(N7880) );
nand2 gate2178( .a(N5199), .b(N7870), .O(N7885) );

  xor2  gate3428(.a(N7872), .b(N5208), .O(gate2179inter0));
  nand2 gate3429(.a(gate2179inter0), .b(s_160), .O(gate2179inter1));
  and2  gate3430(.a(N7872), .b(N5208), .O(gate2179inter2));
  inv1  gate3431(.a(s_160), .O(gate2179inter3));
  inv1  gate3432(.a(s_161), .O(gate2179inter4));
  nand2 gate3433(.a(gate2179inter4), .b(gate2179inter3), .O(gate2179inter5));
  nor2  gate3434(.a(gate2179inter5), .b(gate2179inter2), .O(gate2179inter6));
  inv1  gate3435(.a(N5208), .O(gate2179inter7));
  inv1  gate3436(.a(N7872), .O(gate2179inter8));
  nand2 gate3437(.a(gate2179inter8), .b(gate2179inter7), .O(gate2179inter9));
  nand2 gate3438(.a(s_161), .b(gate2179inter3), .O(gate2179inter10));
  nor2  gate3439(.a(gate2179inter10), .b(gate2179inter9), .O(gate2179inter11));
  nor2  gate3440(.a(gate2179inter11), .b(gate2179inter6), .O(gate2179inter12));
  nand2 gate3441(.a(gate2179inter12), .b(gate2179inter1), .O(N7886));
nand2 gate2180( .a(N6356), .b(N7874), .O(N7887) );
nand2 gate2181( .a(N7879), .b(N7861), .O(N7890) );
nand2 gate2182( .a(N7880), .b(N7863), .O(N7893) );
inv1 gate2183( .a(N7864), .O(N7896) );
nand2 gate2184( .a(N7864), .b(N6753), .O(N7897) );
inv1 gate2185( .a(N7867), .O(N7898) );

  xor2  gate3246(.a(N6762), .b(N7867), .O(gate2186inter0));
  nand2 gate3247(.a(gate2186inter0), .b(s_134), .O(gate2186inter1));
  and2  gate3248(.a(N6762), .b(N7867), .O(gate2186inter2));
  inv1  gate3249(.a(s_134), .O(gate2186inter3));
  inv1  gate3250(.a(s_135), .O(gate2186inter4));
  nand2 gate3251(.a(gate2186inter4), .b(gate2186inter3), .O(gate2186inter5));
  nor2  gate3252(.a(gate2186inter5), .b(gate2186inter2), .O(gate2186inter6));
  inv1  gate3253(.a(N7867), .O(gate2186inter7));
  inv1  gate3254(.a(N6762), .O(gate2186inter8));
  nand2 gate3255(.a(gate2186inter8), .b(gate2186inter7), .O(gate2186inter9));
  nand2 gate3256(.a(s_135), .b(gate2186inter3), .O(gate2186inter10));
  nor2  gate3257(.a(gate2186inter10), .b(gate2186inter9), .O(gate2186inter11));
  nor2  gate3258(.a(gate2186inter11), .b(gate2186inter6), .O(gate2186inter12));
  nand2 gate3259(.a(gate2186inter12), .b(gate2186inter1), .O(N7899));

  xor2  gate3344(.a(N7871), .b(N7885), .O(gate2187inter0));
  nand2 gate3345(.a(gate2187inter0), .b(s_148), .O(gate2187inter1));
  and2  gate3346(.a(N7871), .b(N7885), .O(gate2187inter2));
  inv1  gate3347(.a(s_148), .O(gate2187inter3));
  inv1  gate3348(.a(s_149), .O(gate2187inter4));
  nand2 gate3349(.a(gate2187inter4), .b(gate2187inter3), .O(gate2187inter5));
  nor2  gate3350(.a(gate2187inter5), .b(gate2187inter2), .O(gate2187inter6));
  inv1  gate3351(.a(N7885), .O(gate2187inter7));
  inv1  gate3352(.a(N7871), .O(gate2187inter8));
  nand2 gate3353(.a(gate2187inter8), .b(gate2187inter7), .O(gate2187inter9));
  nand2 gate3354(.a(s_149), .b(gate2187inter3), .O(gate2187inter10));
  nor2  gate3355(.a(gate2187inter10), .b(gate2187inter9), .O(gate2187inter11));
  nor2  gate3356(.a(gate2187inter11), .b(gate2187inter6), .O(gate2187inter12));
  nand2 gate3357(.a(gate2187inter12), .b(gate2187inter1), .O(N7900));
nand2 gate2188( .a(N7886), .b(N7873), .O(N7903) );

  xor2  gate3050(.a(N7875), .b(N7887), .O(gate2189inter0));
  nand2 gate3051(.a(gate2189inter0), .b(s_106), .O(gate2189inter1));
  and2  gate3052(.a(N7875), .b(N7887), .O(gate2189inter2));
  inv1  gate3053(.a(s_106), .O(gate2189inter3));
  inv1  gate3054(.a(s_107), .O(gate2189inter4));
  nand2 gate3055(.a(gate2189inter4), .b(gate2189inter3), .O(gate2189inter5));
  nor2  gate3056(.a(gate2189inter5), .b(gate2189inter2), .O(gate2189inter6));
  inv1  gate3057(.a(N7887), .O(gate2189inter7));
  inv1  gate3058(.a(N7875), .O(gate2189inter8));
  nand2 gate3059(.a(gate2189inter8), .b(gate2189inter7), .O(gate2189inter9));
  nand2 gate3060(.a(s_107), .b(gate2189inter3), .O(gate2189inter10));
  nor2  gate3061(.a(gate2189inter10), .b(gate2189inter9), .O(gate2189inter11));
  nor2  gate3062(.a(gate2189inter11), .b(gate2189inter6), .O(gate2189inter12));
  nand2 gate3063(.a(gate2189inter12), .b(gate2189inter1), .O(N7906));
inv1 gate2190( .a(N7876), .O(N7909) );

  xor2  gate3554(.a(N6791), .b(N7876), .O(gate2191inter0));
  nand2 gate3555(.a(gate2191inter0), .b(s_178), .O(gate2191inter1));
  and2  gate3556(.a(N6791), .b(N7876), .O(gate2191inter2));
  inv1  gate3557(.a(s_178), .O(gate2191inter3));
  inv1  gate3558(.a(s_179), .O(gate2191inter4));
  nand2 gate3559(.a(gate2191inter4), .b(gate2191inter3), .O(gate2191inter5));
  nor2  gate3560(.a(gate2191inter5), .b(gate2191inter2), .O(gate2191inter6));
  inv1  gate3561(.a(N7876), .O(gate2191inter7));
  inv1  gate3562(.a(N6791), .O(gate2191inter8));
  nand2 gate3563(.a(gate2191inter8), .b(gate2191inter7), .O(gate2191inter9));
  nand2 gate3564(.a(s_179), .b(gate2191inter3), .O(gate2191inter10));
  nor2  gate3565(.a(gate2191inter10), .b(gate2191inter9), .O(gate2191inter11));
  nor2  gate3566(.a(gate2191inter11), .b(gate2191inter6), .O(gate2191inter12));
  nand2 gate3567(.a(gate2191inter12), .b(gate2191inter1), .O(N7910));

  xor2  gate3484(.a(N7896), .b(N6301), .O(gate2192inter0));
  nand2 gate3485(.a(gate2192inter0), .b(s_168), .O(gate2192inter1));
  and2  gate3486(.a(N7896), .b(N6301), .O(gate2192inter2));
  inv1  gate3487(.a(s_168), .O(gate2192inter3));
  inv1  gate3488(.a(s_169), .O(gate2192inter4));
  nand2 gate3489(.a(gate2192inter4), .b(gate2192inter3), .O(gate2192inter5));
  nor2  gate3490(.a(gate2192inter5), .b(gate2192inter2), .O(gate2192inter6));
  inv1  gate3491(.a(N6301), .O(gate2192inter7));
  inv1  gate3492(.a(N7896), .O(gate2192inter8));
  nand2 gate3493(.a(gate2192inter8), .b(gate2192inter7), .O(gate2192inter9));
  nand2 gate3494(.a(s_169), .b(gate2192inter3), .O(gate2192inter10));
  nor2  gate3495(.a(gate2192inter10), .b(gate2192inter9), .O(gate2192inter11));
  nor2  gate3496(.a(gate2192inter11), .b(gate2192inter6), .O(gate2192inter12));
  nand2 gate3497(.a(gate2192inter12), .b(gate2192inter1), .O(N7917));

  xor2  gate3666(.a(N7898), .b(N6319), .O(gate2193inter0));
  nand2 gate3667(.a(gate2193inter0), .b(s_194), .O(gate2193inter1));
  and2  gate3668(.a(N7898), .b(N6319), .O(gate2193inter2));
  inv1  gate3669(.a(s_194), .O(gate2193inter3));
  inv1  gate3670(.a(s_195), .O(gate2193inter4));
  nand2 gate3671(.a(gate2193inter4), .b(gate2193inter3), .O(gate2193inter5));
  nor2  gate3672(.a(gate2193inter5), .b(gate2193inter2), .O(gate2193inter6));
  inv1  gate3673(.a(N6319), .O(gate2193inter7));
  inv1  gate3674(.a(N7898), .O(gate2193inter8));
  nand2 gate3675(.a(gate2193inter8), .b(gate2193inter7), .O(gate2193inter9));
  nand2 gate3676(.a(s_195), .b(gate2193inter3), .O(gate2193inter10));
  nor2  gate3677(.a(gate2193inter10), .b(gate2193inter9), .O(gate2193inter11));
  nor2  gate3678(.a(gate2193inter11), .b(gate2193inter6), .O(gate2193inter12));
  nand2 gate3679(.a(gate2193inter12), .b(gate2193inter1), .O(N7918));
nand2 gate2194( .a(N6367), .b(N7909), .O(N7923) );
inv1 gate2195( .a(N7890), .O(N7924) );
nand2 gate2196( .a(N7890), .b(N6680), .O(N7925) );
inv1 gate2197( .a(N7893), .O(N7926) );
nand2 gate2198( .a(N7893), .b(N6681), .O(N7927) );
inv1 gate2199( .a(N7900), .O(N7928) );

  xor2  gate2574(.a(N5690), .b(N7900), .O(gate2200inter0));
  nand2 gate2575(.a(gate2200inter0), .b(s_38), .O(gate2200inter1));
  and2  gate2576(.a(N5690), .b(N7900), .O(gate2200inter2));
  inv1  gate2577(.a(s_38), .O(gate2200inter3));
  inv1  gate2578(.a(s_39), .O(gate2200inter4));
  nand2 gate2579(.a(gate2200inter4), .b(gate2200inter3), .O(gate2200inter5));
  nor2  gate2580(.a(gate2200inter5), .b(gate2200inter2), .O(gate2200inter6));
  inv1  gate2581(.a(N7900), .O(gate2200inter7));
  inv1  gate2582(.a(N5690), .O(gate2200inter8));
  nand2 gate2583(.a(gate2200inter8), .b(gate2200inter7), .O(gate2200inter9));
  nand2 gate2584(.a(s_39), .b(gate2200inter3), .O(gate2200inter10));
  nor2  gate2585(.a(gate2200inter10), .b(gate2200inter9), .O(gate2200inter11));
  nor2  gate2586(.a(gate2200inter11), .b(gate2200inter6), .O(gate2200inter12));
  nand2 gate2587(.a(gate2200inter12), .b(gate2200inter1), .O(N7929));
inv1 gate2201( .a(N7903), .O(N7930) );
nand2 gate2202( .a(N7903), .b(N5691), .O(N7931) );

  xor2  gate3778(.a(N7897), .b(N7917), .O(gate2203inter0));
  nand2 gate3779(.a(gate2203inter0), .b(s_210), .O(gate2203inter1));
  and2  gate3780(.a(N7897), .b(N7917), .O(gate2203inter2));
  inv1  gate3781(.a(s_210), .O(gate2203inter3));
  inv1  gate3782(.a(s_211), .O(gate2203inter4));
  nand2 gate3783(.a(gate2203inter4), .b(gate2203inter3), .O(gate2203inter5));
  nor2  gate3784(.a(gate2203inter5), .b(gate2203inter2), .O(gate2203inter6));
  inv1  gate3785(.a(N7917), .O(gate2203inter7));
  inv1  gate3786(.a(N7897), .O(gate2203inter8));
  nand2 gate3787(.a(gate2203inter8), .b(gate2203inter7), .O(gate2203inter9));
  nand2 gate3788(.a(s_211), .b(gate2203inter3), .O(gate2203inter10));
  nor2  gate3789(.a(gate2203inter10), .b(gate2203inter9), .O(gate2203inter11));
  nor2  gate3790(.a(gate2203inter11), .b(gate2203inter6), .O(gate2203inter12));
  nand2 gate3791(.a(gate2203inter12), .b(gate2203inter1), .O(N7932));
nand2 gate2204( .a(N7918), .b(N7899), .O(N7935) );
inv1 gate2205( .a(N7906), .O(N7938) );
nand2 gate2206( .a(N7906), .b(N6784), .O(N7939) );
nand2 gate2207( .a(N7923), .b(N7910), .O(N7940) );
nand2 gate2208( .a(N6280), .b(N7924), .O(N7943) );

  xor2  gate2868(.a(N7926), .b(N6292), .O(gate2209inter0));
  nand2 gate2869(.a(gate2209inter0), .b(s_80), .O(gate2209inter1));
  and2  gate2870(.a(N7926), .b(N6292), .O(gate2209inter2));
  inv1  gate2871(.a(s_80), .O(gate2209inter3));
  inv1  gate2872(.a(s_81), .O(gate2209inter4));
  nand2 gate2873(.a(gate2209inter4), .b(gate2209inter3), .O(gate2209inter5));
  nor2  gate2874(.a(gate2209inter5), .b(gate2209inter2), .O(gate2209inter6));
  inv1  gate2875(.a(N6292), .O(gate2209inter7));
  inv1  gate2876(.a(N7926), .O(gate2209inter8));
  nand2 gate2877(.a(gate2209inter8), .b(gate2209inter7), .O(gate2209inter9));
  nand2 gate2878(.a(s_81), .b(gate2209inter3), .O(gate2209inter10));
  nor2  gate2879(.a(gate2209inter10), .b(gate2209inter9), .O(gate2209inter11));
  nor2  gate2880(.a(gate2209inter11), .b(gate2209inter6), .O(gate2209inter12));
  nand2 gate2881(.a(gate2209inter12), .b(gate2209inter1), .O(N7944));
nand2 gate2210( .a(N5202), .b(N7928), .O(N7945) );
nand2 gate2211( .a(N5211), .b(N7930), .O(N7946) );
nand2 gate2212( .a(N6359), .b(N7938), .O(N7951) );
nand2 gate2213( .a(N7943), .b(N7925), .O(N7954) );
nand2 gate2214( .a(N7944), .b(N7927), .O(N7957) );

  xor2  gate2770(.a(N7929), .b(N7945), .O(gate2215inter0));
  nand2 gate2771(.a(gate2215inter0), .b(s_66), .O(gate2215inter1));
  and2  gate2772(.a(N7929), .b(N7945), .O(gate2215inter2));
  inv1  gate2773(.a(s_66), .O(gate2215inter3));
  inv1  gate2774(.a(s_67), .O(gate2215inter4));
  nand2 gate2775(.a(gate2215inter4), .b(gate2215inter3), .O(gate2215inter5));
  nor2  gate2776(.a(gate2215inter5), .b(gate2215inter2), .O(gate2215inter6));
  inv1  gate2777(.a(N7945), .O(gate2215inter7));
  inv1  gate2778(.a(N7929), .O(gate2215inter8));
  nand2 gate2779(.a(gate2215inter8), .b(gate2215inter7), .O(gate2215inter9));
  nand2 gate2780(.a(s_67), .b(gate2215inter3), .O(gate2215inter10));
  nor2  gate2781(.a(gate2215inter10), .b(gate2215inter9), .O(gate2215inter11));
  nor2  gate2782(.a(gate2215inter11), .b(gate2215inter6), .O(gate2215inter12));
  nand2 gate2783(.a(gate2215inter12), .b(gate2215inter1), .O(N7960));

  xor2  gate2406(.a(N7931), .b(N7946), .O(gate2216inter0));
  nand2 gate2407(.a(gate2216inter0), .b(s_14), .O(gate2216inter1));
  and2  gate2408(.a(N7931), .b(N7946), .O(gate2216inter2));
  inv1  gate2409(.a(s_14), .O(gate2216inter3));
  inv1  gate2410(.a(s_15), .O(gate2216inter4));
  nand2 gate2411(.a(gate2216inter4), .b(gate2216inter3), .O(gate2216inter5));
  nor2  gate2412(.a(gate2216inter5), .b(gate2216inter2), .O(gate2216inter6));
  inv1  gate2413(.a(N7946), .O(gate2216inter7));
  inv1  gate2414(.a(N7931), .O(gate2216inter8));
  nand2 gate2415(.a(gate2216inter8), .b(gate2216inter7), .O(gate2216inter9));
  nand2 gate2416(.a(s_15), .b(gate2216inter3), .O(gate2216inter10));
  nor2  gate2417(.a(gate2216inter10), .b(gate2216inter9), .O(gate2216inter11));
  nor2  gate2418(.a(gate2216inter11), .b(gate2216inter6), .O(gate2216inter12));
  nand2 gate2419(.a(gate2216inter12), .b(gate2216inter1), .O(N7963));
inv1 gate2217( .a(N7932), .O(N7966) );
nand2 gate2218( .a(N7932), .b(N6754), .O(N7967) );
inv1 gate2219( .a(N7935), .O(N7968) );
nand2 gate2220( .a(N7935), .b(N6755), .O(N7969) );
nand2 gate2221( .a(N7951), .b(N7939), .O(N7970) );
inv1 gate2222( .a(N7940), .O(N7973) );

  xor2  gate3330(.a(N6785), .b(N7940), .O(gate2223inter0));
  nand2 gate3331(.a(gate2223inter0), .b(s_146), .O(gate2223inter1));
  and2  gate3332(.a(N6785), .b(N7940), .O(gate2223inter2));
  inv1  gate3333(.a(s_146), .O(gate2223inter3));
  inv1  gate3334(.a(s_147), .O(gate2223inter4));
  nand2 gate3335(.a(gate2223inter4), .b(gate2223inter3), .O(gate2223inter5));
  nor2  gate3336(.a(gate2223inter5), .b(gate2223inter2), .O(gate2223inter6));
  inv1  gate3337(.a(N7940), .O(gate2223inter7));
  inv1  gate3338(.a(N6785), .O(gate2223inter8));
  nand2 gate3339(.a(gate2223inter8), .b(gate2223inter7), .O(gate2223inter9));
  nand2 gate3340(.a(s_147), .b(gate2223inter3), .O(gate2223inter10));
  nor2  gate3341(.a(gate2223inter10), .b(gate2223inter9), .O(gate2223inter11));
  nor2  gate3342(.a(gate2223inter11), .b(gate2223inter6), .O(gate2223inter12));
  nand2 gate3343(.a(gate2223inter12), .b(gate2223inter1), .O(N7974));
nand2 gate2224( .a(N6304), .b(N7966), .O(N7984) );
nand2 gate2225( .a(N6322), .b(N7968), .O(N7985) );

  xor2  gate2448(.a(N7973), .b(N6370), .O(gate2226inter0));
  nand2 gate2449(.a(gate2226inter0), .b(s_20), .O(gate2226inter1));
  and2  gate2450(.a(N7973), .b(N6370), .O(gate2226inter2));
  inv1  gate2451(.a(s_20), .O(gate2226inter3));
  inv1  gate2452(.a(s_21), .O(gate2226inter4));
  nand2 gate2453(.a(gate2226inter4), .b(gate2226inter3), .O(gate2226inter5));
  nor2  gate2454(.a(gate2226inter5), .b(gate2226inter2), .O(gate2226inter6));
  inv1  gate2455(.a(N6370), .O(gate2226inter7));
  inv1  gate2456(.a(N7973), .O(gate2226inter8));
  nand2 gate2457(.a(gate2226inter8), .b(gate2226inter7), .O(gate2226inter9));
  nand2 gate2458(.a(s_21), .b(gate2226inter3), .O(gate2226inter10));
  nor2  gate2459(.a(gate2226inter10), .b(gate2226inter9), .O(gate2226inter11));
  nor2  gate2460(.a(gate2226inter11), .b(gate2226inter6), .O(gate2226inter12));
  nand2 gate2461(.a(gate2226inter12), .b(gate2226inter1), .O(N7987));
and3 gate2227( .a(N7957), .b(N6831), .c(N1157), .O(N7988) );
and3 gate2228( .a(N7954), .b(N6415), .c(N1157), .O(N7989) );
and3 gate2229( .a(N7957), .b(N7041), .c(N566), .O(N7990) );
and3 gate2230( .a(N7954), .b(N7177), .c(N566), .O(N7991) );
inv1 gate2231( .a(N7970), .O(N7992) );
nand2 gate2232( .a(N7970), .b(N6448), .O(N7993) );
and3 gate2233( .a(N7963), .b(N6857), .c(N1219), .O(N7994) );
and3 gate2234( .a(N7960), .b(N6441), .c(N1219), .O(N7995) );
and3 gate2235( .a(N7963), .b(N7065), .c(N583), .O(N7996) );
and3 gate2236( .a(N7960), .b(N7182), .c(N583), .O(N7997) );
nand2 gate2237( .a(N7984), .b(N7967), .O(N7998) );
nand2 gate2238( .a(N7985), .b(N7969), .O(N8001) );
nand2 gate2239( .a(N7987), .b(N7974), .O(N8004) );
nand2 gate2240( .a(N6051), .b(N7992), .O(N8009) );
or4 gate2241( .a(N7988), .b(N7989), .c(N7990), .d(N7991), .O(N8013) );
or4 gate2242( .a(N7994), .b(N7995), .c(N7996), .d(N7997), .O(N8017) );
inv1 gate2243( .a(N7998), .O(N8020) );

  xor2  gate3610(.a(N6682), .b(N7998), .O(gate2244inter0));
  nand2 gate3611(.a(gate2244inter0), .b(s_186), .O(gate2244inter1));
  and2  gate3612(.a(N6682), .b(N7998), .O(gate2244inter2));
  inv1  gate3613(.a(s_186), .O(gate2244inter3));
  inv1  gate3614(.a(s_187), .O(gate2244inter4));
  nand2 gate3615(.a(gate2244inter4), .b(gate2244inter3), .O(gate2244inter5));
  nor2  gate3616(.a(gate2244inter5), .b(gate2244inter2), .O(gate2244inter6));
  inv1  gate3617(.a(N7998), .O(gate2244inter7));
  inv1  gate3618(.a(N6682), .O(gate2244inter8));
  nand2 gate3619(.a(gate2244inter8), .b(gate2244inter7), .O(gate2244inter9));
  nand2 gate3620(.a(s_187), .b(gate2244inter3), .O(gate2244inter10));
  nor2  gate3621(.a(gate2244inter10), .b(gate2244inter9), .O(gate2244inter11));
  nor2  gate3622(.a(gate2244inter11), .b(gate2244inter6), .O(gate2244inter12));
  nand2 gate3623(.a(gate2244inter12), .b(gate2244inter1), .O(N8021));
inv1 gate2245( .a(N8001), .O(N8022) );
nand2 gate2246( .a(N8001), .b(N6683), .O(N8023) );
nand2 gate2247( .a(N8009), .b(N7993), .O(N8025) );
inv1 gate2248( .a(N8004), .O(N8026) );

  xor2  gate2364(.a(N6449), .b(N8004), .O(gate2249inter0));
  nand2 gate2365(.a(gate2249inter0), .b(s_8), .O(gate2249inter1));
  and2  gate2366(.a(N6449), .b(N8004), .O(gate2249inter2));
  inv1  gate2367(.a(s_8), .O(gate2249inter3));
  inv1  gate2368(.a(s_9), .O(gate2249inter4));
  nand2 gate2369(.a(gate2249inter4), .b(gate2249inter3), .O(gate2249inter5));
  nor2  gate2370(.a(gate2249inter5), .b(gate2249inter2), .O(gate2249inter6));
  inv1  gate2371(.a(N8004), .O(gate2249inter7));
  inv1  gate2372(.a(N6449), .O(gate2249inter8));
  nand2 gate2373(.a(gate2249inter8), .b(gate2249inter7), .O(gate2249inter9));
  nand2 gate2374(.a(s_9), .b(gate2249inter3), .O(gate2249inter10));
  nor2  gate2375(.a(gate2249inter10), .b(gate2249inter9), .O(gate2249inter11));
  nor2  gate2376(.a(gate2249inter11), .b(gate2249inter6), .O(gate2249inter12));
  nand2 gate2377(.a(gate2249inter12), .b(gate2249inter1), .O(N8027));
nand2 gate2250( .a(N6307), .b(N8020), .O(N8031) );

  xor2  gate2840(.a(N8022), .b(N6310), .O(gate2251inter0));
  nand2 gate2841(.a(gate2251inter0), .b(s_76), .O(gate2251inter1));
  and2  gate2842(.a(N8022), .b(N6310), .O(gate2251inter2));
  inv1  gate2843(.a(s_76), .O(gate2251inter3));
  inv1  gate2844(.a(s_77), .O(gate2251inter4));
  nand2 gate2845(.a(gate2251inter4), .b(gate2251inter3), .O(gate2251inter5));
  nor2  gate2846(.a(gate2251inter5), .b(gate2251inter2), .O(gate2251inter6));
  inv1  gate2847(.a(N6310), .O(gate2251inter7));
  inv1  gate2848(.a(N8022), .O(gate2251inter8));
  nand2 gate2849(.a(gate2251inter8), .b(gate2251inter7), .O(gate2251inter9));
  nand2 gate2850(.a(s_77), .b(gate2251inter3), .O(gate2251inter10));
  nor2  gate2851(.a(gate2251inter10), .b(gate2251inter9), .O(gate2251inter11));
  nor2  gate2852(.a(gate2251inter11), .b(gate2251inter6), .O(gate2251inter12));
  nand2 gate2853(.a(gate2251inter12), .b(gate2251inter1), .O(N8032));
inv1 gate2252( .a(N8013), .O(N8033) );

  xor2  gate2826(.a(N8026), .b(N6054), .O(gate2253inter0));
  nand2 gate2827(.a(gate2253inter0), .b(s_74), .O(gate2253inter1));
  and2  gate2828(.a(N8026), .b(N6054), .O(gate2253inter2));
  inv1  gate2829(.a(s_74), .O(gate2253inter3));
  inv1  gate2830(.a(s_75), .O(gate2253inter4));
  nand2 gate2831(.a(gate2253inter4), .b(gate2253inter3), .O(gate2253inter5));
  nor2  gate2832(.a(gate2253inter5), .b(gate2253inter2), .O(gate2253inter6));
  inv1  gate2833(.a(N6054), .O(gate2253inter7));
  inv1  gate2834(.a(N8026), .O(gate2253inter8));
  nand2 gate2835(.a(gate2253inter8), .b(gate2253inter7), .O(gate2253inter9));
  nand2 gate2836(.a(s_75), .b(gate2253inter3), .O(gate2253inter10));
  nor2  gate2837(.a(gate2253inter10), .b(gate2253inter9), .O(gate2253inter11));
  nor2  gate2838(.a(gate2253inter11), .b(gate2253inter6), .O(gate2253inter12));
  nand2 gate2839(.a(gate2253inter12), .b(gate2253inter1), .O(N8034));
and2 gate2254( .a(N583), .b(N8025), .O(N8035) );
inv1 gate2255( .a(N8017), .O(N8036) );
nand2 gate2256( .a(N8031), .b(N8021), .O(N8037) );
nand2 gate2257( .a(N8032), .b(N8023), .O(N8038) );
nand2 gate2258( .a(N8034), .b(N8027), .O(N8039) );
inv1 gate2259( .a(N8038), .O(N8040) );
and2 gate2260( .a(N566), .b(N8037), .O(N8041) );
inv1 gate2261( .a(N8039), .O(N8042) );
and2 gate2262( .a(N8040), .b(N1157), .O(N8043) );
and2 gate2263( .a(N8042), .b(N1219), .O(N8044) );
or2 gate2264( .a(N8043), .b(N8041), .O(N8045) );
or2 gate2265( .a(N8044), .b(N8035), .O(N8048) );
nand2 gate2266( .a(N8045), .b(N8033), .O(N8055) );
inv1 gate2267( .a(N8045), .O(N8056) );
nand2 gate2268( .a(N8048), .b(N8036), .O(N8057) );
inv1 gate2269( .a(N8048), .O(N8058) );

  xor2  gate3358(.a(N8056), .b(N8013), .O(gate2270inter0));
  nand2 gate3359(.a(gate2270inter0), .b(s_150), .O(gate2270inter1));
  and2  gate3360(.a(N8056), .b(N8013), .O(gate2270inter2));
  inv1  gate3361(.a(s_150), .O(gate2270inter3));
  inv1  gate3362(.a(s_151), .O(gate2270inter4));
  nand2 gate3363(.a(gate2270inter4), .b(gate2270inter3), .O(gate2270inter5));
  nor2  gate3364(.a(gate2270inter5), .b(gate2270inter2), .O(gate2270inter6));
  inv1  gate3365(.a(N8013), .O(gate2270inter7));
  inv1  gate3366(.a(N8056), .O(gate2270inter8));
  nand2 gate3367(.a(gate2270inter8), .b(gate2270inter7), .O(gate2270inter9));
  nand2 gate3368(.a(s_151), .b(gate2270inter3), .O(gate2270inter10));
  nor2  gate3369(.a(gate2270inter10), .b(gate2270inter9), .O(gate2270inter11));
  nor2  gate3370(.a(gate2270inter11), .b(gate2270inter6), .O(gate2270inter12));
  nand2 gate3371(.a(gate2270inter12), .b(gate2270inter1), .O(N8059));
nand2 gate2271( .a(N8017), .b(N8058), .O(N8060) );
nand2 gate2272( .a(N8055), .b(N8059), .O(N8061) );
nand2 gate2273( .a(N8057), .b(N8060), .O(N8064) );
and3 gate2274( .a(N8064), .b(N1777), .c(N3130), .O(N8071) );
and3 gate2275( .a(N8061), .b(N1761), .c(N3108), .O(N8072) );
inv1 gate2276( .a(N8061), .O(N8073) );
inv1 gate2277( .a(N8064), .O(N8074) );
or4 gate2278( .a(N7526), .b(N8071), .c(N3659), .d(N2625), .O(N8075) );
or4 gate2279( .a(N7636), .b(N8072), .c(N3661), .d(N2627), .O(N8076) );
and2 gate2280( .a(N8073), .b(N1727), .O(N8077) );
and2 gate2281( .a(N8074), .b(N1727), .O(N8078) );
or2 gate2282( .a(N7530), .b(N8077), .O(N8079) );
or2 gate2283( .a(N7479), .b(N8078), .O(N8082) );
and2 gate2284( .a(N8079), .b(N3063), .O(N8089) );
and2 gate2285( .a(N8082), .b(N3063), .O(N8090) );
and2 gate2286( .a(N8079), .b(N3063), .O(N8091) );
and2 gate2287( .a(N8082), .b(N3063), .O(N8092) );
or2 gate2288( .a(N8089), .b(N3071), .O(N8093) );
or2 gate2289( .a(N8090), .b(N3072), .O(N8096) );
or2 gate2290( .a(N8091), .b(N3073), .O(N8099) );
or2 gate2291( .a(N8092), .b(N3074), .O(N8102) );
and3 gate2292( .a(N8102), .b(N2779), .c(N2790), .O(N8113) );
and3 gate2293( .a(N8099), .b(N1327), .c(N2790), .O(N8114) );
and3 gate2294( .a(N8102), .b(N2801), .c(N2812), .O(N8115) );
and3 gate2295( .a(N8099), .b(N1351), .c(N2812), .O(N8116) );
and3 gate2296( .a(N8096), .b(N2681), .c(N2692), .O(N8117) );
and3 gate2297( .a(N8093), .b(N1185), .c(N2692), .O(N8118) );
and3 gate2298( .a(N8096), .b(N2756), .c(N2767), .O(N8119) );
and3 gate2299( .a(N8093), .b(N1247), .c(N2767), .O(N8120) );
or4 gate2300( .a(N8117), .b(N8118), .c(N3662), .d(N2703), .O(N8121) );
or4 gate2301( .a(N8119), .b(N8120), .c(N3663), .d(N2778), .O(N8122) );
or4 gate2302( .a(N8113), .b(N8114), .c(N3650), .d(N2614), .O(N8123) );
or4 gate2303( .a(N8115), .b(N8116), .c(N3658), .d(N2622), .O(N8124) );
and2 gate2304( .a(N8121), .b(N2675), .O(N8125) );
and2 gate2305( .a(N8122), .b(N2750), .O(N8126) );
inv1 gate2306( .a(N8125), .O(N8127) );
inv1 gate2307( .a(N8126), .O(N8128) );

endmodule