module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate380inter0, gate380inter1, gate380inter2, gate380inter3, gate380inter4, gate380inter5, gate380inter6, gate380inter7, gate380inter8, gate380inter9, gate380inter10, gate380inter11, gate380inter12, gate523inter0, gate523inter1, gate523inter2, gate523inter3, gate523inter4, gate523inter5, gate523inter6, gate523inter7, gate523inter8, gate523inter9, gate523inter10, gate523inter11, gate523inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate583inter0, gate583inter1, gate583inter2, gate583inter3, gate583inter4, gate583inter5, gate583inter6, gate583inter7, gate583inter8, gate583inter9, gate583inter10, gate583inter11, gate583inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate824inter0, gate824inter1, gate824inter2, gate824inter3, gate824inter4, gate824inter5, gate824inter6, gate824inter7, gate824inter8, gate824inter9, gate824inter10, gate824inter11, gate824inter12, gate357inter0, gate357inter1, gate357inter2, gate357inter3, gate357inter4, gate357inter5, gate357inter6, gate357inter7, gate357inter8, gate357inter9, gate357inter10, gate357inter11, gate357inter12, gate561inter0, gate561inter1, gate561inter2, gate561inter3, gate561inter4, gate561inter5, gate561inter6, gate561inter7, gate561inter8, gate561inter9, gate561inter10, gate561inter11, gate561inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate542inter0, gate542inter1, gate542inter2, gate542inter3, gate542inter4, gate542inter5, gate542inter6, gate542inter7, gate542inter8, gate542inter9, gate542inter10, gate542inter11, gate542inter12, gate797inter0, gate797inter1, gate797inter2, gate797inter3, gate797inter4, gate797inter5, gate797inter6, gate797inter7, gate797inter8, gate797inter9, gate797inter10, gate797inter11, gate797inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate650inter0, gate650inter1, gate650inter2, gate650inter3, gate650inter4, gate650inter5, gate650inter6, gate650inter7, gate650inter8, gate650inter9, gate650inter10, gate650inter11, gate650inter12, gate303inter0, gate303inter1, gate303inter2, gate303inter3, gate303inter4, gate303inter5, gate303inter6, gate303inter7, gate303inter8, gate303inter9, gate303inter10, gate303inter11, gate303inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate864inter0, gate864inter1, gate864inter2, gate864inter3, gate864inter4, gate864inter5, gate864inter6, gate864inter7, gate864inter8, gate864inter9, gate864inter10, gate864inter11, gate864inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate649inter0, gate649inter1, gate649inter2, gate649inter3, gate649inter4, gate649inter5, gate649inter6, gate649inter7, gate649inter8, gate649inter9, gate649inter10, gate649inter11, gate649inter12, gate608inter0, gate608inter1, gate608inter2, gate608inter3, gate608inter4, gate608inter5, gate608inter6, gate608inter7, gate608inter8, gate608inter9, gate608inter10, gate608inter11, gate608inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate835inter0, gate835inter1, gate835inter2, gate835inter3, gate835inter4, gate835inter5, gate835inter6, gate835inter7, gate835inter8, gate835inter9, gate835inter10, gate835inter11, gate835inter12, gate808inter0, gate808inter1, gate808inter2, gate808inter3, gate808inter4, gate808inter5, gate808inter6, gate808inter7, gate808inter8, gate808inter9, gate808inter10, gate808inter11, gate808inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate315inter0, gate315inter1, gate315inter2, gate315inter3, gate315inter4, gate315inter5, gate315inter6, gate315inter7, gate315inter8, gate315inter9, gate315inter10, gate315inter11, gate315inter12, gate605inter0, gate605inter1, gate605inter2, gate605inter3, gate605inter4, gate605inter5, gate605inter6, gate605inter7, gate605inter8, gate605inter9, gate605inter10, gate605inter11, gate605inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate679inter0, gate679inter1, gate679inter2, gate679inter3, gate679inter4, gate679inter5, gate679inter6, gate679inter7, gate679inter8, gate679inter9, gate679inter10, gate679inter11, gate679inter12, gate319inter0, gate319inter1, gate319inter2, gate319inter3, gate319inter4, gate319inter5, gate319inter6, gate319inter7, gate319inter8, gate319inter9, gate319inter10, gate319inter11, gate319inter12, gate682inter0, gate682inter1, gate682inter2, gate682inter3, gate682inter4, gate682inter5, gate682inter6, gate682inter7, gate682inter8, gate682inter9, gate682inter10, gate682inter11, gate682inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate537inter0, gate537inter1, gate537inter2, gate537inter3, gate537inter4, gate537inter5, gate537inter6, gate537inter7, gate537inter8, gate537inter9, gate537inter10, gate537inter11, gate537inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate636inter0, gate636inter1, gate636inter2, gate636inter3, gate636inter4, gate636inter5, gate636inter6, gate636inter7, gate636inter8, gate636inter9, gate636inter10, gate636inter11, gate636inter12, gate850inter0, gate850inter1, gate850inter2, gate850inter3, gate850inter4, gate850inter5, gate850inter6, gate850inter7, gate850inter8, gate850inter9, gate850inter10, gate850inter11, gate850inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate623inter0, gate623inter1, gate623inter2, gate623inter3, gate623inter4, gate623inter5, gate623inter6, gate623inter7, gate623inter8, gate623inter9, gate623inter10, gate623inter11, gate623inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate681inter0, gate681inter1, gate681inter2, gate681inter3, gate681inter4, gate681inter5, gate681inter6, gate681inter7, gate681inter8, gate681inter9, gate681inter10, gate681inter11, gate681inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate304inter0, gate304inter1, gate304inter2, gate304inter3, gate304inter4, gate304inter5, gate304inter6, gate304inter7, gate304inter8, gate304inter9, gate304inter10, gate304inter11, gate304inter12, gate363inter0, gate363inter1, gate363inter2, gate363inter3, gate363inter4, gate363inter5, gate363inter6, gate363inter7, gate363inter8, gate363inter9, gate363inter10, gate363inter11, gate363inter12, gate798inter0, gate798inter1, gate798inter2, gate798inter3, gate798inter4, gate798inter5, gate798inter6, gate798inter7, gate798inter8, gate798inter9, gate798inter10, gate798inter11, gate798inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate760inter0, gate760inter1, gate760inter2, gate760inter3, gate760inter4, gate760inter5, gate760inter6, gate760inter7, gate760inter8, gate760inter9, gate760inter10, gate760inter11, gate760inter12, gate822inter0, gate822inter1, gate822inter2, gate822inter3, gate822inter4, gate822inter5, gate822inter6, gate822inter7, gate822inter8, gate822inter9, gate822inter10, gate822inter11, gate822inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate837inter0, gate837inter1, gate837inter2, gate837inter3, gate837inter4, gate837inter5, gate837inter6, gate837inter7, gate837inter8, gate837inter9, gate837inter10, gate837inter11, gate837inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate820inter0, gate820inter1, gate820inter2, gate820inter3, gate820inter4, gate820inter5, gate820inter6, gate820inter7, gate820inter8, gate820inter9, gate820inter10, gate820inter11, gate820inter12, gate683inter0, gate683inter1, gate683inter2, gate683inter3, gate683inter4, gate683inter5, gate683inter6, gate683inter7, gate683inter8, gate683inter9, gate683inter10, gate683inter11, gate683inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12;



inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );

  xor2  gate1847(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate1848(.a(gate77inter0), .b(s_138), .O(gate77inter1));
  and2  gate1849(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate1850(.a(s_138), .O(gate77inter3));
  inv1  gate1851(.a(s_139), .O(gate77inter4));
  nand2 gate1852(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1853(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1854(.a(N306), .O(gate77inter7));
  inv1  gate1855(.a(N331), .O(gate77inter8));
  nand2 gate1856(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1857(.a(s_139), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1858(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1859(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1860(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );

  xor2  gate1007(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate1008(.a(gate99inter0), .b(s_18), .O(gate99inter1));
  and2  gate1009(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate1010(.a(s_18), .O(gate99inter3));
  inv1  gate1011(.a(s_19), .O(gate99inter4));
  nand2 gate1012(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1013(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1014(.a(N260), .O(gate99inter7));
  inv1  gate1015(.a(N300), .O(gate99inter8));
  nand2 gate1016(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1017(.a(s_19), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1018(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1019(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1020(.a(gate99inter12), .b(gate99inter1), .O(N608));

  xor2  gate1595(.a(N300), .b(N256), .O(gate100inter0));
  nand2 gate1596(.a(gate100inter0), .b(s_102), .O(gate100inter1));
  and2  gate1597(.a(N300), .b(N256), .O(gate100inter2));
  inv1  gate1598(.a(s_102), .O(gate100inter3));
  inv1  gate1599(.a(s_103), .O(gate100inter4));
  nand2 gate1600(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1601(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1602(.a(N256), .O(gate100inter7));
  inv1  gate1603(.a(N300), .O(gate100inter8));
  nand2 gate1604(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1605(.a(s_103), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1606(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1607(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1608(.a(gate100inter12), .b(gate100inter1), .O(N612));
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );

  xor2  gate1273(.a(N889), .b(N616), .O(gate234inter0));
  nand2 gate1274(.a(gate234inter0), .b(s_56), .O(gate234inter1));
  and2  gate1275(.a(N889), .b(N616), .O(gate234inter2));
  inv1  gate1276(.a(s_56), .O(gate234inter3));
  inv1  gate1277(.a(s_57), .O(gate234inter4));
  nand2 gate1278(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1279(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1280(.a(N616), .O(gate234inter7));
  inv1  gate1281(.a(N889), .O(gate234inter8));
  nand2 gate1282(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1283(.a(s_57), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1284(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1285(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1286(.a(gate234inter12), .b(gate234inter1), .O(N1055));
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );

  xor2  gate1567(.a(N895), .b(N655), .O(gate237inter0));
  nand2 gate1568(.a(gate237inter0), .b(s_98), .O(gate237inter1));
  and2  gate1569(.a(N895), .b(N655), .O(gate237inter2));
  inv1  gate1570(.a(s_98), .O(gate237inter3));
  inv1  gate1571(.a(s_99), .O(gate237inter4));
  nand2 gate1572(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1573(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1574(.a(N655), .O(gate237inter7));
  inv1  gate1575(.a(N895), .O(gate237inter8));
  nand2 gate1576(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1577(.a(s_99), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1578(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1579(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1580(.a(gate237inter12), .b(gate237inter1), .O(N1067));

  xor2  gate951(.a(N896), .b(N652), .O(gate238inter0));
  nand2 gate952(.a(gate238inter0), .b(s_10), .O(gate238inter1));
  and2  gate953(.a(N896), .b(N652), .O(gate238inter2));
  inv1  gate954(.a(s_10), .O(gate238inter3));
  inv1  gate955(.a(s_11), .O(gate238inter4));
  nand2 gate956(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate957(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate958(.a(N652), .O(gate238inter7));
  inv1  gate959(.a(N896), .O(gate238inter8));
  nand2 gate960(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate961(.a(s_11), .b(gate238inter3), .O(gate238inter10));
  nor2  gate962(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate963(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate964(.a(gate238inter12), .b(gate238inter1), .O(N1068));
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );

  xor2  gate1931(.a(N991), .b(N727), .O(gate241inter0));
  nand2 gate1932(.a(gate241inter0), .b(s_150), .O(gate241inter1));
  and2  gate1933(.a(N991), .b(N727), .O(gate241inter2));
  inv1  gate1934(.a(s_150), .O(gate241inter3));
  inv1  gate1935(.a(s_151), .O(gate241inter4));
  nand2 gate1936(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1937(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1938(.a(N727), .O(gate241inter7));
  inv1  gate1939(.a(N991), .O(gate241inter8));
  nand2 gate1940(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1941(.a(s_151), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1942(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1943(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1944(.a(gate241inter12), .b(gate241inter1), .O(N1121));
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );

  xor2  gate1497(.a(N1055), .b(N1054), .O(gate251inter0));
  nand2 gate1498(.a(gate251inter0), .b(s_88), .O(gate251inter1));
  and2  gate1499(.a(N1055), .b(N1054), .O(gate251inter2));
  inv1  gate1500(.a(s_88), .O(gate251inter3));
  inv1  gate1501(.a(s_89), .O(gate251inter4));
  nand2 gate1502(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1503(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1504(.a(N1054), .O(gate251inter7));
  inv1  gate1505(.a(N1055), .O(gate251inter8));
  nand2 gate1506(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1507(.a(s_89), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1508(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1509(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1510(.a(gate251inter12), .b(gate251inter1), .O(N1150));
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );

  xor2  gate1889(.a(N1068), .b(N1067), .O(gate263inter0));
  nand2 gate1890(.a(gate263inter0), .b(s_144), .O(gate263inter1));
  and2  gate1891(.a(N1068), .b(N1067), .O(gate263inter2));
  inv1  gate1892(.a(s_144), .O(gate263inter3));
  inv1  gate1893(.a(s_145), .O(gate263inter4));
  nand2 gate1894(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1895(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1896(.a(N1067), .O(gate263inter7));
  inv1  gate1897(.a(N1068), .O(gate263inter8));
  nand2 gate1898(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1899(.a(s_145), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1900(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1901(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1902(.a(gate263inter12), .b(gate263inter1), .O(N1162));
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate1147(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate1148(.a(gate275inter0), .b(s_38), .O(gate275inter1));
  and2  gate1149(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate1150(.a(s_38), .O(gate275inter3));
  inv1  gate1151(.a(s_39), .O(gate275inter4));
  nand2 gate1152(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1153(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1154(.a(N1016), .O(gate275inter7));
  inv1  gate1155(.a(N946), .O(gate275inter8));
  nand2 gate1156(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1157(.a(s_39), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1158(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1159(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1160(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );

  xor2  gate1385(.a(N958), .b(N1025), .O(gate281inter0));
  nand2 gate1386(.a(gate281inter0), .b(s_72), .O(gate281inter1));
  and2  gate1387(.a(N958), .b(N1025), .O(gate281inter2));
  inv1  gate1388(.a(s_72), .O(gate281inter3));
  inv1  gate1389(.a(s_73), .O(gate281inter4));
  nand2 gate1390(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1391(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1392(.a(N1025), .O(gate281inter7));
  inv1  gate1393(.a(N958), .O(gate281inter8));
  nand2 gate1394(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1395(.a(s_73), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1396(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1397(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1398(.a(gate281inter12), .b(gate281inter1), .O(N1216));
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );

  xor2  gate1441(.a(N984), .b(N981), .O(gate296inter0));
  nand2 gate1442(.a(gate296inter0), .b(s_80), .O(gate296inter1));
  and2  gate1443(.a(N984), .b(N981), .O(gate296inter2));
  inv1  gate1444(.a(s_80), .O(gate296inter3));
  inv1  gate1445(.a(s_81), .O(gate296inter4));
  nand2 gate1446(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1447(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1448(.a(N981), .O(gate296inter7));
  inv1  gate1449(.a(N984), .O(gate296inter8));
  nand2 gate1450(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1451(.a(s_81), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1452(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1453(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1454(.a(gate296inter12), .b(gate296inter1), .O(N1231));

  xor2  gate965(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate966(.a(gate297inter0), .b(s_12), .O(gate297inter1));
  and2  gate967(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate968(.a(s_12), .O(gate297inter3));
  inv1  gate969(.a(s_13), .O(gate297inter4));
  nand2 gate970(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate971(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate972(.a(N1119), .O(gate297inter7));
  inv1  gate973(.a(N1120), .O(gate297inter8));
  nand2 gate974(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate975(.a(s_13), .b(gate297inter3), .O(gate297inter10));
  nor2  gate976(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate977(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate978(.a(gate297inter12), .b(gate297inter1), .O(N1232));

  xor2  gate1399(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate1400(.a(gate298inter0), .b(s_74), .O(gate298inter1));
  and2  gate1401(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate1402(.a(s_74), .O(gate298inter3));
  inv1  gate1403(.a(s_75), .O(gate298inter4));
  nand2 gate1404(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate1405(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate1406(.a(N1121), .O(gate298inter7));
  inv1  gate1407(.a(N1122), .O(gate298inter8));
  nand2 gate1408(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate1409(.a(s_75), .b(gate298inter3), .O(gate298inter10));
  nor2  gate1410(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate1411(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate1412(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );

  xor2  gate1217(.a(N1001), .b(N1049), .O(gate303inter0));
  nand2 gate1218(.a(gate303inter0), .b(s_48), .O(gate303inter1));
  and2  gate1219(.a(N1001), .b(N1049), .O(gate303inter2));
  inv1  gate1220(.a(s_48), .O(gate303inter3));
  inv1  gate1221(.a(s_49), .O(gate303inter4));
  nand2 gate1222(.a(gate303inter4), .b(gate303inter3), .O(gate303inter5));
  nor2  gate1223(.a(gate303inter5), .b(gate303inter2), .O(gate303inter6));
  inv1  gate1224(.a(N1049), .O(gate303inter7));
  inv1  gate1225(.a(N1001), .O(gate303inter8));
  nand2 gate1226(.a(gate303inter8), .b(gate303inter7), .O(gate303inter9));
  nand2 gate1227(.a(s_49), .b(gate303inter3), .O(gate303inter10));
  nor2  gate1228(.a(gate303inter10), .b(gate303inter9), .O(gate303inter11));
  nor2  gate1229(.a(gate303inter11), .b(gate303inter6), .O(gate303inter12));
  nand2 gate1230(.a(gate303inter12), .b(gate303inter1), .O(N1242));

  xor2  gate1805(.a(N1129), .b(N1128), .O(gate304inter0));
  nand2 gate1806(.a(gate304inter0), .b(s_132), .O(gate304inter1));
  and2  gate1807(.a(N1129), .b(N1128), .O(gate304inter2));
  inv1  gate1808(.a(s_132), .O(gate304inter3));
  inv1  gate1809(.a(s_133), .O(gate304inter4));
  nand2 gate1810(.a(gate304inter4), .b(gate304inter3), .O(gate304inter5));
  nor2  gate1811(.a(gate304inter5), .b(gate304inter2), .O(gate304inter6));
  inv1  gate1812(.a(N1128), .O(gate304inter7));
  inv1  gate1813(.a(N1129), .O(gate304inter8));
  nand2 gate1814(.a(gate304inter8), .b(gate304inter7), .O(gate304inter9));
  nand2 gate1815(.a(s_133), .b(gate304inter3), .O(gate304inter10));
  nor2  gate1816(.a(gate304inter10), .b(gate304inter9), .O(gate304inter11));
  nor2  gate1817(.a(gate304inter11), .b(gate304inter6), .O(gate304inter12));
  nand2 gate1818(.a(gate304inter12), .b(gate304inter1), .O(N1243));
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );

  xor2  gate1469(.a(N1209), .b(N694), .O(gate315inter0));
  nand2 gate1470(.a(gate315inter0), .b(s_84), .O(gate315inter1));
  and2  gate1471(.a(N1209), .b(N694), .O(gate315inter2));
  inv1  gate1472(.a(s_84), .O(gate315inter3));
  inv1  gate1473(.a(s_85), .O(gate315inter4));
  nand2 gate1474(.a(gate315inter4), .b(gate315inter3), .O(gate315inter5));
  nor2  gate1475(.a(gate315inter5), .b(gate315inter2), .O(gate315inter6));
  inv1  gate1476(.a(N694), .O(gate315inter7));
  inv1  gate1477(.a(N1209), .O(gate315inter8));
  nand2 gate1478(.a(gate315inter8), .b(gate315inter7), .O(gate315inter9));
  nand2 gate1479(.a(s_85), .b(gate315inter3), .O(gate315inter10));
  nor2  gate1480(.a(gate315inter10), .b(gate315inter9), .O(gate315inter11));
  nor2  gate1481(.a(gate315inter11), .b(gate315inter6), .O(gate315inter12));
  nand2 gate1482(.a(gate315inter12), .b(gate315inter1), .O(N1311));
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );

  xor2  gate1539(.a(N1220), .b(N706), .O(gate319inter0));
  nand2 gate1540(.a(gate319inter0), .b(s_94), .O(gate319inter1));
  and2  gate1541(.a(N1220), .b(N706), .O(gate319inter2));
  inv1  gate1542(.a(s_94), .O(gate319inter3));
  inv1  gate1543(.a(s_95), .O(gate319inter4));
  nand2 gate1544(.a(gate319inter4), .b(gate319inter3), .O(gate319inter5));
  nor2  gate1545(.a(gate319inter5), .b(gate319inter2), .O(gate319inter6));
  inv1  gate1546(.a(N706), .O(gate319inter7));
  inv1  gate1547(.a(N1220), .O(gate319inter8));
  nand2 gate1548(.a(gate319inter8), .b(gate319inter7), .O(gate319inter9));
  nand2 gate1549(.a(s_95), .b(gate319inter3), .O(gate319inter10));
  nor2  gate1550(.a(gate319inter10), .b(gate319inter9), .O(gate319inter11));
  nor2  gate1551(.a(gate319inter11), .b(gate319inter6), .O(gate319inter12));
  nand2 gate1552(.a(gate319inter12), .b(gate319inter1), .O(N1315));
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );

  xor2  gate1091(.a(N1160), .b(N1267), .O(gate328inter0));
  nand2 gate1092(.a(gate328inter0), .b(s_30), .O(gate328inter1));
  and2  gate1093(.a(N1160), .b(N1267), .O(gate328inter2));
  inv1  gate1094(.a(s_30), .O(gate328inter3));
  inv1  gate1095(.a(s_31), .O(gate328inter4));
  nand2 gate1096(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate1097(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate1098(.a(N1267), .O(gate328inter7));
  inv1  gate1099(.a(N1160), .O(gate328inter8));
  nand2 gate1100(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate1101(.a(s_31), .b(gate328inter3), .O(gate328inter10));
  nor2  gate1102(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate1103(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate1104(.a(gate328inter12), .b(gate328inter1), .O(N1344));
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate1189(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate1190(.a(gate347inter0), .b(s_44), .O(gate347inter1));
  and2  gate1191(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate1192(.a(s_44), .O(gate347inter3));
  inv1  gate1193(.a(s_45), .O(gate347inter4));
  nand2 gate1194(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate1195(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate1196(.a(N1232), .O(gate347inter7));
  inv1  gate1197(.a(N990), .O(gate347inter8));
  nand2 gate1198(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate1199(.a(s_45), .b(gate347inter3), .O(gate347inter10));
  nor2  gate1200(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate1201(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate1202(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );

  xor2  gate1119(.a(N1346), .b(N649), .O(gate357inter0));
  nand2 gate1120(.a(gate357inter0), .b(s_34), .O(gate357inter1));
  and2  gate1121(.a(N1346), .b(N649), .O(gate357inter2));
  inv1  gate1122(.a(s_34), .O(gate357inter3));
  inv1  gate1123(.a(s_35), .O(gate357inter4));
  nand2 gate1124(.a(gate357inter4), .b(gate357inter3), .O(gate357inter5));
  nor2  gate1125(.a(gate357inter5), .b(gate357inter2), .O(gate357inter6));
  inv1  gate1126(.a(N649), .O(gate357inter7));
  inv1  gate1127(.a(N1346), .O(gate357inter8));
  nand2 gate1128(.a(gate357inter8), .b(gate357inter7), .O(gate357inter9));
  nand2 gate1129(.a(s_35), .b(gate357inter3), .O(gate357inter10));
  nor2  gate1130(.a(gate357inter10), .b(gate357inter9), .O(gate357inter11));
  nor2  gate1131(.a(gate357inter11), .b(gate357inter6), .O(gate357inter12));
  nand2 gate1132(.a(gate357inter12), .b(gate357inter1), .O(N1412));
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );

  xor2  gate1819(.a(N1396), .b(N640), .O(gate363inter0));
  nand2 gate1820(.a(gate363inter0), .b(s_134), .O(gate363inter1));
  and2  gate1821(.a(N1396), .b(N640), .O(gate363inter2));
  inv1  gate1822(.a(s_134), .O(gate363inter3));
  inv1  gate1823(.a(s_135), .O(gate363inter4));
  nand2 gate1824(.a(gate363inter4), .b(gate363inter3), .O(gate363inter5));
  nor2  gate1825(.a(gate363inter5), .b(gate363inter2), .O(gate363inter6));
  inv1  gate1826(.a(N640), .O(gate363inter7));
  inv1  gate1827(.a(N1396), .O(gate363inter8));
  nand2 gate1828(.a(gate363inter8), .b(gate363inter7), .O(gate363inter9));
  nand2 gate1829(.a(s_135), .b(gate363inter3), .O(gate363inter10));
  nor2  gate1830(.a(gate363inter10), .b(gate363inter9), .O(gate363inter11));
  nor2  gate1831(.a(gate363inter11), .b(gate363inter6), .O(gate363inter12));
  nand2 gate1832(.a(gate363inter12), .b(gate363inter1), .O(N1438));
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );

  xor2  gate881(.a(N1157), .b(N1379), .O(gate380inter0));
  nand2 gate882(.a(gate380inter0), .b(s_0), .O(gate380inter1));
  and2  gate883(.a(N1157), .b(N1379), .O(gate380inter2));
  inv1  gate884(.a(s_0), .O(gate380inter3));
  inv1  gate885(.a(s_1), .O(gate380inter4));
  nand2 gate886(.a(gate380inter4), .b(gate380inter3), .O(gate380inter5));
  nor2  gate887(.a(gate380inter5), .b(gate380inter2), .O(gate380inter6));
  inv1  gate888(.a(N1379), .O(gate380inter7));
  inv1  gate889(.a(N1157), .O(gate380inter8));
  nand2 gate890(.a(gate380inter8), .b(gate380inter7), .O(gate380inter9));
  nand2 gate891(.a(s_1), .b(gate380inter3), .O(gate380inter10));
  nor2  gate892(.a(gate380inter10), .b(gate380inter9), .O(gate380inter11));
  nor2  gate893(.a(gate380inter11), .b(gate380inter6), .O(gate380inter12));
  nand2 gate894(.a(gate380inter12), .b(gate380inter1), .O(N1459));
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );

  xor2  gate1231(.a(N1438), .b(N1397), .O(gate395inter0));
  nand2 gate1232(.a(gate395inter0), .b(s_50), .O(gate395inter1));
  and2  gate1233(.a(N1438), .b(N1397), .O(gate395inter2));
  inv1  gate1234(.a(s_50), .O(gate395inter3));
  inv1  gate1235(.a(s_51), .O(gate395inter4));
  nand2 gate1236(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1237(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1238(.a(N1397), .O(gate395inter7));
  inv1  gate1239(.a(N1438), .O(gate395inter8));
  nand2 gate1240(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1241(.a(s_51), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1242(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1243(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1244(.a(gate395inter12), .b(gate395inter1), .O(N1484));
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );

  xor2  gate1721(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate1722(.a(gate402inter0), .b(s_120), .O(gate402inter1));
  and2  gate1723(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate1724(.a(s_120), .O(gate402inter3));
  inv1  gate1725(.a(s_121), .O(gate402inter4));
  nand2 gate1726(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1727(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1728(.a(N955), .O(gate402inter7));
  inv1  gate1729(.a(N1454), .O(gate402inter8));
  nand2 gate1730(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1731(.a(s_121), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1732(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1733(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1734(.a(gate402inter12), .b(gate402inter1), .O(N1493));
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );

  xor2  gate1035(.a(N1458), .b(N969), .O(gate404inter0));
  nand2 gate1036(.a(gate404inter0), .b(s_22), .O(gate404inter1));
  and2  gate1037(.a(N1458), .b(N969), .O(gate404inter2));
  inv1  gate1038(.a(s_22), .O(gate404inter3));
  inv1  gate1039(.a(s_23), .O(gate404inter4));
  nand2 gate1040(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1041(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1042(.a(N969), .O(gate404inter7));
  inv1  gate1043(.a(N1458), .O(gate404inter8));
  nand2 gate1044(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1045(.a(s_23), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1046(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1047(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1048(.a(gate404inter12), .b(gate404inter1), .O(N1495));
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );

  xor2  gate1287(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate1288(.a(gate406inter0), .b(s_58), .O(gate406inter1));
  and2  gate1289(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate1290(.a(s_58), .O(gate406inter3));
  inv1  gate1291(.a(s_59), .O(gate406inter4));
  nand2 gate1292(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1293(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1294(.a(N998), .O(gate406inter7));
  inv1  gate1295(.a(N1463), .O(gate406inter8));
  nand2 gate1296(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1297(.a(s_59), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1298(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1299(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1300(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );

  xor2  gate1791(.a(N1470), .b(N973), .O(gate409inter0));
  nand2 gate1792(.a(gate409inter0), .b(s_130), .O(gate409inter1));
  and2  gate1793(.a(N1470), .b(N973), .O(gate409inter2));
  inv1  gate1794(.a(s_130), .O(gate409inter3));
  inv1  gate1795(.a(s_131), .O(gate409inter4));
  nand2 gate1796(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1797(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1798(.a(N973), .O(gate409inter7));
  inv1  gate1799(.a(N1470), .O(gate409inter8));
  nand2 gate1800(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1801(.a(s_131), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1802(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1803(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1804(.a(gate409inter12), .b(gate409inter1), .O(N1501));
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );

  xor2  gate1245(.a(N1487), .b(N1443), .O(gate412inter0));
  nand2 gate1246(.a(gate412inter0), .b(s_52), .O(gate412inter1));
  and2  gate1247(.a(N1487), .b(N1443), .O(gate412inter2));
  inv1  gate1248(.a(s_52), .O(gate412inter3));
  inv1  gate1249(.a(s_53), .O(gate412inter4));
  nand2 gate1250(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1251(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1252(.a(N1443), .O(gate412inter7));
  inv1  gate1253(.a(N1487), .O(gate412inter8));
  nand2 gate1254(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1255(.a(s_53), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1256(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1257(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1258(.a(gate412inter12), .b(gate412inter1), .O(N1513));
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );

  xor2  gate1679(.a(N1495), .b(N1457), .O(gate418inter0));
  nand2 gate1680(.a(gate418inter0), .b(s_114), .O(gate418inter1));
  and2  gate1681(.a(N1495), .b(N1457), .O(gate418inter2));
  inv1  gate1682(.a(s_114), .O(gate418inter3));
  inv1  gate1683(.a(s_115), .O(gate418inter4));
  nand2 gate1684(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1685(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1686(.a(N1457), .O(gate418inter7));
  inv1  gate1687(.a(N1495), .O(gate418inter8));
  nand2 gate1688(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1689(.a(s_115), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1690(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1691(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1692(.a(gate418inter12), .b(gate418inter1), .O(N1526));
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate1735(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate1736(.a(gate421inter0), .b(s_122), .O(gate421inter1));
  and2  gate1737(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate1738(.a(s_122), .O(gate421inter3));
  inv1  gate1739(.a(s_123), .O(gate421inter4));
  nand2 gate1740(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1741(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1742(.a(N1462), .O(gate421inter7));
  inv1  gate1743(.a(N1498), .O(gate421inter8));
  nand2 gate1744(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1745(.a(s_123), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1746(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1747(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1748(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );

  xor2  gate1049(.a(N1504), .b(N1476), .O(gate427inter0));
  nand2 gate1050(.a(gate427inter0), .b(s_24), .O(gate427inter1));
  and2  gate1051(.a(N1504), .b(N1476), .O(gate427inter2));
  inv1  gate1052(.a(s_24), .O(gate427inter3));
  inv1  gate1053(.a(s_25), .O(gate427inter4));
  nand2 gate1054(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1055(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1056(.a(N1476), .O(gate427inter7));
  inv1  gate1057(.a(N1504), .O(gate427inter8));
  nand2 gate1058(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1059(.a(s_25), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1060(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1061(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1062(.a(gate427inter12), .b(gate427inter1), .O(N1540));
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );

  xor2  gate909(.a(N1531), .b(N1484), .O(gate432inter0));
  nand2 gate910(.a(gate432inter0), .b(s_4), .O(gate432inter1));
  and2  gate911(.a(N1531), .b(N1484), .O(gate432inter2));
  inv1  gate912(.a(s_4), .O(gate432inter3));
  inv1  gate913(.a(s_5), .O(gate432inter4));
  nand2 gate914(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate915(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate916(.a(N1484), .O(gate432inter7));
  inv1  gate917(.a(N1531), .O(gate432inter8));
  nand2 gate918(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate919(.a(s_5), .b(gate432inter3), .O(gate432inter10));
  nor2  gate920(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate921(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate922(.a(gate432inter12), .b(gate432inter1), .O(N1567));
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );

  xor2  gate1651(.a(N1595), .b(N1478), .O(gate452inter0));
  nand2 gate1652(.a(gate452inter0), .b(s_110), .O(gate452inter1));
  and2  gate1653(.a(N1595), .b(N1478), .O(gate452inter2));
  inv1  gate1654(.a(s_110), .O(gate452inter3));
  inv1  gate1655(.a(s_111), .O(gate452inter4));
  nand2 gate1656(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1657(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1658(.a(N1478), .O(gate452inter7));
  inv1  gate1659(.a(N1595), .O(gate452inter8));
  nand2 gate1660(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1661(.a(s_111), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1662(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1663(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1664(.a(gate452inter12), .b(gate452inter1), .O(N1636));
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );

  xor2  gate1259(.a(N893), .b(N1596), .O(gate462inter0));
  nand2 gate1260(.a(gate462inter0), .b(s_54), .O(gate462inter1));
  and2  gate1261(.a(N893), .b(N1596), .O(gate462inter2));
  inv1  gate1262(.a(s_54), .O(gate462inter3));
  inv1  gate1263(.a(s_55), .O(gate462inter4));
  nand2 gate1264(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1265(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1266(.a(N1596), .O(gate462inter7));
  inv1  gate1267(.a(N893), .O(gate462inter8));
  nand2 gate1268(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1269(.a(s_55), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1270(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1271(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1272(.a(gate462inter12), .b(gate462inter1), .O(N1671));
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );

  xor2  gate1329(.a(N1217), .b(N1606), .O(gate466inter0));
  nand2 gate1330(.a(gate466inter0), .b(s_64), .O(gate466inter1));
  and2  gate1331(.a(N1217), .b(N1606), .O(gate466inter2));
  inv1  gate1332(.a(s_64), .O(gate466inter3));
  inv1  gate1333(.a(s_65), .O(gate466inter4));
  nand2 gate1334(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1335(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1336(.a(N1606), .O(gate466inter7));
  inv1  gate1337(.a(N1217), .O(gate466inter8));
  nand2 gate1338(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1339(.a(s_65), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1340(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1341(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1342(.a(gate466inter12), .b(gate466inter1), .O(N1678));
inv1 gate467( .a(N1606), .O(N1679) );

  xor2  gate1063(.a(N1219), .b(N1609), .O(gate468inter0));
  nand2 gate1064(.a(gate468inter0), .b(s_26), .O(gate468inter1));
  and2  gate1065(.a(N1219), .b(N1609), .O(gate468inter2));
  inv1  gate1066(.a(s_26), .O(gate468inter3));
  inv1  gate1067(.a(s_27), .O(gate468inter4));
  nand2 gate1068(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1069(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1070(.a(N1609), .O(gate468inter7));
  inv1  gate1071(.a(N1219), .O(gate468inter8));
  nand2 gate1072(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1073(.a(s_27), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1074(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1075(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1076(.a(gate468inter12), .b(gate468inter1), .O(N1680));
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );

  xor2  gate1077(.a(N1636), .b(N1594), .O(gate472inter0));
  nand2 gate1078(.a(gate472inter0), .b(s_28), .O(gate472inter1));
  and2  gate1079(.a(N1636), .b(N1594), .O(gate472inter2));
  inv1  gate1080(.a(s_28), .O(gate472inter3));
  inv1  gate1081(.a(s_29), .O(gate472inter4));
  nand2 gate1082(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1083(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1084(.a(N1594), .O(gate472inter7));
  inv1  gate1085(.a(N1636), .O(gate472inter8));
  nand2 gate1086(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1087(.a(s_29), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1088(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1089(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1090(.a(gate472inter12), .b(gate472inter1), .O(N1685));
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );

  xor2  gate1315(.a(N1672), .b(N643), .O(gate476inter0));
  nand2 gate1316(.a(gate476inter0), .b(s_62), .O(gate476inter1));
  and2  gate1317(.a(N1672), .b(N643), .O(gate476inter2));
  inv1  gate1318(.a(s_62), .O(gate476inter3));
  inv1  gate1319(.a(s_63), .O(gate476inter4));
  nand2 gate1320(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1321(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1322(.a(N643), .O(gate476inter7));
  inv1  gate1323(.a(N1672), .O(gate476inter8));
  nand2 gate1324(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1325(.a(s_63), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1326(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1327(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1328(.a(gate476inter12), .b(gate476inter1), .O(N1706));
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );

  xor2  gate1609(.a(N1679), .b(N1028), .O(gate482inter0));
  nand2 gate1610(.a(gate482inter0), .b(s_104), .O(gate482inter1));
  and2  gate1611(.a(N1679), .b(N1028), .O(gate482inter2));
  inv1  gate1612(.a(s_104), .O(gate482inter3));
  inv1  gate1613(.a(s_105), .O(gate482inter4));
  nand2 gate1614(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1615(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1616(.a(N1028), .O(gate482inter7));
  inv1  gate1617(.a(N1679), .O(gate482inter8));
  nand2 gate1618(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1619(.a(s_105), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1620(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1621(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1622(.a(gate482inter12), .b(gate482inter1), .O(N1712));
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );

  xor2  gate1763(.a(N1746), .b(N1708), .O(gate510inter0));
  nand2 gate1764(.a(gate510inter0), .b(s_126), .O(gate510inter1));
  and2  gate1765(.a(N1746), .b(N1708), .O(gate510inter2));
  inv1  gate1766(.a(s_126), .O(gate510inter3));
  inv1  gate1767(.a(s_127), .O(gate510inter4));
  nand2 gate1768(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1769(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1770(.a(N1708), .O(gate510inter7));
  inv1  gate1771(.a(N1746), .O(gate510inter8));
  nand2 gate1772(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1773(.a(s_127), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1774(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1775(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1776(.a(gate510inter12), .b(gate510inter1), .O(N1774));
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );

  xor2  gate895(.a(N1773), .b(N1334), .O(gate523inter0));
  nand2 gate896(.a(gate523inter0), .b(s_2), .O(gate523inter1));
  and2  gate897(.a(N1773), .b(N1334), .O(gate523inter2));
  inv1  gate898(.a(s_2), .O(gate523inter3));
  inv1  gate899(.a(s_3), .O(gate523inter4));
  nand2 gate900(.a(gate523inter4), .b(gate523inter3), .O(gate523inter5));
  nor2  gate901(.a(gate523inter5), .b(gate523inter2), .O(gate523inter6));
  inv1  gate902(.a(N1334), .O(gate523inter7));
  inv1  gate903(.a(N1773), .O(gate523inter8));
  nand2 gate904(.a(gate523inter8), .b(gate523inter7), .O(gate523inter9));
  nand2 gate905(.a(s_3), .b(gate523inter3), .O(gate523inter10));
  nor2  gate906(.a(gate523inter10), .b(gate523inter9), .O(gate523inter11));
  nor2  gate907(.a(gate523inter11), .b(gate523inter6), .O(gate523inter12));
  nand2 gate908(.a(gate523inter12), .b(gate523inter1), .O(N1801));
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate1511(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate1512(.a(gate532inter0), .b(s_90), .O(gate532inter1));
  and2  gate1513(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate1514(.a(s_90), .O(gate532inter3));
  inv1  gate1515(.a(s_91), .O(gate532inter4));
  nand2 gate1516(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate1517(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate1518(.a(N1777), .O(gate532inter7));
  inv1  gate1519(.a(N1490), .O(gate532inter8));
  nand2 gate1520(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate1521(.a(s_91), .b(gate532inter3), .O(gate532inter10));
  nor2  gate1522(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate1523(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate1524(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );

  xor2  gate1581(.a(N1409), .b(N1788), .O(gate537inter0));
  nand2 gate1582(.a(gate537inter0), .b(s_100), .O(gate537inter1));
  and2  gate1583(.a(N1409), .b(N1788), .O(gate537inter2));
  inv1  gate1584(.a(s_100), .O(gate537inter3));
  inv1  gate1585(.a(s_101), .O(gate537inter4));
  nand2 gate1586(.a(gate537inter4), .b(gate537inter3), .O(gate537inter5));
  nor2  gate1587(.a(gate537inter5), .b(gate537inter2), .O(gate537inter6));
  inv1  gate1588(.a(N1788), .O(gate537inter7));
  inv1  gate1589(.a(N1409), .O(gate537inter8));
  nand2 gate1590(.a(gate537inter8), .b(gate537inter7), .O(gate537inter9));
  nand2 gate1591(.a(s_101), .b(gate537inter3), .O(gate537inter10));
  nor2  gate1592(.a(gate537inter10), .b(gate537inter9), .O(gate537inter11));
  nor2  gate1593(.a(gate537inter11), .b(gate537inter6), .O(gate537inter12));
  nand2 gate1594(.a(gate537inter12), .b(gate537inter1), .O(N1826));
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );

  xor2  gate1161(.a(N1787), .b(N1810), .O(gate542inter0));
  nand2 gate1162(.a(gate542inter0), .b(s_40), .O(gate542inter1));
  and2  gate1163(.a(N1787), .b(N1810), .O(gate542inter2));
  inv1  gate1164(.a(s_40), .O(gate542inter3));
  inv1  gate1165(.a(s_41), .O(gate542inter4));
  nand2 gate1166(.a(gate542inter4), .b(gate542inter3), .O(gate542inter5));
  nor2  gate1167(.a(gate542inter5), .b(gate542inter2), .O(gate542inter6));
  inv1  gate1168(.a(N1810), .O(gate542inter7));
  inv1  gate1169(.a(N1787), .O(gate542inter8));
  nand2 gate1170(.a(gate542inter8), .b(gate542inter7), .O(gate542inter9));
  nand2 gate1171(.a(s_41), .b(gate542inter3), .O(gate542inter10));
  nor2  gate1172(.a(gate542inter10), .b(gate542inter9), .O(gate542inter11));
  nor2  gate1173(.a(gate542inter11), .b(gate542inter6), .O(gate542inter12));
  nand2 gate1174(.a(gate542inter12), .b(gate542inter1), .O(N1841));
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );

  xor2  gate1903(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate1904(.a(gate547inter0), .b(s_146), .O(gate547inter1));
  and2  gate1905(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate1906(.a(s_146), .O(gate547inter3));
  inv1  gate1907(.a(s_147), .O(gate547inter4));
  nand2 gate1908(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate1909(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate1910(.a(N1815), .O(gate547inter7));
  inv1  gate1911(.a(N1707), .O(gate547inter8));
  nand2 gate1912(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate1913(.a(s_147), .b(gate547inter3), .O(gate547inter10));
  nor2  gate1914(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate1915(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate1916(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );

  xor2  gate993(.a(N1768), .b(N1841), .O(gate559inter0));
  nand2 gate994(.a(gate559inter0), .b(s_16), .O(gate559inter1));
  and2  gate995(.a(N1768), .b(N1841), .O(gate559inter2));
  inv1  gate996(.a(s_16), .O(gate559inter3));
  inv1  gate997(.a(s_17), .O(gate559inter4));
  nand2 gate998(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate999(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate1000(.a(N1841), .O(gate559inter7));
  inv1  gate1001(.a(N1768), .O(gate559inter8));
  nand2 gate1002(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate1003(.a(s_17), .b(gate559inter3), .O(gate559inter10));
  nor2  gate1004(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate1005(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate1006(.a(gate559inter12), .b(gate559inter1), .O(N1882));
inv1 gate560( .a(N1841), .O(N1883) );

  xor2  gate1133(.a(N1852), .b(N1826), .O(gate561inter0));
  nand2 gate1134(.a(gate561inter0), .b(s_36), .O(gate561inter1));
  and2  gate1135(.a(N1852), .b(N1826), .O(gate561inter2));
  inv1  gate1136(.a(s_36), .O(gate561inter3));
  inv1  gate1137(.a(s_37), .O(gate561inter4));
  nand2 gate1138(.a(gate561inter4), .b(gate561inter3), .O(gate561inter5));
  nor2  gate1139(.a(gate561inter5), .b(gate561inter2), .O(gate561inter6));
  inv1  gate1140(.a(N1826), .O(gate561inter7));
  inv1  gate1141(.a(N1852), .O(gate561inter8));
  nand2 gate1142(.a(gate561inter8), .b(gate561inter7), .O(gate561inter9));
  nand2 gate1143(.a(s_37), .b(gate561inter3), .O(gate561inter10));
  nor2  gate1144(.a(gate561inter10), .b(gate561inter9), .O(gate561inter11));
  nor2  gate1145(.a(gate561inter11), .b(gate561inter6), .O(gate561inter12));
  nand2 gate1146(.a(gate561inter12), .b(gate561inter1), .O(N1884));
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );

  xor2  gate1665(.a(N1864), .b(N1640), .O(gate566inter0));
  nand2 gate1666(.a(gate566inter0), .b(s_112), .O(gate566inter1));
  and2  gate1667(.a(N1864), .b(N1640), .O(gate566inter2));
  inv1  gate1668(.a(s_112), .O(gate566inter3));
  inv1  gate1669(.a(s_113), .O(gate566inter4));
  nand2 gate1670(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate1671(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate1672(.a(N1640), .O(gate566inter7));
  inv1  gate1673(.a(N1864), .O(gate566inter8));
  nand2 gate1674(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate1675(.a(s_113), .b(gate566inter3), .O(gate566inter10));
  nor2  gate1676(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate1677(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate1678(.a(gate566inter12), .b(gate566inter1), .O(N1897));
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );

  xor2  gate979(.a(N1911), .b(N1882), .O(gate583inter0));
  nand2 gate980(.a(gate583inter0), .b(s_14), .O(gate583inter1));
  and2  gate981(.a(N1911), .b(N1882), .O(gate583inter2));
  inv1  gate982(.a(s_14), .O(gate583inter3));
  inv1  gate983(.a(s_15), .O(gate583inter4));
  nand2 gate984(.a(gate583inter4), .b(gate583inter3), .O(gate583inter5));
  nor2  gate985(.a(gate583inter5), .b(gate583inter2), .O(gate583inter6));
  inv1  gate986(.a(N1882), .O(gate583inter7));
  inv1  gate987(.a(N1911), .O(gate583inter8));
  nand2 gate988(.a(gate583inter8), .b(gate583inter7), .O(gate583inter9));
  nand2 gate989(.a(s_15), .b(gate583inter3), .O(gate583inter10));
  nor2  gate990(.a(gate583inter10), .b(gate583inter9), .O(gate583inter11));
  nor2  gate991(.a(gate583inter11), .b(gate583inter6), .O(gate583inter12));
  nand2 gate992(.a(gate583inter12), .b(gate583inter1), .O(N1936));
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );

  xor2  gate1455(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate1456(.a(gate601inter0), .b(s_82), .O(gate601inter1));
  and2  gate1457(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate1458(.a(s_82), .O(gate601inter3));
  inv1  gate1459(.a(s_83), .O(gate601inter4));
  nand2 gate1460(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate1461(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate1462(.a(N1921), .O(gate601inter7));
  inv1  gate1463(.a(N1942), .O(gate601inter8));
  nand2 gate1464(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate1465(.a(s_83), .b(gate601inter3), .O(gate601inter10));
  nor2  gate1466(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate1467(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate1468(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );

  xor2  gate1483(.a(N1937), .b(N1944), .O(gate605inter0));
  nand2 gate1484(.a(gate605inter0), .b(s_86), .O(gate605inter1));
  and2  gate1485(.a(N1937), .b(N1944), .O(gate605inter2));
  inv1  gate1486(.a(s_86), .O(gate605inter3));
  inv1  gate1487(.a(s_87), .O(gate605inter4));
  nand2 gate1488(.a(gate605inter4), .b(gate605inter3), .O(gate605inter5));
  nor2  gate1489(.a(gate605inter5), .b(gate605inter2), .O(gate605inter6));
  inv1  gate1490(.a(N1944), .O(gate605inter7));
  inv1  gate1491(.a(N1937), .O(gate605inter8));
  nand2 gate1492(.a(gate605inter8), .b(gate605inter7), .O(gate605inter9));
  nand2 gate1493(.a(s_87), .b(gate605inter3), .O(gate605inter10));
  nor2  gate1494(.a(gate605inter10), .b(gate605inter9), .O(gate605inter11));
  nor2  gate1495(.a(gate605inter11), .b(gate605inter6), .O(gate605inter12));
  nand2 gate1496(.a(gate605inter12), .b(gate605inter1), .O(N2000));
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );

  xor2  gate1357(.a(N1350), .b(N1953), .O(gate608inter0));
  nand2 gate1358(.a(gate608inter0), .b(s_68), .O(gate608inter1));
  and2  gate1359(.a(N1350), .b(N1953), .O(gate608inter2));
  inv1  gate1360(.a(s_68), .O(gate608inter3));
  inv1  gate1361(.a(s_69), .O(gate608inter4));
  nand2 gate1362(.a(gate608inter4), .b(gate608inter3), .O(gate608inter5));
  nor2  gate1363(.a(gate608inter5), .b(gate608inter2), .O(gate608inter6));
  inv1  gate1364(.a(N1953), .O(gate608inter7));
  inv1  gate1365(.a(N1350), .O(gate608inter8));
  nand2 gate1366(.a(gate608inter8), .b(gate608inter7), .O(gate608inter9));
  nand2 gate1367(.a(s_69), .b(gate608inter3), .O(gate608inter10));
  nor2  gate1368(.a(gate608inter10), .b(gate608inter9), .O(gate608inter11));
  nor2  gate1369(.a(gate608inter11), .b(gate608inter6), .O(gate608inter12));
  nand2 gate1370(.a(gate608inter12), .b(gate608inter1), .O(N2004));
inv1 gate609( .a(N1953), .O(N2005) );

  xor2  gate1707(.a(N1351), .b(N1950), .O(gate610inter0));
  nand2 gate1708(.a(gate610inter0), .b(s_118), .O(gate610inter1));
  and2  gate1709(.a(N1351), .b(N1950), .O(gate610inter2));
  inv1  gate1710(.a(s_118), .O(gate610inter3));
  inv1  gate1711(.a(s_119), .O(gate610inter4));
  nand2 gate1712(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate1713(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate1714(.a(N1950), .O(gate610inter7));
  inv1  gate1715(.a(N1351), .O(gate610inter8));
  nand2 gate1716(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate1717(.a(s_119), .b(gate610inter3), .O(gate610inter10));
  nor2  gate1718(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate1719(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate1720(.a(gate610inter12), .b(gate610inter1), .O(N2006));
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );

  xor2  gate1749(.a(N1591), .b(N1987), .O(gate623inter0));
  nand2 gate1750(.a(gate623inter0), .b(s_124), .O(gate623inter1));
  and2  gate1751(.a(N1591), .b(N1987), .O(gate623inter2));
  inv1  gate1752(.a(s_124), .O(gate623inter3));
  inv1  gate1753(.a(s_125), .O(gate623inter4));
  nand2 gate1754(.a(gate623inter4), .b(gate623inter3), .O(gate623inter5));
  nor2  gate1755(.a(gate623inter5), .b(gate623inter2), .O(gate623inter6));
  inv1  gate1756(.a(N1987), .O(gate623inter7));
  inv1  gate1757(.a(N1591), .O(gate623inter8));
  nand2 gate1758(.a(gate623inter8), .b(gate623inter7), .O(gate623inter9));
  nand2 gate1759(.a(s_125), .b(gate623inter3), .O(gate623inter10));
  nor2  gate1760(.a(gate623inter10), .b(gate623inter9), .O(gate623inter11));
  nor2  gate1761(.a(gate623inter11), .b(gate623inter6), .O(gate623inter12));
  nand2 gate1762(.a(gate623inter12), .b(gate623inter1), .O(N2022));
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );

  xor2  gate923(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate924(.a(gate634inter0), .b(s_6), .O(gate634inter1));
  and2  gate925(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate926(.a(s_6), .O(gate634inter3));
  inv1  gate927(.a(s_7), .O(gate634inter4));
  nand2 gate928(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate929(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate930(.a(N1534), .O(gate634inter7));
  inv1  gate931(.a(N2021), .O(gate634inter8));
  nand2 gate932(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate933(.a(s_7), .b(gate634inter3), .O(gate634inter10));
  nor2  gate934(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate935(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate936(.a(gate634inter12), .b(gate634inter1), .O(N2039));
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );

  xor2  gate1623(.a(N2024), .b(N2004), .O(gate636inter0));
  nand2 gate1624(.a(gate636inter0), .b(s_106), .O(gate636inter1));
  and2  gate1625(.a(N2024), .b(N2004), .O(gate636inter2));
  inv1  gate1626(.a(s_106), .O(gate636inter3));
  inv1  gate1627(.a(s_107), .O(gate636inter4));
  nand2 gate1628(.a(gate636inter4), .b(gate636inter3), .O(gate636inter5));
  nor2  gate1629(.a(gate636inter5), .b(gate636inter2), .O(gate636inter6));
  inv1  gate1630(.a(N2004), .O(gate636inter7));
  inv1  gate1631(.a(N2024), .O(gate636inter8));
  nand2 gate1632(.a(gate636inter8), .b(gate636inter7), .O(gate636inter9));
  nand2 gate1633(.a(s_107), .b(gate636inter3), .O(gate636inter10));
  nor2  gate1634(.a(gate636inter10), .b(gate636inter9), .O(gate636inter11));
  nor2  gate1635(.a(gate636inter11), .b(gate636inter6), .O(gate636inter12));
  nand2 gate1636(.a(gate636inter12), .b(gate636inter1), .O(N2041));
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );

  xor2  gate1343(.a(N290), .b(N2060), .O(gate649inter0));
  nand2 gate1344(.a(gate649inter0), .b(s_66), .O(gate649inter1));
  and2  gate1345(.a(N290), .b(N2060), .O(gate649inter2));
  inv1  gate1346(.a(s_66), .O(gate649inter3));
  inv1  gate1347(.a(s_67), .O(gate649inter4));
  nand2 gate1348(.a(gate649inter4), .b(gate649inter3), .O(gate649inter5));
  nor2  gate1349(.a(gate649inter5), .b(gate649inter2), .O(gate649inter6));
  inv1  gate1350(.a(N2060), .O(gate649inter7));
  inv1  gate1351(.a(N290), .O(gate649inter8));
  nand2 gate1352(.a(gate649inter8), .b(gate649inter7), .O(gate649inter9));
  nand2 gate1353(.a(s_67), .b(gate649inter3), .O(gate649inter10));
  nor2  gate1354(.a(gate649inter10), .b(gate649inter9), .O(gate649inter11));
  nor2  gate1355(.a(gate649inter11), .b(gate649inter6), .O(gate649inter12));
  nand2 gate1356(.a(gate649inter12), .b(gate649inter1), .O(N2078));

  xor2  gate1203(.a(N290), .b(N2061), .O(gate650inter0));
  nand2 gate1204(.a(gate650inter0), .b(s_46), .O(gate650inter1));
  and2  gate1205(.a(N290), .b(N2061), .O(gate650inter2));
  inv1  gate1206(.a(s_46), .O(gate650inter3));
  inv1  gate1207(.a(s_47), .O(gate650inter4));
  nand2 gate1208(.a(gate650inter4), .b(gate650inter3), .O(gate650inter5));
  nor2  gate1209(.a(gate650inter5), .b(gate650inter2), .O(gate650inter6));
  inv1  gate1210(.a(N2061), .O(gate650inter7));
  inv1  gate1211(.a(N290), .O(gate650inter8));
  nand2 gate1212(.a(gate650inter8), .b(gate650inter7), .O(gate650inter9));
  nand2 gate1213(.a(s_47), .b(gate650inter3), .O(gate650inter10));
  nor2  gate1214(.a(gate650inter10), .b(gate650inter9), .O(gate650inter11));
  nor2  gate1215(.a(gate650inter11), .b(gate650inter6), .O(gate650inter12));
  nand2 gate1216(.a(gate650inter12), .b(gate650inter1), .O(N2081));
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate1021(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate1022(.a(gate671inter0), .b(s_20), .O(gate671inter1));
  and2  gate1023(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate1024(.a(s_20), .O(gate671inter3));
  inv1  gate1025(.a(s_21), .O(gate671inter4));
  nand2 gate1026(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate1027(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate1028(.a(N2205), .O(gate671inter7));
  inv1  gate1029(.a(N913), .O(gate671inter8));
  nand2 gate1030(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate1031(.a(s_21), .b(gate671inter3), .O(gate671inter10));
  nor2  gate1032(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate1033(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate1034(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );

  xor2  gate1525(.a(N2227), .b(N661), .O(gate679inter0));
  nand2 gate1526(.a(gate679inter0), .b(s_92), .O(gate679inter1));
  and2  gate1527(.a(N2227), .b(N661), .O(gate679inter2));
  inv1  gate1528(.a(s_92), .O(gate679inter3));
  inv1  gate1529(.a(s_93), .O(gate679inter4));
  nand2 gate1530(.a(gate679inter4), .b(gate679inter3), .O(gate679inter5));
  nor2  gate1531(.a(gate679inter5), .b(gate679inter2), .O(gate679inter6));
  inv1  gate1532(.a(N661), .O(gate679inter7));
  inv1  gate1533(.a(N2227), .O(gate679inter8));
  nand2 gate1534(.a(gate679inter8), .b(gate679inter7), .O(gate679inter9));
  nand2 gate1535(.a(s_93), .b(gate679inter3), .O(gate679inter10));
  nor2  gate1536(.a(gate679inter10), .b(gate679inter9), .O(gate679inter11));
  nor2  gate1537(.a(gate679inter11), .b(gate679inter6), .O(gate679inter12));
  nand2 gate1538(.a(gate679inter12), .b(gate679inter1), .O(N2234));
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );

  xor2  gate1777(.a(N2230), .b(N2214), .O(gate681inter0));
  nand2 gate1778(.a(gate681inter0), .b(s_128), .O(gate681inter1));
  and2  gate1779(.a(N2230), .b(N2214), .O(gate681inter2));
  inv1  gate1780(.a(s_128), .O(gate681inter3));
  inv1  gate1781(.a(s_129), .O(gate681inter4));
  nand2 gate1782(.a(gate681inter4), .b(gate681inter3), .O(gate681inter5));
  nor2  gate1783(.a(gate681inter5), .b(gate681inter2), .O(gate681inter6));
  inv1  gate1784(.a(N2214), .O(gate681inter7));
  inv1  gate1785(.a(N2230), .O(gate681inter8));
  nand2 gate1786(.a(gate681inter8), .b(gate681inter7), .O(gate681inter9));
  nand2 gate1787(.a(s_129), .b(gate681inter3), .O(gate681inter10));
  nor2  gate1788(.a(gate681inter10), .b(gate681inter9), .O(gate681inter11));
  nor2  gate1789(.a(gate681inter11), .b(gate681inter6), .O(gate681inter12));
  nand2 gate1790(.a(gate681inter12), .b(gate681inter1), .O(N2236));

  xor2  gate1553(.a(N2231), .b(N2216), .O(gate682inter0));
  nand2 gate1554(.a(gate682inter0), .b(s_96), .O(gate682inter1));
  and2  gate1555(.a(N2231), .b(N2216), .O(gate682inter2));
  inv1  gate1556(.a(s_96), .O(gate682inter3));
  inv1  gate1557(.a(s_97), .O(gate682inter4));
  nand2 gate1558(.a(gate682inter4), .b(gate682inter3), .O(gate682inter5));
  nor2  gate1559(.a(gate682inter5), .b(gate682inter2), .O(gate682inter6));
  inv1  gate1560(.a(N2216), .O(gate682inter7));
  inv1  gate1561(.a(N2231), .O(gate682inter8));
  nand2 gate1562(.a(gate682inter8), .b(gate682inter7), .O(gate682inter9));
  nand2 gate1563(.a(s_97), .b(gate682inter3), .O(gate682inter10));
  nor2  gate1564(.a(gate682inter10), .b(gate682inter9), .O(gate682inter11));
  nor2  gate1565(.a(gate682inter11), .b(gate682inter6), .O(gate682inter12));
  nand2 gate1566(.a(gate682inter12), .b(gate682inter1), .O(N2237));

  xor2  gate1987(.a(N2232), .b(N2222), .O(gate683inter0));
  nand2 gate1988(.a(gate683inter0), .b(s_158), .O(gate683inter1));
  and2  gate1989(.a(N2232), .b(N2222), .O(gate683inter2));
  inv1  gate1990(.a(s_158), .O(gate683inter3));
  inv1  gate1991(.a(s_159), .O(gate683inter4));
  nand2 gate1992(.a(gate683inter4), .b(gate683inter3), .O(gate683inter5));
  nor2  gate1993(.a(gate683inter5), .b(gate683inter2), .O(gate683inter6));
  inv1  gate1994(.a(N2222), .O(gate683inter7));
  inv1  gate1995(.a(N2232), .O(gate683inter8));
  nand2 gate1996(.a(gate683inter8), .b(gate683inter7), .O(gate683inter9));
  nand2 gate1997(.a(s_159), .b(gate683inter3), .O(gate683inter10));
  nor2  gate1998(.a(gate683inter10), .b(gate683inter9), .O(gate683inter11));
  nor2  gate1999(.a(gate683inter11), .b(gate683inter6), .O(gate683inter12));
  nand2 gate2000(.a(gate683inter12), .b(gate683inter1), .O(N2240));

  xor2  gate1371(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate1372(.a(gate684inter0), .b(s_70), .O(gate684inter1));
  and2  gate1373(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate1374(.a(s_70), .O(gate684inter3));
  inv1  gate1375(.a(s_71), .O(gate684inter4));
  nand2 gate1376(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate1377(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate1378(.a(N2224), .O(gate684inter7));
  inv1  gate1379(.a(N2233), .O(gate684inter8));
  nand2 gate1380(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate1381(.a(s_71), .b(gate684inter3), .O(gate684inter10));
  nor2  gate1382(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate1383(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate1384(.a(gate684inter12), .b(gate684inter1), .O(N2241));
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );

  xor2  gate1861(.a(N548), .b(N2573), .O(gate760inter0));
  nand2 gate1862(.a(gate760inter0), .b(s_140), .O(gate760inter1));
  and2  gate1863(.a(N548), .b(N2573), .O(gate760inter2));
  inv1  gate1864(.a(s_140), .O(gate760inter3));
  inv1  gate1865(.a(s_141), .O(gate760inter4));
  nand2 gate1866(.a(gate760inter4), .b(gate760inter3), .O(gate760inter5));
  nor2  gate1867(.a(gate760inter5), .b(gate760inter2), .O(gate760inter6));
  inv1  gate1868(.a(N2573), .O(gate760inter7));
  inv1  gate1869(.a(N548), .O(gate760inter8));
  nand2 gate1870(.a(gate760inter8), .b(gate760inter7), .O(gate760inter9));
  nand2 gate1871(.a(s_141), .b(gate760inter3), .O(gate760inter10));
  nor2  gate1872(.a(gate760inter10), .b(gate760inter9), .O(gate760inter11));
  nor2  gate1873(.a(gate760inter11), .b(gate760inter6), .O(gate760inter12));
  nand2 gate1874(.a(gate760inter12), .b(gate760inter1), .O(N2688));
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );

  xor2  gate1175(.a(N2723), .b(N2675), .O(gate797inter0));
  nand2 gate1176(.a(gate797inter0), .b(s_42), .O(gate797inter1));
  and2  gate1177(.a(N2723), .b(N2675), .O(gate797inter2));
  inv1  gate1178(.a(s_42), .O(gate797inter3));
  inv1  gate1179(.a(s_43), .O(gate797inter4));
  nand2 gate1180(.a(gate797inter4), .b(gate797inter3), .O(gate797inter5));
  nor2  gate1181(.a(gate797inter5), .b(gate797inter2), .O(gate797inter6));
  inv1  gate1182(.a(N2675), .O(gate797inter7));
  inv1  gate1183(.a(N2723), .O(gate797inter8));
  nand2 gate1184(.a(gate797inter8), .b(gate797inter7), .O(gate797inter9));
  nand2 gate1185(.a(s_43), .b(gate797inter3), .O(gate797inter10));
  nor2  gate1186(.a(gate797inter10), .b(gate797inter9), .O(gate797inter11));
  nor2  gate1187(.a(gate797inter11), .b(gate797inter6), .O(gate797inter12));
  nand2 gate1188(.a(gate797inter12), .b(gate797inter1), .O(N2756));

  xor2  gate1833(.a(N2725), .b(N355), .O(gate798inter0));
  nand2 gate1834(.a(gate798inter0), .b(s_136), .O(gate798inter1));
  and2  gate1835(.a(N2725), .b(N355), .O(gate798inter2));
  inv1  gate1836(.a(s_136), .O(gate798inter3));
  inv1  gate1837(.a(s_137), .O(gate798inter4));
  nand2 gate1838(.a(gate798inter4), .b(gate798inter3), .O(gate798inter5));
  nor2  gate1839(.a(gate798inter5), .b(gate798inter2), .O(gate798inter6));
  inv1  gate1840(.a(N355), .O(gate798inter7));
  inv1  gate1841(.a(N2725), .O(gate798inter8));
  nand2 gate1842(.a(gate798inter8), .b(gate798inter7), .O(gate798inter9));
  nand2 gate1843(.a(s_137), .b(gate798inter3), .O(gate798inter10));
  nor2  gate1844(.a(gate798inter10), .b(gate798inter9), .O(gate798inter11));
  nor2  gate1845(.a(gate798inter11), .b(gate798inter6), .O(gate798inter12));
  nand2 gate1846(.a(gate798inter12), .b(gate798inter1), .O(N2757));
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );

  xor2  gate1427(.a(N2743), .b(N2688), .O(gate808inter0));
  nand2 gate1428(.a(gate808inter0), .b(s_78), .O(gate808inter1));
  and2  gate1429(.a(N2743), .b(N2688), .O(gate808inter2));
  inv1  gate1430(.a(s_78), .O(gate808inter3));
  inv1  gate1431(.a(s_79), .O(gate808inter4));
  nand2 gate1432(.a(gate808inter4), .b(gate808inter3), .O(gate808inter5));
  nor2  gate1433(.a(gate808inter5), .b(gate808inter2), .O(gate808inter6));
  inv1  gate1434(.a(N2688), .O(gate808inter7));
  inv1  gate1435(.a(N2743), .O(gate808inter8));
  nand2 gate1436(.a(gate808inter8), .b(gate808inter7), .O(gate808inter9));
  nand2 gate1437(.a(s_79), .b(gate808inter3), .O(gate808inter10));
  nor2  gate1438(.a(gate808inter10), .b(gate808inter9), .O(gate808inter11));
  nor2  gate1439(.a(gate808inter11), .b(gate808inter6), .O(gate808inter12));
  nand2 gate1440(.a(gate808inter12), .b(gate808inter1), .O(N2767));
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );

  xor2  gate1973(.a(N2766), .b(N2741), .O(gate820inter0));
  nand2 gate1974(.a(gate820inter0), .b(s_156), .O(gate820inter1));
  and2  gate1975(.a(N2766), .b(N2741), .O(gate820inter2));
  inv1  gate1976(.a(s_156), .O(gate820inter3));
  inv1  gate1977(.a(s_157), .O(gate820inter4));
  nand2 gate1978(.a(gate820inter4), .b(gate820inter3), .O(gate820inter5));
  nor2  gate1979(.a(gate820inter5), .b(gate820inter2), .O(gate820inter6));
  inv1  gate1980(.a(N2741), .O(gate820inter7));
  inv1  gate1981(.a(N2766), .O(gate820inter8));
  nand2 gate1982(.a(gate820inter8), .b(gate820inter7), .O(gate820inter9));
  nand2 gate1983(.a(s_157), .b(gate820inter3), .O(gate820inter10));
  nor2  gate1984(.a(gate820inter10), .b(gate820inter9), .O(gate820inter11));
  nor2  gate1985(.a(gate820inter11), .b(gate820inter6), .O(gate820inter12));
  nand2 gate1986(.a(gate820inter12), .b(gate820inter1), .O(N2787));
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );

  xor2  gate1875(.a(N2750), .b(N2747), .O(gate822inter0));
  nand2 gate1876(.a(gate822inter0), .b(s_142), .O(gate822inter1));
  and2  gate1877(.a(N2750), .b(N2747), .O(gate822inter2));
  inv1  gate1878(.a(s_142), .O(gate822inter3));
  inv1  gate1879(.a(s_143), .O(gate822inter4));
  nand2 gate1880(.a(gate822inter4), .b(gate822inter3), .O(gate822inter5));
  nor2  gate1881(.a(gate822inter5), .b(gate822inter2), .O(gate822inter6));
  inv1  gate1882(.a(N2747), .O(gate822inter7));
  inv1  gate1883(.a(N2750), .O(gate822inter8));
  nand2 gate1884(.a(gate822inter8), .b(gate822inter7), .O(gate822inter9));
  nand2 gate1885(.a(s_143), .b(gate822inter3), .O(gate822inter10));
  nor2  gate1886(.a(gate822inter10), .b(gate822inter9), .O(gate822inter11));
  nor2  gate1887(.a(gate822inter11), .b(gate822inter6), .O(gate822inter12));
  nand2 gate1888(.a(gate822inter12), .b(gate822inter1), .O(N2789));
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );

  xor2  gate1105(.a(N2018), .b(N2773), .O(gate824inter0));
  nand2 gate1106(.a(gate824inter0), .b(s_32), .O(gate824inter1));
  and2  gate1107(.a(N2018), .b(N2773), .O(gate824inter2));
  inv1  gate1108(.a(s_32), .O(gate824inter3));
  inv1  gate1109(.a(s_33), .O(gate824inter4));
  nand2 gate1110(.a(gate824inter4), .b(gate824inter3), .O(gate824inter5));
  nor2  gate1111(.a(gate824inter5), .b(gate824inter2), .O(gate824inter6));
  inv1  gate1112(.a(N2773), .O(gate824inter7));
  inv1  gate1113(.a(N2018), .O(gate824inter8));
  nand2 gate1114(.a(gate824inter8), .b(gate824inter7), .O(gate824inter9));
  nand2 gate1115(.a(s_33), .b(gate824inter3), .O(gate824inter10));
  nor2  gate1116(.a(gate824inter10), .b(gate824inter9), .O(gate824inter11));
  nor2  gate1117(.a(gate824inter11), .b(gate824inter6), .O(gate824inter12));
  nand2 gate1118(.a(gate824inter12), .b(gate824inter1), .O(N2807));
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );

  xor2  gate1413(.a(N2810), .b(N1968), .O(gate835inter0));
  nand2 gate1414(.a(gate835inter0), .b(s_76), .O(gate835inter1));
  and2  gate1415(.a(N2810), .b(N1968), .O(gate835inter2));
  inv1  gate1416(.a(s_76), .O(gate835inter3));
  inv1  gate1417(.a(s_77), .O(gate835inter4));
  nand2 gate1418(.a(gate835inter4), .b(gate835inter3), .O(gate835inter5));
  nor2  gate1419(.a(gate835inter5), .b(gate835inter2), .O(gate835inter6));
  inv1  gate1420(.a(N1968), .O(gate835inter7));
  inv1  gate1421(.a(N2810), .O(gate835inter8));
  nand2 gate1422(.a(gate835inter8), .b(gate835inter7), .O(gate835inter9));
  nand2 gate1423(.a(s_77), .b(gate835inter3), .O(gate835inter10));
  nor2  gate1424(.a(gate835inter10), .b(gate835inter9), .O(gate835inter11));
  nor2  gate1425(.a(gate835inter11), .b(gate835inter6), .O(gate835inter12));
  nand2 gate1426(.a(gate835inter12), .b(gate835inter1), .O(N2828));
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );

  xor2  gate1945(.a(N2827), .b(N2807), .O(gate837inter0));
  nand2 gate1946(.a(gate837inter0), .b(s_152), .O(gate837inter1));
  and2  gate1947(.a(N2827), .b(N2807), .O(gate837inter2));
  inv1  gate1948(.a(s_152), .O(gate837inter3));
  inv1  gate1949(.a(s_153), .O(gate837inter4));
  nand2 gate1950(.a(gate837inter4), .b(gate837inter3), .O(gate837inter5));
  nor2  gate1951(.a(gate837inter5), .b(gate837inter2), .O(gate837inter6));
  inv1  gate1952(.a(N2807), .O(gate837inter7));
  inv1  gate1953(.a(N2827), .O(gate837inter8));
  nand2 gate1954(.a(gate837inter8), .b(gate837inter7), .O(gate837inter9));
  nand2 gate1955(.a(s_153), .b(gate837inter3), .O(gate837inter10));
  nor2  gate1956(.a(gate837inter10), .b(gate837inter9), .O(gate837inter11));
  nor2  gate1957(.a(gate837inter11), .b(gate837inter6), .O(gate837inter12));
  nand2 gate1958(.a(gate837inter12), .b(gate837inter1), .O(N2843));
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );

  xor2  gate937(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate938(.a(gate839inter0), .b(s_8), .O(gate839inter1));
  and2  gate939(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate940(.a(s_8), .O(gate839inter3));
  inv1  gate941(.a(s_9), .O(gate839inter4));
  nand2 gate942(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate943(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate944(.a(N2812), .O(gate839inter7));
  inv1  gate945(.a(N2076), .O(gate839inter8));
  nand2 gate946(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate947(.a(s_9), .b(gate839inter3), .O(gate839inter10));
  nor2  gate948(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate949(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate950(.a(gate839inter12), .b(gate839inter1), .O(N2850));

  xor2  gate2001(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate2002(.a(gate840inter0), .b(s_160), .O(gate840inter1));
  and2  gate2003(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate2004(.a(s_160), .O(gate840inter3));
  inv1  gate2005(.a(s_161), .O(gate840inter4));
  nand2 gate2006(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate2007(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate2008(.a(N2815), .O(gate840inter7));
  inv1  gate2009(.a(N2077), .O(gate840inter8));
  nand2 gate2010(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate2011(.a(s_161), .b(gate840inter3), .O(gate840inter10));
  nor2  gate2012(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate2013(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate2014(.a(gate840inter12), .b(gate840inter1), .O(N2851));
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );

  xor2  gate1637(.a(N1985), .b(N2829), .O(gate850inter0));
  nand2 gate1638(.a(gate850inter0), .b(s_108), .O(gate850inter1));
  and2  gate1639(.a(N1985), .b(N2829), .O(gate850inter2));
  inv1  gate1640(.a(s_108), .O(gate850inter3));
  inv1  gate1641(.a(s_109), .O(gate850inter4));
  nand2 gate1642(.a(gate850inter4), .b(gate850inter3), .O(gate850inter5));
  nor2  gate1643(.a(gate850inter5), .b(gate850inter2), .O(gate850inter6));
  inv1  gate1644(.a(N2829), .O(gate850inter7));
  inv1  gate1645(.a(N1985), .O(gate850inter8));
  nand2 gate1646(.a(gate850inter8), .b(gate850inter7), .O(gate850inter9));
  nand2 gate1647(.a(s_109), .b(gate850inter3), .O(gate850inter10));
  nor2  gate1648(.a(gate850inter10), .b(gate850inter9), .O(gate850inter11));
  nor2  gate1649(.a(gate850inter11), .b(gate850inter6), .O(gate850inter12));
  nand2 gate1650(.a(gate850inter12), .b(gate850inter1), .O(N2863));
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate1693(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate1694(.a(gate860inter0), .b(s_116), .O(gate860inter1));
  and2  gate1695(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate1696(.a(s_116), .O(gate860inter3));
  inv1  gate1697(.a(s_117), .O(gate860inter4));
  nand2 gate1698(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate1699(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate1700(.a(N1933), .O(gate860inter7));
  inv1  gate1701(.a(N2862), .O(gate860inter8));
  nand2 gate1702(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate1703(.a(s_117), .b(gate860inter3), .O(gate860inter10));
  nor2  gate1704(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate1705(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate1706(.a(gate860inter12), .b(gate860inter1), .O(N2875));
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );

  xor2  gate1301(.a(N2853), .b(N2869), .O(gate864inter0));
  nand2 gate1302(.a(gate864inter0), .b(s_60), .O(gate864inter1));
  and2  gate1303(.a(N2853), .b(N2869), .O(gate864inter2));
  inv1  gate1304(.a(s_60), .O(gate864inter3));
  inv1  gate1305(.a(s_61), .O(gate864inter4));
  nand2 gate1306(.a(gate864inter4), .b(gate864inter3), .O(gate864inter5));
  nor2  gate1307(.a(gate864inter5), .b(gate864inter2), .O(gate864inter6));
  inv1  gate1308(.a(N2869), .O(gate864inter7));
  inv1  gate1309(.a(N2853), .O(gate864inter8));
  nand2 gate1310(.a(gate864inter8), .b(gate864inter7), .O(gate864inter9));
  nand2 gate1311(.a(s_61), .b(gate864inter3), .O(gate864inter10));
  nor2  gate1312(.a(gate864inter10), .b(gate864inter9), .O(gate864inter11));
  nor2  gate1313(.a(gate864inter11), .b(gate864inter6), .O(gate864inter12));
  nand2 gate1314(.a(gate864inter12), .b(gate864inter1), .O(N2879));

  xor2  gate1959(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate1960(.a(gate865inter0), .b(s_154), .O(gate865inter1));
  and2  gate1961(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate1962(.a(s_154), .O(gate865inter3));
  inv1  gate1963(.a(s_155), .O(gate865inter4));
  nand2 gate1964(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate1965(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate1966(.a(N2870), .O(gate865inter7));
  inv1  gate1967(.a(N2854), .O(gate865inter8));
  nand2 gate1968(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate1969(.a(s_155), .b(gate865inter3), .O(gate865inter10));
  nor2  gate1970(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate1971(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate1972(.a(gate865inter12), .b(gate865inter1), .O(N2880));
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate1917(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate1918(.a(gate874inter0), .b(s_148), .O(gate874inter1));
  and2  gate1919(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate1920(.a(s_148), .O(gate874inter3));
  inv1  gate1921(.a(s_149), .O(gate874inter4));
  nand2 gate1922(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate1923(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate1924(.a(N2871), .O(gate874inter7));
  inv1  gate1925(.a(N2881), .O(gate874inter8));
  nand2 gate1926(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate1927(.a(s_149), .b(gate874inter3), .O(gate874inter10));
  nor2  gate1928(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate1929(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate1930(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule