module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate589(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate590(.a(gate24inter0), .b(s_6), .O(gate24inter1));
  and2  gate591(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate592(.a(s_6), .O(gate24inter3));
  inv1  gate593(.a(s_7), .O(gate24inter4));
  nand2 gate594(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate595(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate596(.a(G31), .O(gate24inter7));
  inv1  gate597(.a(G32), .O(gate24inter8));
  nand2 gate598(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate599(.a(s_7), .b(gate24inter3), .O(gate24inter10));
  nor2  gate600(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate601(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate602(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1387(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1388(.a(gate25inter0), .b(s_120), .O(gate25inter1));
  and2  gate1389(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1390(.a(s_120), .O(gate25inter3));
  inv1  gate1391(.a(s_121), .O(gate25inter4));
  nand2 gate1392(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1393(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1394(.a(G1), .O(gate25inter7));
  inv1  gate1395(.a(G5), .O(gate25inter8));
  nand2 gate1396(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1397(.a(s_121), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1398(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1399(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1400(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate575(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate576(.a(gate40inter0), .b(s_4), .O(gate40inter1));
  and2  gate577(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate578(.a(s_4), .O(gate40inter3));
  inv1  gate579(.a(s_5), .O(gate40inter4));
  nand2 gate580(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate581(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate582(.a(G28), .O(gate40inter7));
  inv1  gate583(.a(G32), .O(gate40inter8));
  nand2 gate584(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate585(.a(s_5), .b(gate40inter3), .O(gate40inter10));
  nor2  gate586(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate587(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate588(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate911(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate912(.a(gate49inter0), .b(s_52), .O(gate49inter1));
  and2  gate913(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate914(.a(s_52), .O(gate49inter3));
  inv1  gate915(.a(s_53), .O(gate49inter4));
  nand2 gate916(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate917(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate918(.a(G9), .O(gate49inter7));
  inv1  gate919(.a(G278), .O(gate49inter8));
  nand2 gate920(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate921(.a(s_53), .b(gate49inter3), .O(gate49inter10));
  nor2  gate922(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate923(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate924(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1275(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1276(.a(gate56inter0), .b(s_104), .O(gate56inter1));
  and2  gate1277(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1278(.a(s_104), .O(gate56inter3));
  inv1  gate1279(.a(s_105), .O(gate56inter4));
  nand2 gate1280(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1281(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1282(.a(G16), .O(gate56inter7));
  inv1  gate1283(.a(G287), .O(gate56inter8));
  nand2 gate1284(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1285(.a(s_105), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1286(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1287(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1288(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate631(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate632(.a(gate58inter0), .b(s_12), .O(gate58inter1));
  and2  gate633(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate634(.a(s_12), .O(gate58inter3));
  inv1  gate635(.a(s_13), .O(gate58inter4));
  nand2 gate636(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate637(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate638(.a(G18), .O(gate58inter7));
  inv1  gate639(.a(G290), .O(gate58inter8));
  nand2 gate640(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate641(.a(s_13), .b(gate58inter3), .O(gate58inter10));
  nor2  gate642(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate643(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate644(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate743(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate744(.a(gate63inter0), .b(s_28), .O(gate63inter1));
  and2  gate745(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate746(.a(s_28), .O(gate63inter3));
  inv1  gate747(.a(s_29), .O(gate63inter4));
  nand2 gate748(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate749(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate750(.a(G23), .O(gate63inter7));
  inv1  gate751(.a(G299), .O(gate63inter8));
  nand2 gate752(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate753(.a(s_29), .b(gate63inter3), .O(gate63inter10));
  nor2  gate754(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate755(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate756(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate855(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate856(.a(gate72inter0), .b(s_44), .O(gate72inter1));
  and2  gate857(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate858(.a(s_44), .O(gate72inter3));
  inv1  gate859(.a(s_45), .O(gate72inter4));
  nand2 gate860(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate861(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate862(.a(G32), .O(gate72inter7));
  inv1  gate863(.a(G311), .O(gate72inter8));
  nand2 gate864(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate865(.a(s_45), .b(gate72inter3), .O(gate72inter10));
  nor2  gate866(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate867(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate868(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1065(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1066(.a(gate77inter0), .b(s_74), .O(gate77inter1));
  and2  gate1067(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1068(.a(s_74), .O(gate77inter3));
  inv1  gate1069(.a(s_75), .O(gate77inter4));
  nand2 gate1070(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1071(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1072(.a(G2), .O(gate77inter7));
  inv1  gate1073(.a(G320), .O(gate77inter8));
  nand2 gate1074(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1075(.a(s_75), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1076(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1077(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1078(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate757(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate758(.a(gate79inter0), .b(s_30), .O(gate79inter1));
  and2  gate759(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate760(.a(s_30), .O(gate79inter3));
  inv1  gate761(.a(s_31), .O(gate79inter4));
  nand2 gate762(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate763(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate764(.a(G10), .O(gate79inter7));
  inv1  gate765(.a(G323), .O(gate79inter8));
  nand2 gate766(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate767(.a(s_31), .b(gate79inter3), .O(gate79inter10));
  nor2  gate768(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate769(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate770(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1177(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1178(.a(gate84inter0), .b(s_90), .O(gate84inter1));
  and2  gate1179(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1180(.a(s_90), .O(gate84inter3));
  inv1  gate1181(.a(s_91), .O(gate84inter4));
  nand2 gate1182(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1183(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1184(.a(G15), .O(gate84inter7));
  inv1  gate1185(.a(G329), .O(gate84inter8));
  nand2 gate1186(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1187(.a(s_91), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1188(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1189(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1190(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate869(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate870(.a(gate86inter0), .b(s_46), .O(gate86inter1));
  and2  gate871(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate872(.a(s_46), .O(gate86inter3));
  inv1  gate873(.a(s_47), .O(gate86inter4));
  nand2 gate874(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate875(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate876(.a(G8), .O(gate86inter7));
  inv1  gate877(.a(G332), .O(gate86inter8));
  nand2 gate878(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate879(.a(s_47), .b(gate86inter3), .O(gate86inter10));
  nor2  gate880(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate881(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate882(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1205(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1206(.a(gate98inter0), .b(s_94), .O(gate98inter1));
  and2  gate1207(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1208(.a(s_94), .O(gate98inter3));
  inv1  gate1209(.a(s_95), .O(gate98inter4));
  nand2 gate1210(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1211(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1212(.a(G23), .O(gate98inter7));
  inv1  gate1213(.a(G350), .O(gate98inter8));
  nand2 gate1214(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1215(.a(s_95), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1216(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1217(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1218(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1149(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1150(.a(gate99inter0), .b(s_86), .O(gate99inter1));
  and2  gate1151(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1152(.a(s_86), .O(gate99inter3));
  inv1  gate1153(.a(s_87), .O(gate99inter4));
  nand2 gate1154(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1155(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1156(.a(G27), .O(gate99inter7));
  inv1  gate1157(.a(G353), .O(gate99inter8));
  nand2 gate1158(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1159(.a(s_87), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1160(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1161(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1162(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate645(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate646(.a(gate101inter0), .b(s_14), .O(gate101inter1));
  and2  gate647(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate648(.a(s_14), .O(gate101inter3));
  inv1  gate649(.a(s_15), .O(gate101inter4));
  nand2 gate650(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate651(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate652(.a(G20), .O(gate101inter7));
  inv1  gate653(.a(G356), .O(gate101inter8));
  nand2 gate654(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate655(.a(s_15), .b(gate101inter3), .O(gate101inter10));
  nor2  gate656(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate657(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate658(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1415(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1416(.a(gate108inter0), .b(s_124), .O(gate108inter1));
  and2  gate1417(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1418(.a(s_124), .O(gate108inter3));
  inv1  gate1419(.a(s_125), .O(gate108inter4));
  nand2 gate1420(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1421(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1422(.a(G368), .O(gate108inter7));
  inv1  gate1423(.a(G369), .O(gate108inter8));
  nand2 gate1424(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1425(.a(s_125), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1426(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1427(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1428(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1429(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1430(.a(gate113inter0), .b(s_126), .O(gate113inter1));
  and2  gate1431(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1432(.a(s_126), .O(gate113inter3));
  inv1  gate1433(.a(s_127), .O(gate113inter4));
  nand2 gate1434(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1435(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1436(.a(G378), .O(gate113inter7));
  inv1  gate1437(.a(G379), .O(gate113inter8));
  nand2 gate1438(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1439(.a(s_127), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1440(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1441(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1442(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate659(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate660(.a(gate130inter0), .b(s_16), .O(gate130inter1));
  and2  gate661(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate662(.a(s_16), .O(gate130inter3));
  inv1  gate663(.a(s_17), .O(gate130inter4));
  nand2 gate664(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate665(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate666(.a(G412), .O(gate130inter7));
  inv1  gate667(.a(G413), .O(gate130inter8));
  nand2 gate668(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate669(.a(s_17), .b(gate130inter3), .O(gate130inter10));
  nor2  gate670(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate671(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate672(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate715(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate716(.a(gate133inter0), .b(s_24), .O(gate133inter1));
  and2  gate717(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate718(.a(s_24), .O(gate133inter3));
  inv1  gate719(.a(s_25), .O(gate133inter4));
  nand2 gate720(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate721(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate722(.a(G418), .O(gate133inter7));
  inv1  gate723(.a(G419), .O(gate133inter8));
  nand2 gate724(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate725(.a(s_25), .b(gate133inter3), .O(gate133inter10));
  nor2  gate726(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate727(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate728(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate813(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate814(.a(gate134inter0), .b(s_38), .O(gate134inter1));
  and2  gate815(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate816(.a(s_38), .O(gate134inter3));
  inv1  gate817(.a(s_39), .O(gate134inter4));
  nand2 gate818(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate819(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate820(.a(G420), .O(gate134inter7));
  inv1  gate821(.a(G421), .O(gate134inter8));
  nand2 gate822(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate823(.a(s_39), .b(gate134inter3), .O(gate134inter10));
  nor2  gate824(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate825(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate826(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate547(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate548(.a(gate150inter0), .b(s_0), .O(gate150inter1));
  and2  gate549(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate550(.a(s_0), .O(gate150inter3));
  inv1  gate551(.a(s_1), .O(gate150inter4));
  nand2 gate552(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate553(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate554(.a(G504), .O(gate150inter7));
  inv1  gate555(.a(G507), .O(gate150inter8));
  nand2 gate556(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate557(.a(s_1), .b(gate150inter3), .O(gate150inter10));
  nor2  gate558(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate559(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate560(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate673(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate674(.a(gate160inter0), .b(s_18), .O(gate160inter1));
  and2  gate675(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate676(.a(s_18), .O(gate160inter3));
  inv1  gate677(.a(s_19), .O(gate160inter4));
  nand2 gate678(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate679(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate680(.a(G447), .O(gate160inter7));
  inv1  gate681(.a(G531), .O(gate160inter8));
  nand2 gate682(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate683(.a(s_19), .b(gate160inter3), .O(gate160inter10));
  nor2  gate684(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate685(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate686(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate967(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate968(.a(gate161inter0), .b(s_60), .O(gate161inter1));
  and2  gate969(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate970(.a(s_60), .O(gate161inter3));
  inv1  gate971(.a(s_61), .O(gate161inter4));
  nand2 gate972(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate973(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate974(.a(G450), .O(gate161inter7));
  inv1  gate975(.a(G534), .O(gate161inter8));
  nand2 gate976(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate977(.a(s_61), .b(gate161inter3), .O(gate161inter10));
  nor2  gate978(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate979(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate980(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1107(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1108(.a(gate162inter0), .b(s_80), .O(gate162inter1));
  and2  gate1109(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1110(.a(s_80), .O(gate162inter3));
  inv1  gate1111(.a(s_81), .O(gate162inter4));
  nand2 gate1112(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1113(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1114(.a(G453), .O(gate162inter7));
  inv1  gate1115(.a(G534), .O(gate162inter8));
  nand2 gate1116(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1117(.a(s_81), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1118(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1119(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1120(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1359(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1360(.a(gate170inter0), .b(s_116), .O(gate170inter1));
  and2  gate1361(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1362(.a(s_116), .O(gate170inter3));
  inv1  gate1363(.a(s_117), .O(gate170inter4));
  nand2 gate1364(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1365(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1366(.a(G477), .O(gate170inter7));
  inv1  gate1367(.a(G546), .O(gate170inter8));
  nand2 gate1368(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1369(.a(s_117), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1370(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1371(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1372(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate561(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate562(.a(gate183inter0), .b(s_2), .O(gate183inter1));
  and2  gate563(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate564(.a(s_2), .O(gate183inter3));
  inv1  gate565(.a(s_3), .O(gate183inter4));
  nand2 gate566(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate567(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate568(.a(G516), .O(gate183inter7));
  inv1  gate569(.a(G567), .O(gate183inter8));
  nand2 gate570(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate571(.a(s_3), .b(gate183inter3), .O(gate183inter10));
  nor2  gate572(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate573(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate574(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate701(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate702(.a(gate188inter0), .b(s_22), .O(gate188inter1));
  and2  gate703(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate704(.a(s_22), .O(gate188inter3));
  inv1  gate705(.a(s_23), .O(gate188inter4));
  nand2 gate706(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate707(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate708(.a(G576), .O(gate188inter7));
  inv1  gate709(.a(G577), .O(gate188inter8));
  nand2 gate710(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate711(.a(s_23), .b(gate188inter3), .O(gate188inter10));
  nor2  gate712(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate713(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate714(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate925(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate926(.a(gate190inter0), .b(s_54), .O(gate190inter1));
  and2  gate927(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate928(.a(s_54), .O(gate190inter3));
  inv1  gate929(.a(s_55), .O(gate190inter4));
  nand2 gate930(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate931(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate932(.a(G580), .O(gate190inter7));
  inv1  gate933(.a(G581), .O(gate190inter8));
  nand2 gate934(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate935(.a(s_55), .b(gate190inter3), .O(gate190inter10));
  nor2  gate936(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate937(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate938(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1135(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1136(.a(gate195inter0), .b(s_84), .O(gate195inter1));
  and2  gate1137(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1138(.a(s_84), .O(gate195inter3));
  inv1  gate1139(.a(s_85), .O(gate195inter4));
  nand2 gate1140(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1141(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1142(.a(G590), .O(gate195inter7));
  inv1  gate1143(.a(G591), .O(gate195inter8));
  nand2 gate1144(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1145(.a(s_85), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1146(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1147(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1148(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate827(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate828(.a(gate196inter0), .b(s_40), .O(gate196inter1));
  and2  gate829(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate830(.a(s_40), .O(gate196inter3));
  inv1  gate831(.a(s_41), .O(gate196inter4));
  nand2 gate832(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate833(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate834(.a(G592), .O(gate196inter7));
  inv1  gate835(.a(G593), .O(gate196inter8));
  nand2 gate836(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate837(.a(s_41), .b(gate196inter3), .O(gate196inter10));
  nor2  gate838(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate839(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate840(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1079(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1080(.a(gate202inter0), .b(s_76), .O(gate202inter1));
  and2  gate1081(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1082(.a(s_76), .O(gate202inter3));
  inv1  gate1083(.a(s_77), .O(gate202inter4));
  nand2 gate1084(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1085(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1086(.a(G612), .O(gate202inter7));
  inv1  gate1087(.a(G617), .O(gate202inter8));
  nand2 gate1088(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1089(.a(s_77), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1090(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1091(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1092(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1457(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1458(.a(gate205inter0), .b(s_130), .O(gate205inter1));
  and2  gate1459(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1460(.a(s_130), .O(gate205inter3));
  inv1  gate1461(.a(s_131), .O(gate205inter4));
  nand2 gate1462(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1463(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1464(.a(G622), .O(gate205inter7));
  inv1  gate1465(.a(G627), .O(gate205inter8));
  nand2 gate1466(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1467(.a(s_131), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1468(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1469(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1470(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1051(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1052(.a(gate213inter0), .b(s_72), .O(gate213inter1));
  and2  gate1053(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1054(.a(s_72), .O(gate213inter3));
  inv1  gate1055(.a(s_73), .O(gate213inter4));
  nand2 gate1056(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1057(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1058(.a(G602), .O(gate213inter7));
  inv1  gate1059(.a(G672), .O(gate213inter8));
  nand2 gate1060(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1061(.a(s_73), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1062(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1063(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1064(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1093(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1094(.a(gate216inter0), .b(s_78), .O(gate216inter1));
  and2  gate1095(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1096(.a(s_78), .O(gate216inter3));
  inv1  gate1097(.a(s_79), .O(gate216inter4));
  nand2 gate1098(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1099(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1100(.a(G617), .O(gate216inter7));
  inv1  gate1101(.a(G675), .O(gate216inter8));
  nand2 gate1102(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1103(.a(s_79), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1104(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1105(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1106(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1037(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1038(.a(gate227inter0), .b(s_70), .O(gate227inter1));
  and2  gate1039(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1040(.a(s_70), .O(gate227inter3));
  inv1  gate1041(.a(s_71), .O(gate227inter4));
  nand2 gate1042(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1043(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1044(.a(G694), .O(gate227inter7));
  inv1  gate1045(.a(G695), .O(gate227inter8));
  nand2 gate1046(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1047(.a(s_71), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1048(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1049(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1050(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1191(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1192(.a(gate247inter0), .b(s_92), .O(gate247inter1));
  and2  gate1193(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1194(.a(s_92), .O(gate247inter3));
  inv1  gate1195(.a(s_93), .O(gate247inter4));
  nand2 gate1196(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1197(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1198(.a(G251), .O(gate247inter7));
  inv1  gate1199(.a(G739), .O(gate247inter8));
  nand2 gate1200(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1201(.a(s_93), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1202(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1203(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1204(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate995(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate996(.a(gate248inter0), .b(s_64), .O(gate248inter1));
  and2  gate997(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate998(.a(s_64), .O(gate248inter3));
  inv1  gate999(.a(s_65), .O(gate248inter4));
  nand2 gate1000(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1001(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1002(.a(G727), .O(gate248inter7));
  inv1  gate1003(.a(G739), .O(gate248inter8));
  nand2 gate1004(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1005(.a(s_65), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1006(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1007(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1008(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate841(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate842(.a(gate254inter0), .b(s_42), .O(gate254inter1));
  and2  gate843(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate844(.a(s_42), .O(gate254inter3));
  inv1  gate845(.a(s_43), .O(gate254inter4));
  nand2 gate846(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate847(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate848(.a(G712), .O(gate254inter7));
  inv1  gate849(.a(G748), .O(gate254inter8));
  nand2 gate850(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate851(.a(s_43), .b(gate254inter3), .O(gate254inter10));
  nor2  gate852(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate853(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate854(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1331(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1332(.a(gate259inter0), .b(s_112), .O(gate259inter1));
  and2  gate1333(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1334(.a(s_112), .O(gate259inter3));
  inv1  gate1335(.a(s_113), .O(gate259inter4));
  nand2 gate1336(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1337(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1338(.a(G758), .O(gate259inter7));
  inv1  gate1339(.a(G759), .O(gate259inter8));
  nand2 gate1340(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1341(.a(s_113), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1342(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1343(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1344(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate617(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate618(.a(gate272inter0), .b(s_10), .O(gate272inter1));
  and2  gate619(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate620(.a(s_10), .O(gate272inter3));
  inv1  gate621(.a(s_11), .O(gate272inter4));
  nand2 gate622(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate623(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate624(.a(G663), .O(gate272inter7));
  inv1  gate625(.a(G791), .O(gate272inter8));
  nand2 gate626(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate627(.a(s_11), .b(gate272inter3), .O(gate272inter10));
  nor2  gate628(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate629(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate630(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate771(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate772(.a(gate276inter0), .b(s_32), .O(gate276inter1));
  and2  gate773(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate774(.a(s_32), .O(gate276inter3));
  inv1  gate775(.a(s_33), .O(gate276inter4));
  nand2 gate776(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate777(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate778(.a(G773), .O(gate276inter7));
  inv1  gate779(.a(G797), .O(gate276inter8));
  nand2 gate780(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate781(.a(s_33), .b(gate276inter3), .O(gate276inter10));
  nor2  gate782(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate783(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate784(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate785(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate786(.a(gate282inter0), .b(s_34), .O(gate282inter1));
  and2  gate787(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate788(.a(s_34), .O(gate282inter3));
  inv1  gate789(.a(s_35), .O(gate282inter4));
  nand2 gate790(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate791(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate792(.a(G782), .O(gate282inter7));
  inv1  gate793(.a(G806), .O(gate282inter8));
  nand2 gate794(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate795(.a(s_35), .b(gate282inter3), .O(gate282inter10));
  nor2  gate796(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate797(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate798(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate603(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate604(.a(gate287inter0), .b(s_8), .O(gate287inter1));
  and2  gate605(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate606(.a(s_8), .O(gate287inter3));
  inv1  gate607(.a(s_9), .O(gate287inter4));
  nand2 gate608(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate609(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate610(.a(G663), .O(gate287inter7));
  inv1  gate611(.a(G815), .O(gate287inter8));
  nand2 gate612(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate613(.a(s_9), .b(gate287inter3), .O(gate287inter10));
  nor2  gate614(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate615(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate616(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1121(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1122(.a(gate401inter0), .b(s_82), .O(gate401inter1));
  and2  gate1123(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1124(.a(s_82), .O(gate401inter3));
  inv1  gate1125(.a(s_83), .O(gate401inter4));
  nand2 gate1126(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1127(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1128(.a(G15), .O(gate401inter7));
  inv1  gate1129(.a(G1078), .O(gate401inter8));
  nand2 gate1130(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1131(.a(s_83), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1132(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1133(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1134(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1401(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1402(.a(gate406inter0), .b(s_122), .O(gate406inter1));
  and2  gate1403(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1404(.a(s_122), .O(gate406inter3));
  inv1  gate1405(.a(s_123), .O(gate406inter4));
  nand2 gate1406(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1407(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1408(.a(G20), .O(gate406inter7));
  inv1  gate1409(.a(G1093), .O(gate406inter8));
  nand2 gate1410(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1411(.a(s_123), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1412(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1413(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1414(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate981(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate982(.a(gate415inter0), .b(s_62), .O(gate415inter1));
  and2  gate983(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate984(.a(s_62), .O(gate415inter3));
  inv1  gate985(.a(s_63), .O(gate415inter4));
  nand2 gate986(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate987(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate988(.a(G29), .O(gate415inter7));
  inv1  gate989(.a(G1120), .O(gate415inter8));
  nand2 gate990(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate991(.a(s_63), .b(gate415inter3), .O(gate415inter10));
  nor2  gate992(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate993(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate994(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate883(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate884(.a(gate417inter0), .b(s_48), .O(gate417inter1));
  and2  gate885(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate886(.a(s_48), .O(gate417inter3));
  inv1  gate887(.a(s_49), .O(gate417inter4));
  nand2 gate888(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate889(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate890(.a(G31), .O(gate417inter7));
  inv1  gate891(.a(G1126), .O(gate417inter8));
  nand2 gate892(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate893(.a(s_49), .b(gate417inter3), .O(gate417inter10));
  nor2  gate894(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate895(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate896(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1373(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1374(.a(gate420inter0), .b(s_118), .O(gate420inter1));
  and2  gate1375(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1376(.a(s_118), .O(gate420inter3));
  inv1  gate1377(.a(s_119), .O(gate420inter4));
  nand2 gate1378(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1379(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1380(.a(G1036), .O(gate420inter7));
  inv1  gate1381(.a(G1132), .O(gate420inter8));
  nand2 gate1382(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1383(.a(s_119), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1384(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1385(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1386(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate687(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate688(.a(gate425inter0), .b(s_20), .O(gate425inter1));
  and2  gate689(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate690(.a(s_20), .O(gate425inter3));
  inv1  gate691(.a(s_21), .O(gate425inter4));
  nand2 gate692(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate693(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate694(.a(G4), .O(gate425inter7));
  inv1  gate695(.a(G1141), .O(gate425inter8));
  nand2 gate696(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate697(.a(s_21), .b(gate425inter3), .O(gate425inter10));
  nor2  gate698(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate699(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate700(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate939(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate940(.a(gate426inter0), .b(s_56), .O(gate426inter1));
  and2  gate941(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate942(.a(s_56), .O(gate426inter3));
  inv1  gate943(.a(s_57), .O(gate426inter4));
  nand2 gate944(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate945(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate946(.a(G1045), .O(gate426inter7));
  inv1  gate947(.a(G1141), .O(gate426inter8));
  nand2 gate948(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate949(.a(s_57), .b(gate426inter3), .O(gate426inter10));
  nor2  gate950(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate951(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate952(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1233(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1234(.a(gate431inter0), .b(s_98), .O(gate431inter1));
  and2  gate1235(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1236(.a(s_98), .O(gate431inter3));
  inv1  gate1237(.a(s_99), .O(gate431inter4));
  nand2 gate1238(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1239(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1240(.a(G7), .O(gate431inter7));
  inv1  gate1241(.a(G1150), .O(gate431inter8));
  nand2 gate1242(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1243(.a(s_99), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1244(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1245(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1246(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1261(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1262(.a(gate432inter0), .b(s_102), .O(gate432inter1));
  and2  gate1263(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1264(.a(s_102), .O(gate432inter3));
  inv1  gate1265(.a(s_103), .O(gate432inter4));
  nand2 gate1266(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1267(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1268(.a(G1054), .O(gate432inter7));
  inv1  gate1269(.a(G1150), .O(gate432inter8));
  nand2 gate1270(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1271(.a(s_103), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1272(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1273(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1274(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1443(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1444(.a(gate435inter0), .b(s_128), .O(gate435inter1));
  and2  gate1445(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1446(.a(s_128), .O(gate435inter3));
  inv1  gate1447(.a(s_129), .O(gate435inter4));
  nand2 gate1448(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1449(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1450(.a(G9), .O(gate435inter7));
  inv1  gate1451(.a(G1156), .O(gate435inter8));
  nand2 gate1452(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1453(.a(s_129), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1454(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1455(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1456(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1317(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1318(.a(gate437inter0), .b(s_110), .O(gate437inter1));
  and2  gate1319(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1320(.a(s_110), .O(gate437inter3));
  inv1  gate1321(.a(s_111), .O(gate437inter4));
  nand2 gate1322(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1323(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1324(.a(G10), .O(gate437inter7));
  inv1  gate1325(.a(G1159), .O(gate437inter8));
  nand2 gate1326(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1327(.a(s_111), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1328(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1329(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1330(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1219(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1220(.a(gate438inter0), .b(s_96), .O(gate438inter1));
  and2  gate1221(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1222(.a(s_96), .O(gate438inter3));
  inv1  gate1223(.a(s_97), .O(gate438inter4));
  nand2 gate1224(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1225(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1226(.a(G1063), .O(gate438inter7));
  inv1  gate1227(.a(G1159), .O(gate438inter8));
  nand2 gate1228(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1229(.a(s_97), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1230(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1231(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1232(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1345(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1346(.a(gate441inter0), .b(s_114), .O(gate441inter1));
  and2  gate1347(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1348(.a(s_114), .O(gate441inter3));
  inv1  gate1349(.a(s_115), .O(gate441inter4));
  nand2 gate1350(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1351(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1352(.a(G12), .O(gate441inter7));
  inv1  gate1353(.a(G1165), .O(gate441inter8));
  nand2 gate1354(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1355(.a(s_115), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1356(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1357(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1358(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1289(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1290(.a(gate444inter0), .b(s_106), .O(gate444inter1));
  and2  gate1291(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1292(.a(s_106), .O(gate444inter3));
  inv1  gate1293(.a(s_107), .O(gate444inter4));
  nand2 gate1294(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1295(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1296(.a(G1072), .O(gate444inter7));
  inv1  gate1297(.a(G1168), .O(gate444inter8));
  nand2 gate1298(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1299(.a(s_107), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1300(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1301(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1302(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1247(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1248(.a(gate450inter0), .b(s_100), .O(gate450inter1));
  and2  gate1249(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1250(.a(s_100), .O(gate450inter3));
  inv1  gate1251(.a(s_101), .O(gate450inter4));
  nand2 gate1252(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1253(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1254(.a(G1081), .O(gate450inter7));
  inv1  gate1255(.a(G1177), .O(gate450inter8));
  nand2 gate1256(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1257(.a(s_101), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1258(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1259(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1260(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1303(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1304(.a(gate456inter0), .b(s_108), .O(gate456inter1));
  and2  gate1305(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1306(.a(s_108), .O(gate456inter3));
  inv1  gate1307(.a(s_109), .O(gate456inter4));
  nand2 gate1308(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1309(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1310(.a(G1090), .O(gate456inter7));
  inv1  gate1311(.a(G1186), .O(gate456inter8));
  nand2 gate1312(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1313(.a(s_109), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1314(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1315(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1316(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate799(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate800(.a(gate460inter0), .b(s_36), .O(gate460inter1));
  and2  gate801(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate802(.a(s_36), .O(gate460inter3));
  inv1  gate803(.a(s_37), .O(gate460inter4));
  nand2 gate804(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate805(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate806(.a(G1096), .O(gate460inter7));
  inv1  gate807(.a(G1192), .O(gate460inter8));
  nand2 gate808(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate809(.a(s_37), .b(gate460inter3), .O(gate460inter10));
  nor2  gate810(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate811(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate812(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1009(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1010(.a(gate466inter0), .b(s_66), .O(gate466inter1));
  and2  gate1011(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1012(.a(s_66), .O(gate466inter3));
  inv1  gate1013(.a(s_67), .O(gate466inter4));
  nand2 gate1014(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1015(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1016(.a(G1105), .O(gate466inter7));
  inv1  gate1017(.a(G1201), .O(gate466inter8));
  nand2 gate1018(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1019(.a(s_67), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1020(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1021(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1022(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate729(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate730(.a(gate476inter0), .b(s_26), .O(gate476inter1));
  and2  gate731(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate732(.a(s_26), .O(gate476inter3));
  inv1  gate733(.a(s_27), .O(gate476inter4));
  nand2 gate734(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate735(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate736(.a(G1120), .O(gate476inter7));
  inv1  gate737(.a(G1216), .O(gate476inter8));
  nand2 gate738(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate739(.a(s_27), .b(gate476inter3), .O(gate476inter10));
  nor2  gate740(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate741(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate742(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate953(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate954(.a(gate488inter0), .b(s_58), .O(gate488inter1));
  and2  gate955(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate956(.a(s_58), .O(gate488inter3));
  inv1  gate957(.a(s_59), .O(gate488inter4));
  nand2 gate958(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate959(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate960(.a(G1238), .O(gate488inter7));
  inv1  gate961(.a(G1239), .O(gate488inter8));
  nand2 gate962(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate963(.a(s_59), .b(gate488inter3), .O(gate488inter10));
  nor2  gate964(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate965(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate966(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1023(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1024(.a(gate491inter0), .b(s_68), .O(gate491inter1));
  and2  gate1025(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1026(.a(s_68), .O(gate491inter3));
  inv1  gate1027(.a(s_69), .O(gate491inter4));
  nand2 gate1028(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1029(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1030(.a(G1244), .O(gate491inter7));
  inv1  gate1031(.a(G1245), .O(gate491inter8));
  nand2 gate1032(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1033(.a(s_69), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1034(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1035(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1036(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate897(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate898(.a(gate499inter0), .b(s_50), .O(gate499inter1));
  and2  gate899(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate900(.a(s_50), .O(gate499inter3));
  inv1  gate901(.a(s_51), .O(gate499inter4));
  nand2 gate902(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate903(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate904(.a(G1260), .O(gate499inter7));
  inv1  gate905(.a(G1261), .O(gate499inter8));
  nand2 gate906(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate907(.a(s_51), .b(gate499inter3), .O(gate499inter10));
  nor2  gate908(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate909(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate910(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1163(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1164(.a(gate510inter0), .b(s_88), .O(gate510inter1));
  and2  gate1165(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1166(.a(s_88), .O(gate510inter3));
  inv1  gate1167(.a(s_89), .O(gate510inter4));
  nand2 gate1168(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1169(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1170(.a(G1282), .O(gate510inter7));
  inv1  gate1171(.a(G1283), .O(gate510inter8));
  nand2 gate1172(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1173(.a(s_89), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1174(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1175(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1176(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule