module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate687(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate688(.a(gate11inter0), .b(s_20), .O(gate11inter1));
  and2  gate689(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate690(.a(s_20), .O(gate11inter3));
  inv1  gate691(.a(s_21), .O(gate11inter4));
  nand2 gate692(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate693(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate694(.a(G5), .O(gate11inter7));
  inv1  gate695(.a(G6), .O(gate11inter8));
  nand2 gate696(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate697(.a(s_21), .b(gate11inter3), .O(gate11inter10));
  nor2  gate698(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate699(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate700(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate715(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate716(.a(gate12inter0), .b(s_24), .O(gate12inter1));
  and2  gate717(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate718(.a(s_24), .O(gate12inter3));
  inv1  gate719(.a(s_25), .O(gate12inter4));
  nand2 gate720(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate721(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate722(.a(G7), .O(gate12inter7));
  inv1  gate723(.a(G8), .O(gate12inter8));
  nand2 gate724(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate725(.a(s_25), .b(gate12inter3), .O(gate12inter10));
  nor2  gate726(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate727(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate728(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate939(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate940(.a(gate22inter0), .b(s_56), .O(gate22inter1));
  and2  gate941(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate942(.a(s_56), .O(gate22inter3));
  inv1  gate943(.a(s_57), .O(gate22inter4));
  nand2 gate944(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate945(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate946(.a(G27), .O(gate22inter7));
  inv1  gate947(.a(G28), .O(gate22inter8));
  nand2 gate948(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate949(.a(s_57), .b(gate22inter3), .O(gate22inter10));
  nor2  gate950(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate951(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate952(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate799(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate800(.a(gate25inter0), .b(s_36), .O(gate25inter1));
  and2  gate801(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate802(.a(s_36), .O(gate25inter3));
  inv1  gate803(.a(s_37), .O(gate25inter4));
  nand2 gate804(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate805(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate806(.a(G1), .O(gate25inter7));
  inv1  gate807(.a(G5), .O(gate25inter8));
  nand2 gate808(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate809(.a(s_37), .b(gate25inter3), .O(gate25inter10));
  nor2  gate810(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate811(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate812(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1079(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1080(.a(gate26inter0), .b(s_76), .O(gate26inter1));
  and2  gate1081(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1082(.a(s_76), .O(gate26inter3));
  inv1  gate1083(.a(s_77), .O(gate26inter4));
  nand2 gate1084(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1085(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1086(.a(G9), .O(gate26inter7));
  inv1  gate1087(.a(G13), .O(gate26inter8));
  nand2 gate1088(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1089(.a(s_77), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1090(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1091(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1092(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1009(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1010(.a(gate31inter0), .b(s_66), .O(gate31inter1));
  and2  gate1011(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1012(.a(s_66), .O(gate31inter3));
  inv1  gate1013(.a(s_67), .O(gate31inter4));
  nand2 gate1014(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1015(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1016(.a(G4), .O(gate31inter7));
  inv1  gate1017(.a(G8), .O(gate31inter8));
  nand2 gate1018(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1019(.a(s_67), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1020(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1021(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1022(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1345(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1346(.a(gate54inter0), .b(s_114), .O(gate54inter1));
  and2  gate1347(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1348(.a(s_114), .O(gate54inter3));
  inv1  gate1349(.a(s_115), .O(gate54inter4));
  nand2 gate1350(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1351(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1352(.a(G14), .O(gate54inter7));
  inv1  gate1353(.a(G284), .O(gate54inter8));
  nand2 gate1354(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1355(.a(s_115), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1356(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1357(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1358(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1177(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1178(.a(gate55inter0), .b(s_90), .O(gate55inter1));
  and2  gate1179(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1180(.a(s_90), .O(gate55inter3));
  inv1  gate1181(.a(s_91), .O(gate55inter4));
  nand2 gate1182(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1183(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1184(.a(G15), .O(gate55inter7));
  inv1  gate1185(.a(G287), .O(gate55inter8));
  nand2 gate1186(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1187(.a(s_91), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1188(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1189(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1190(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate967(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate968(.a(gate60inter0), .b(s_60), .O(gate60inter1));
  and2  gate969(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate970(.a(s_60), .O(gate60inter3));
  inv1  gate971(.a(s_61), .O(gate60inter4));
  nand2 gate972(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate973(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate974(.a(G20), .O(gate60inter7));
  inv1  gate975(.a(G293), .O(gate60inter8));
  nand2 gate976(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate977(.a(s_61), .b(gate60inter3), .O(gate60inter10));
  nor2  gate978(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate979(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate980(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1275(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1276(.a(gate61inter0), .b(s_104), .O(gate61inter1));
  and2  gate1277(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1278(.a(s_104), .O(gate61inter3));
  inv1  gate1279(.a(s_105), .O(gate61inter4));
  nand2 gate1280(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1281(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1282(.a(G21), .O(gate61inter7));
  inv1  gate1283(.a(G296), .O(gate61inter8));
  nand2 gate1284(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1285(.a(s_105), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1286(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1287(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1288(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate897(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate898(.a(gate65inter0), .b(s_50), .O(gate65inter1));
  and2  gate899(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate900(.a(s_50), .O(gate65inter3));
  inv1  gate901(.a(s_51), .O(gate65inter4));
  nand2 gate902(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate903(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate904(.a(G25), .O(gate65inter7));
  inv1  gate905(.a(G302), .O(gate65inter8));
  nand2 gate906(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate907(.a(s_51), .b(gate65inter3), .O(gate65inter10));
  nor2  gate908(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate909(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate910(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1093(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1094(.a(gate68inter0), .b(s_78), .O(gate68inter1));
  and2  gate1095(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1096(.a(s_78), .O(gate68inter3));
  inv1  gate1097(.a(s_79), .O(gate68inter4));
  nand2 gate1098(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1099(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1100(.a(G28), .O(gate68inter7));
  inv1  gate1101(.a(G305), .O(gate68inter8));
  nand2 gate1102(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1103(.a(s_79), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1104(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1105(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1106(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate841(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate842(.a(gate76inter0), .b(s_42), .O(gate76inter1));
  and2  gate843(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate844(.a(s_42), .O(gate76inter3));
  inv1  gate845(.a(s_43), .O(gate76inter4));
  nand2 gate846(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate847(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate848(.a(G13), .O(gate76inter7));
  inv1  gate849(.a(G317), .O(gate76inter8));
  nand2 gate850(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate851(.a(s_43), .b(gate76inter3), .O(gate76inter10));
  nor2  gate852(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate853(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate854(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1247(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1248(.a(gate98inter0), .b(s_100), .O(gate98inter1));
  and2  gate1249(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1250(.a(s_100), .O(gate98inter3));
  inv1  gate1251(.a(s_101), .O(gate98inter4));
  nand2 gate1252(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1253(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1254(.a(G23), .O(gate98inter7));
  inv1  gate1255(.a(G350), .O(gate98inter8));
  nand2 gate1256(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1257(.a(s_101), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1258(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1259(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1260(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1303(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1304(.a(gate103inter0), .b(s_108), .O(gate103inter1));
  and2  gate1305(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1306(.a(s_108), .O(gate103inter3));
  inv1  gate1307(.a(s_109), .O(gate103inter4));
  nand2 gate1308(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1309(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1310(.a(G28), .O(gate103inter7));
  inv1  gate1311(.a(G359), .O(gate103inter8));
  nand2 gate1312(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1313(.a(s_109), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1314(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1315(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1316(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate953(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate954(.a(gate120inter0), .b(s_58), .O(gate120inter1));
  and2  gate955(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate956(.a(s_58), .O(gate120inter3));
  inv1  gate957(.a(s_59), .O(gate120inter4));
  nand2 gate958(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate959(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate960(.a(G392), .O(gate120inter7));
  inv1  gate961(.a(G393), .O(gate120inter8));
  nand2 gate962(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate963(.a(s_59), .b(gate120inter3), .O(gate120inter10));
  nor2  gate964(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate965(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate966(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1163(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1164(.a(gate123inter0), .b(s_88), .O(gate123inter1));
  and2  gate1165(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1166(.a(s_88), .O(gate123inter3));
  inv1  gate1167(.a(s_89), .O(gate123inter4));
  nand2 gate1168(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1169(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1170(.a(G398), .O(gate123inter7));
  inv1  gate1171(.a(G399), .O(gate123inter8));
  nand2 gate1172(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1173(.a(s_89), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1174(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1175(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1176(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate925(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate926(.a(gate128inter0), .b(s_54), .O(gate128inter1));
  and2  gate927(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate928(.a(s_54), .O(gate128inter3));
  inv1  gate929(.a(s_55), .O(gate128inter4));
  nand2 gate930(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate931(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate932(.a(G408), .O(gate128inter7));
  inv1  gate933(.a(G409), .O(gate128inter8));
  nand2 gate934(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate935(.a(s_55), .b(gate128inter3), .O(gate128inter10));
  nor2  gate936(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate937(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate938(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate869(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate870(.a(gate141inter0), .b(s_46), .O(gate141inter1));
  and2  gate871(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate872(.a(s_46), .O(gate141inter3));
  inv1  gate873(.a(s_47), .O(gate141inter4));
  nand2 gate874(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate875(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate876(.a(G450), .O(gate141inter7));
  inv1  gate877(.a(G453), .O(gate141inter8));
  nand2 gate878(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate879(.a(s_47), .b(gate141inter3), .O(gate141inter10));
  nor2  gate880(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate881(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate882(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1191(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1192(.a(gate144inter0), .b(s_92), .O(gate144inter1));
  and2  gate1193(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1194(.a(s_92), .O(gate144inter3));
  inv1  gate1195(.a(s_93), .O(gate144inter4));
  nand2 gate1196(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1197(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1198(.a(G468), .O(gate144inter7));
  inv1  gate1199(.a(G471), .O(gate144inter8));
  nand2 gate1200(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1201(.a(s_93), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1202(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1203(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1204(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate995(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate996(.a(gate150inter0), .b(s_64), .O(gate150inter1));
  and2  gate997(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate998(.a(s_64), .O(gate150inter3));
  inv1  gate999(.a(s_65), .O(gate150inter4));
  nand2 gate1000(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1001(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1002(.a(G504), .O(gate150inter7));
  inv1  gate1003(.a(G507), .O(gate150inter8));
  nand2 gate1004(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1005(.a(s_65), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1006(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1007(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1008(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate645(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate646(.a(gate153inter0), .b(s_14), .O(gate153inter1));
  and2  gate647(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate648(.a(s_14), .O(gate153inter3));
  inv1  gate649(.a(s_15), .O(gate153inter4));
  nand2 gate650(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate651(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate652(.a(G426), .O(gate153inter7));
  inv1  gate653(.a(G522), .O(gate153inter8));
  nand2 gate654(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate655(.a(s_15), .b(gate153inter3), .O(gate153inter10));
  nor2  gate656(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate657(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate658(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate827(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate828(.a(gate154inter0), .b(s_40), .O(gate154inter1));
  and2  gate829(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate830(.a(s_40), .O(gate154inter3));
  inv1  gate831(.a(s_41), .O(gate154inter4));
  nand2 gate832(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate833(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate834(.a(G429), .O(gate154inter7));
  inv1  gate835(.a(G522), .O(gate154inter8));
  nand2 gate836(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate837(.a(s_41), .b(gate154inter3), .O(gate154inter10));
  nor2  gate838(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate839(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate840(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate771(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate772(.a(gate162inter0), .b(s_32), .O(gate162inter1));
  and2  gate773(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate774(.a(s_32), .O(gate162inter3));
  inv1  gate775(.a(s_33), .O(gate162inter4));
  nand2 gate776(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate777(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate778(.a(G453), .O(gate162inter7));
  inv1  gate779(.a(G534), .O(gate162inter8));
  nand2 gate780(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate781(.a(s_33), .b(gate162inter3), .O(gate162inter10));
  nor2  gate782(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate783(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate784(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate729(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate730(.a(gate164inter0), .b(s_26), .O(gate164inter1));
  and2  gate731(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate732(.a(s_26), .O(gate164inter3));
  inv1  gate733(.a(s_27), .O(gate164inter4));
  nand2 gate734(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate735(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate736(.a(G459), .O(gate164inter7));
  inv1  gate737(.a(G537), .O(gate164inter8));
  nand2 gate738(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate739(.a(s_27), .b(gate164inter3), .O(gate164inter10));
  nor2  gate740(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate741(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate742(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1219(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1220(.a(gate169inter0), .b(s_96), .O(gate169inter1));
  and2  gate1221(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1222(.a(s_96), .O(gate169inter3));
  inv1  gate1223(.a(s_97), .O(gate169inter4));
  nand2 gate1224(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1225(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1226(.a(G474), .O(gate169inter7));
  inv1  gate1227(.a(G546), .O(gate169inter8));
  nand2 gate1228(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1229(.a(s_97), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1230(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1231(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1232(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1121(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1122(.a(gate179inter0), .b(s_82), .O(gate179inter1));
  and2  gate1123(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1124(.a(s_82), .O(gate179inter3));
  inv1  gate1125(.a(s_83), .O(gate179inter4));
  nand2 gate1126(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1127(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1128(.a(G504), .O(gate179inter7));
  inv1  gate1129(.a(G561), .O(gate179inter8));
  nand2 gate1130(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1131(.a(s_83), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1132(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1133(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1134(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate659(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate660(.a(gate181inter0), .b(s_16), .O(gate181inter1));
  and2  gate661(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate662(.a(s_16), .O(gate181inter3));
  inv1  gate663(.a(s_17), .O(gate181inter4));
  nand2 gate664(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate665(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate666(.a(G510), .O(gate181inter7));
  inv1  gate667(.a(G564), .O(gate181inter8));
  nand2 gate668(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate669(.a(s_17), .b(gate181inter3), .O(gate181inter10));
  nor2  gate670(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate671(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate672(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1317(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1318(.a(gate184inter0), .b(s_110), .O(gate184inter1));
  and2  gate1319(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1320(.a(s_110), .O(gate184inter3));
  inv1  gate1321(.a(s_111), .O(gate184inter4));
  nand2 gate1322(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1323(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1324(.a(G519), .O(gate184inter7));
  inv1  gate1325(.a(G567), .O(gate184inter8));
  nand2 gate1326(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1327(.a(s_111), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1328(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1329(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1330(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1289(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1290(.a(gate188inter0), .b(s_106), .O(gate188inter1));
  and2  gate1291(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1292(.a(s_106), .O(gate188inter3));
  inv1  gate1293(.a(s_107), .O(gate188inter4));
  nand2 gate1294(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1295(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1296(.a(G576), .O(gate188inter7));
  inv1  gate1297(.a(G577), .O(gate188inter8));
  nand2 gate1298(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1299(.a(s_107), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1300(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1301(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1302(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1037(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1038(.a(gate222inter0), .b(s_70), .O(gate222inter1));
  and2  gate1039(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1040(.a(s_70), .O(gate222inter3));
  inv1  gate1041(.a(s_71), .O(gate222inter4));
  nand2 gate1042(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1043(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1044(.a(G632), .O(gate222inter7));
  inv1  gate1045(.a(G684), .O(gate222inter8));
  nand2 gate1046(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1047(.a(s_71), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1048(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1049(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1050(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1149(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1150(.a(gate225inter0), .b(s_86), .O(gate225inter1));
  and2  gate1151(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1152(.a(s_86), .O(gate225inter3));
  inv1  gate1153(.a(s_87), .O(gate225inter4));
  nand2 gate1154(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1155(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1156(.a(G690), .O(gate225inter7));
  inv1  gate1157(.a(G691), .O(gate225inter8));
  nand2 gate1158(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1159(.a(s_87), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1160(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1161(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1162(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1023(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1024(.a(gate228inter0), .b(s_68), .O(gate228inter1));
  and2  gate1025(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1026(.a(s_68), .O(gate228inter3));
  inv1  gate1027(.a(s_69), .O(gate228inter4));
  nand2 gate1028(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1029(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1030(.a(G696), .O(gate228inter7));
  inv1  gate1031(.a(G697), .O(gate228inter8));
  nand2 gate1032(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1033(.a(s_69), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1034(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1035(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1036(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate813(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate814(.a(gate229inter0), .b(s_38), .O(gate229inter1));
  and2  gate815(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate816(.a(s_38), .O(gate229inter3));
  inv1  gate817(.a(s_39), .O(gate229inter4));
  nand2 gate818(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate819(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate820(.a(G698), .O(gate229inter7));
  inv1  gate821(.a(G699), .O(gate229inter8));
  nand2 gate822(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate823(.a(s_39), .b(gate229inter3), .O(gate229inter10));
  nor2  gate824(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate825(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate826(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1107(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1108(.a(gate231inter0), .b(s_80), .O(gate231inter1));
  and2  gate1109(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1110(.a(s_80), .O(gate231inter3));
  inv1  gate1111(.a(s_81), .O(gate231inter4));
  nand2 gate1112(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1113(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1114(.a(G702), .O(gate231inter7));
  inv1  gate1115(.a(G703), .O(gate231inter8));
  nand2 gate1116(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1117(.a(s_81), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1118(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1119(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1120(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate757(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate758(.a(gate256inter0), .b(s_30), .O(gate256inter1));
  and2  gate759(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate760(.a(s_30), .O(gate256inter3));
  inv1  gate761(.a(s_31), .O(gate256inter4));
  nand2 gate762(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate763(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate764(.a(G715), .O(gate256inter7));
  inv1  gate765(.a(G751), .O(gate256inter8));
  nand2 gate766(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate767(.a(s_31), .b(gate256inter3), .O(gate256inter10));
  nor2  gate768(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate769(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate770(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate701(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate702(.a(gate258inter0), .b(s_22), .O(gate258inter1));
  and2  gate703(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate704(.a(s_22), .O(gate258inter3));
  inv1  gate705(.a(s_23), .O(gate258inter4));
  nand2 gate706(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate707(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate708(.a(G756), .O(gate258inter7));
  inv1  gate709(.a(G757), .O(gate258inter8));
  nand2 gate710(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate711(.a(s_23), .b(gate258inter3), .O(gate258inter10));
  nor2  gate712(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate713(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate714(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1051(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1052(.a(gate259inter0), .b(s_72), .O(gate259inter1));
  and2  gate1053(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1054(.a(s_72), .O(gate259inter3));
  inv1  gate1055(.a(s_73), .O(gate259inter4));
  nand2 gate1056(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1057(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1058(.a(G758), .O(gate259inter7));
  inv1  gate1059(.a(G759), .O(gate259inter8));
  nand2 gate1060(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1061(.a(s_73), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1062(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1063(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1064(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate561(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate562(.a(gate260inter0), .b(s_2), .O(gate260inter1));
  and2  gate563(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate564(.a(s_2), .O(gate260inter3));
  inv1  gate565(.a(s_3), .O(gate260inter4));
  nand2 gate566(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate567(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate568(.a(G760), .O(gate260inter7));
  inv1  gate569(.a(G761), .O(gate260inter8));
  nand2 gate570(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate571(.a(s_3), .b(gate260inter3), .O(gate260inter10));
  nor2  gate572(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate573(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate574(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1261(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1262(.a(gate266inter0), .b(s_102), .O(gate266inter1));
  and2  gate1263(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1264(.a(s_102), .O(gate266inter3));
  inv1  gate1265(.a(s_103), .O(gate266inter4));
  nand2 gate1266(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1267(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1268(.a(G645), .O(gate266inter7));
  inv1  gate1269(.a(G773), .O(gate266inter8));
  nand2 gate1270(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1271(.a(s_103), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1272(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1273(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1274(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate855(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate856(.a(gate270inter0), .b(s_44), .O(gate270inter1));
  and2  gate857(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate858(.a(s_44), .O(gate270inter3));
  inv1  gate859(.a(s_45), .O(gate270inter4));
  nand2 gate860(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate861(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate862(.a(G657), .O(gate270inter7));
  inv1  gate863(.a(G785), .O(gate270inter8));
  nand2 gate864(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate865(.a(s_45), .b(gate270inter3), .O(gate270inter10));
  nor2  gate866(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate867(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate868(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate743(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate744(.a(gate271inter0), .b(s_28), .O(gate271inter1));
  and2  gate745(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate746(.a(s_28), .O(gate271inter3));
  inv1  gate747(.a(s_29), .O(gate271inter4));
  nand2 gate748(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate749(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate750(.a(G660), .O(gate271inter7));
  inv1  gate751(.a(G788), .O(gate271inter8));
  nand2 gate752(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate753(.a(s_29), .b(gate271inter3), .O(gate271inter10));
  nor2  gate754(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate755(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate756(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1359(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1360(.a(gate281inter0), .b(s_116), .O(gate281inter1));
  and2  gate1361(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1362(.a(s_116), .O(gate281inter3));
  inv1  gate1363(.a(s_117), .O(gate281inter4));
  nand2 gate1364(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1365(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1366(.a(G654), .O(gate281inter7));
  inv1  gate1367(.a(G806), .O(gate281inter8));
  nand2 gate1368(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1369(.a(s_117), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1370(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1371(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1372(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1065(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1066(.a(gate294inter0), .b(s_74), .O(gate294inter1));
  and2  gate1067(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1068(.a(s_74), .O(gate294inter3));
  inv1  gate1069(.a(s_75), .O(gate294inter4));
  nand2 gate1070(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1071(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1072(.a(G832), .O(gate294inter7));
  inv1  gate1073(.a(G833), .O(gate294inter8));
  nand2 gate1074(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1075(.a(s_75), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1076(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1077(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1078(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate547(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate548(.a(gate387inter0), .b(s_0), .O(gate387inter1));
  and2  gate549(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate550(.a(s_0), .O(gate387inter3));
  inv1  gate551(.a(s_1), .O(gate387inter4));
  nand2 gate552(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate553(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate554(.a(G1), .O(gate387inter7));
  inv1  gate555(.a(G1036), .O(gate387inter8));
  nand2 gate556(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate557(.a(s_1), .b(gate387inter3), .O(gate387inter10));
  nor2  gate558(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate559(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate560(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate981(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate982(.a(gate392inter0), .b(s_62), .O(gate392inter1));
  and2  gate983(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate984(.a(s_62), .O(gate392inter3));
  inv1  gate985(.a(s_63), .O(gate392inter4));
  nand2 gate986(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate987(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate988(.a(G6), .O(gate392inter7));
  inv1  gate989(.a(G1051), .O(gate392inter8));
  nand2 gate990(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate991(.a(s_63), .b(gate392inter3), .O(gate392inter10));
  nor2  gate992(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate993(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate994(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate617(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate618(.a(gate395inter0), .b(s_10), .O(gate395inter1));
  and2  gate619(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate620(.a(s_10), .O(gate395inter3));
  inv1  gate621(.a(s_11), .O(gate395inter4));
  nand2 gate622(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate623(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate624(.a(G9), .O(gate395inter7));
  inv1  gate625(.a(G1060), .O(gate395inter8));
  nand2 gate626(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate627(.a(s_11), .b(gate395inter3), .O(gate395inter10));
  nor2  gate628(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate629(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate630(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate673(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate674(.a(gate418inter0), .b(s_18), .O(gate418inter1));
  and2  gate675(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate676(.a(s_18), .O(gate418inter3));
  inv1  gate677(.a(s_19), .O(gate418inter4));
  nand2 gate678(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate679(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate680(.a(G32), .O(gate418inter7));
  inv1  gate681(.a(G1129), .O(gate418inter8));
  nand2 gate682(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate683(.a(s_19), .b(gate418inter3), .O(gate418inter10));
  nor2  gate684(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate685(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate686(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1135(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1136(.a(gate421inter0), .b(s_84), .O(gate421inter1));
  and2  gate1137(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1138(.a(s_84), .O(gate421inter3));
  inv1  gate1139(.a(s_85), .O(gate421inter4));
  nand2 gate1140(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1141(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1142(.a(G2), .O(gate421inter7));
  inv1  gate1143(.a(G1135), .O(gate421inter8));
  nand2 gate1144(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1145(.a(s_85), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1146(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1147(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1148(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate631(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate632(.a(gate456inter0), .b(s_12), .O(gate456inter1));
  and2  gate633(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate634(.a(s_12), .O(gate456inter3));
  inv1  gate635(.a(s_13), .O(gate456inter4));
  nand2 gate636(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate637(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate638(.a(G1090), .O(gate456inter7));
  inv1  gate639(.a(G1186), .O(gate456inter8));
  nand2 gate640(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate641(.a(s_13), .b(gate456inter3), .O(gate456inter10));
  nor2  gate642(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate643(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate644(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1387(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1388(.a(gate461inter0), .b(s_120), .O(gate461inter1));
  and2  gate1389(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1390(.a(s_120), .O(gate461inter3));
  inv1  gate1391(.a(s_121), .O(gate461inter4));
  nand2 gate1392(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1393(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1394(.a(G22), .O(gate461inter7));
  inv1  gate1395(.a(G1195), .O(gate461inter8));
  nand2 gate1396(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1397(.a(s_121), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1398(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1399(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1400(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1233(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1234(.a(gate472inter0), .b(s_98), .O(gate472inter1));
  and2  gate1235(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1236(.a(s_98), .O(gate472inter3));
  inv1  gate1237(.a(s_99), .O(gate472inter4));
  nand2 gate1238(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1239(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1240(.a(G1114), .O(gate472inter7));
  inv1  gate1241(.a(G1210), .O(gate472inter8));
  nand2 gate1242(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1243(.a(s_99), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1244(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1245(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1246(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate883(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate884(.a(gate478inter0), .b(s_48), .O(gate478inter1));
  and2  gate885(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate886(.a(s_48), .O(gate478inter3));
  inv1  gate887(.a(s_49), .O(gate478inter4));
  nand2 gate888(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate889(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate890(.a(G1123), .O(gate478inter7));
  inv1  gate891(.a(G1219), .O(gate478inter8));
  nand2 gate892(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate893(.a(s_49), .b(gate478inter3), .O(gate478inter10));
  nor2  gate894(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate895(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate896(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate589(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate590(.a(gate482inter0), .b(s_6), .O(gate482inter1));
  and2  gate591(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate592(.a(s_6), .O(gate482inter3));
  inv1  gate593(.a(s_7), .O(gate482inter4));
  nand2 gate594(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate595(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate596(.a(G1129), .O(gate482inter7));
  inv1  gate597(.a(G1225), .O(gate482inter8));
  nand2 gate598(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate599(.a(s_7), .b(gate482inter3), .O(gate482inter10));
  nor2  gate600(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate601(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate602(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1373(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1374(.a(gate484inter0), .b(s_118), .O(gate484inter1));
  and2  gate1375(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1376(.a(s_118), .O(gate484inter3));
  inv1  gate1377(.a(s_119), .O(gate484inter4));
  nand2 gate1378(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1379(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1380(.a(G1230), .O(gate484inter7));
  inv1  gate1381(.a(G1231), .O(gate484inter8));
  nand2 gate1382(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1383(.a(s_119), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1384(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1385(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1386(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1331(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1332(.a(gate487inter0), .b(s_112), .O(gate487inter1));
  and2  gate1333(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1334(.a(s_112), .O(gate487inter3));
  inv1  gate1335(.a(s_113), .O(gate487inter4));
  nand2 gate1336(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1337(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1338(.a(G1236), .O(gate487inter7));
  inv1  gate1339(.a(G1237), .O(gate487inter8));
  nand2 gate1340(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1341(.a(s_113), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1342(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1343(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1344(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate785(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate786(.a(gate493inter0), .b(s_34), .O(gate493inter1));
  and2  gate787(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate788(.a(s_34), .O(gate493inter3));
  inv1  gate789(.a(s_35), .O(gate493inter4));
  nand2 gate790(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate791(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate792(.a(G1248), .O(gate493inter7));
  inv1  gate793(.a(G1249), .O(gate493inter8));
  nand2 gate794(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate795(.a(s_35), .b(gate493inter3), .O(gate493inter10));
  nor2  gate796(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate797(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate798(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1205(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1206(.a(gate495inter0), .b(s_94), .O(gate495inter1));
  and2  gate1207(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1208(.a(s_94), .O(gate495inter3));
  inv1  gate1209(.a(s_95), .O(gate495inter4));
  nand2 gate1210(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1211(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1212(.a(G1252), .O(gate495inter7));
  inv1  gate1213(.a(G1253), .O(gate495inter8));
  nand2 gate1214(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1215(.a(s_95), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1216(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1217(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1218(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate575(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate576(.a(gate497inter0), .b(s_4), .O(gate497inter1));
  and2  gate577(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate578(.a(s_4), .O(gate497inter3));
  inv1  gate579(.a(s_5), .O(gate497inter4));
  nand2 gate580(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate581(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate582(.a(G1256), .O(gate497inter7));
  inv1  gate583(.a(G1257), .O(gate497inter8));
  nand2 gate584(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate585(.a(s_5), .b(gate497inter3), .O(gate497inter10));
  nor2  gate586(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate587(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate588(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate603(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate604(.a(gate499inter0), .b(s_8), .O(gate499inter1));
  and2  gate605(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate606(.a(s_8), .O(gate499inter3));
  inv1  gate607(.a(s_9), .O(gate499inter4));
  nand2 gate608(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate609(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate610(.a(G1260), .O(gate499inter7));
  inv1  gate611(.a(G1261), .O(gate499inter8));
  nand2 gate612(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate613(.a(s_9), .b(gate499inter3), .O(gate499inter10));
  nor2  gate614(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate615(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate616(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate911(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate912(.a(gate501inter0), .b(s_52), .O(gate501inter1));
  and2  gate913(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate914(.a(s_52), .O(gate501inter3));
  inv1  gate915(.a(s_53), .O(gate501inter4));
  nand2 gate916(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate917(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate918(.a(G1264), .O(gate501inter7));
  inv1  gate919(.a(G1265), .O(gate501inter8));
  nand2 gate920(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate921(.a(s_53), .b(gate501inter3), .O(gate501inter10));
  nor2  gate922(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate923(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate924(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule