module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1807(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1808(.a(gate16inter0), .b(s_180), .O(gate16inter1));
  and2  gate1809(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1810(.a(s_180), .O(gate16inter3));
  inv1  gate1811(.a(s_181), .O(gate16inter4));
  nand2 gate1812(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1813(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1814(.a(G15), .O(gate16inter7));
  inv1  gate1815(.a(G16), .O(gate16inter8));
  nand2 gate1816(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1817(.a(s_181), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1818(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1819(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1820(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1611(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1612(.a(gate18inter0), .b(s_152), .O(gate18inter1));
  and2  gate1613(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1614(.a(s_152), .O(gate18inter3));
  inv1  gate1615(.a(s_153), .O(gate18inter4));
  nand2 gate1616(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1617(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1618(.a(G19), .O(gate18inter7));
  inv1  gate1619(.a(G20), .O(gate18inter8));
  nand2 gate1620(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1621(.a(s_153), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1622(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1623(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1624(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate701(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate702(.a(gate19inter0), .b(s_22), .O(gate19inter1));
  and2  gate703(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate704(.a(s_22), .O(gate19inter3));
  inv1  gate705(.a(s_23), .O(gate19inter4));
  nand2 gate706(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate707(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate708(.a(G21), .O(gate19inter7));
  inv1  gate709(.a(G22), .O(gate19inter8));
  nand2 gate710(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate711(.a(s_23), .b(gate19inter3), .O(gate19inter10));
  nor2  gate712(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate713(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate714(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1625(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1626(.a(gate21inter0), .b(s_154), .O(gate21inter1));
  and2  gate1627(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1628(.a(s_154), .O(gate21inter3));
  inv1  gate1629(.a(s_155), .O(gate21inter4));
  nand2 gate1630(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1631(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1632(.a(G25), .O(gate21inter7));
  inv1  gate1633(.a(G26), .O(gate21inter8));
  nand2 gate1634(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1635(.a(s_155), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1636(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1637(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1638(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1569(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1570(.a(gate22inter0), .b(s_146), .O(gate22inter1));
  and2  gate1571(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1572(.a(s_146), .O(gate22inter3));
  inv1  gate1573(.a(s_147), .O(gate22inter4));
  nand2 gate1574(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1575(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1576(.a(G27), .O(gate22inter7));
  inv1  gate1577(.a(G28), .O(gate22inter8));
  nand2 gate1578(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1579(.a(s_147), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1580(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1581(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1582(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1121(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1122(.a(gate24inter0), .b(s_82), .O(gate24inter1));
  and2  gate1123(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1124(.a(s_82), .O(gate24inter3));
  inv1  gate1125(.a(s_83), .O(gate24inter4));
  nand2 gate1126(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1127(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1128(.a(G31), .O(gate24inter7));
  inv1  gate1129(.a(G32), .O(gate24inter8));
  nand2 gate1130(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1131(.a(s_83), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1132(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1133(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1134(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate659(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate660(.a(gate30inter0), .b(s_16), .O(gate30inter1));
  and2  gate661(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate662(.a(s_16), .O(gate30inter3));
  inv1  gate663(.a(s_17), .O(gate30inter4));
  nand2 gate664(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate665(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate666(.a(G11), .O(gate30inter7));
  inv1  gate667(.a(G15), .O(gate30inter8));
  nand2 gate668(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate669(.a(s_17), .b(gate30inter3), .O(gate30inter10));
  nor2  gate670(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate671(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate672(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1401(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1402(.a(gate32inter0), .b(s_122), .O(gate32inter1));
  and2  gate1403(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1404(.a(s_122), .O(gate32inter3));
  inv1  gate1405(.a(s_123), .O(gate32inter4));
  nand2 gate1406(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1407(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1408(.a(G12), .O(gate32inter7));
  inv1  gate1409(.a(G16), .O(gate32inter8));
  nand2 gate1410(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1411(.a(s_123), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1412(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1413(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1414(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1779(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1780(.a(gate35inter0), .b(s_176), .O(gate35inter1));
  and2  gate1781(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1782(.a(s_176), .O(gate35inter3));
  inv1  gate1783(.a(s_177), .O(gate35inter4));
  nand2 gate1784(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1785(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1786(.a(G18), .O(gate35inter7));
  inv1  gate1787(.a(G22), .O(gate35inter8));
  nand2 gate1788(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1789(.a(s_177), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1790(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1791(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1792(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1835(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1836(.a(gate37inter0), .b(s_184), .O(gate37inter1));
  and2  gate1837(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1838(.a(s_184), .O(gate37inter3));
  inv1  gate1839(.a(s_185), .O(gate37inter4));
  nand2 gate1840(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1841(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1842(.a(G19), .O(gate37inter7));
  inv1  gate1843(.a(G23), .O(gate37inter8));
  nand2 gate1844(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1845(.a(s_185), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1846(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1847(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1848(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate841(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate842(.a(gate41inter0), .b(s_42), .O(gate41inter1));
  and2  gate843(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate844(.a(s_42), .O(gate41inter3));
  inv1  gate845(.a(s_43), .O(gate41inter4));
  nand2 gate846(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate847(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate848(.a(G1), .O(gate41inter7));
  inv1  gate849(.a(G266), .O(gate41inter8));
  nand2 gate850(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate851(.a(s_43), .b(gate41inter3), .O(gate41inter10));
  nor2  gate852(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate853(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate854(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1681(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1682(.a(gate43inter0), .b(s_162), .O(gate43inter1));
  and2  gate1683(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1684(.a(s_162), .O(gate43inter3));
  inv1  gate1685(.a(s_163), .O(gate43inter4));
  nand2 gate1686(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1687(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1688(.a(G3), .O(gate43inter7));
  inv1  gate1689(.a(G269), .O(gate43inter8));
  nand2 gate1690(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1691(.a(s_163), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1692(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1693(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1694(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate911(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate912(.a(gate44inter0), .b(s_52), .O(gate44inter1));
  and2  gate913(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate914(.a(s_52), .O(gate44inter3));
  inv1  gate915(.a(s_53), .O(gate44inter4));
  nand2 gate916(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate917(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate918(.a(G4), .O(gate44inter7));
  inv1  gate919(.a(G269), .O(gate44inter8));
  nand2 gate920(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate921(.a(s_53), .b(gate44inter3), .O(gate44inter10));
  nor2  gate922(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate923(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate924(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1289(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1290(.a(gate45inter0), .b(s_106), .O(gate45inter1));
  and2  gate1291(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1292(.a(s_106), .O(gate45inter3));
  inv1  gate1293(.a(s_107), .O(gate45inter4));
  nand2 gate1294(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1295(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1296(.a(G5), .O(gate45inter7));
  inv1  gate1297(.a(G272), .O(gate45inter8));
  nand2 gate1298(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1299(.a(s_107), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1300(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1301(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1302(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1233(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1234(.a(gate46inter0), .b(s_98), .O(gate46inter1));
  and2  gate1235(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1236(.a(s_98), .O(gate46inter3));
  inv1  gate1237(.a(s_99), .O(gate46inter4));
  nand2 gate1238(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1239(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1240(.a(G6), .O(gate46inter7));
  inv1  gate1241(.a(G272), .O(gate46inter8));
  nand2 gate1242(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1243(.a(s_99), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1244(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1245(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1246(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1555(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1556(.a(gate54inter0), .b(s_144), .O(gate54inter1));
  and2  gate1557(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1558(.a(s_144), .O(gate54inter3));
  inv1  gate1559(.a(s_145), .O(gate54inter4));
  nand2 gate1560(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1561(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1562(.a(G14), .O(gate54inter7));
  inv1  gate1563(.a(G284), .O(gate54inter8));
  nand2 gate1564(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1565(.a(s_145), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1566(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1567(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1568(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1821(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1822(.a(gate61inter0), .b(s_182), .O(gate61inter1));
  and2  gate1823(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1824(.a(s_182), .O(gate61inter3));
  inv1  gate1825(.a(s_183), .O(gate61inter4));
  nand2 gate1826(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1827(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1828(.a(G21), .O(gate61inter7));
  inv1  gate1829(.a(G296), .O(gate61inter8));
  nand2 gate1830(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1831(.a(s_183), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1832(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1833(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1834(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1695(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1696(.a(gate63inter0), .b(s_164), .O(gate63inter1));
  and2  gate1697(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1698(.a(s_164), .O(gate63inter3));
  inv1  gate1699(.a(s_165), .O(gate63inter4));
  nand2 gate1700(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1701(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1702(.a(G23), .O(gate63inter7));
  inv1  gate1703(.a(G299), .O(gate63inter8));
  nand2 gate1704(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1705(.a(s_165), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1706(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1707(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1708(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate981(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate982(.a(gate72inter0), .b(s_62), .O(gate72inter1));
  and2  gate983(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate984(.a(s_62), .O(gate72inter3));
  inv1  gate985(.a(s_63), .O(gate72inter4));
  nand2 gate986(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate987(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate988(.a(G32), .O(gate72inter7));
  inv1  gate989(.a(G311), .O(gate72inter8));
  nand2 gate990(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate991(.a(s_63), .b(gate72inter3), .O(gate72inter10));
  nor2  gate992(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate993(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate994(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate589(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate590(.a(gate74inter0), .b(s_6), .O(gate74inter1));
  and2  gate591(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate592(.a(s_6), .O(gate74inter3));
  inv1  gate593(.a(s_7), .O(gate74inter4));
  nand2 gate594(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate595(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate596(.a(G5), .O(gate74inter7));
  inv1  gate597(.a(G314), .O(gate74inter8));
  nand2 gate598(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate599(.a(s_7), .b(gate74inter3), .O(gate74inter10));
  nor2  gate600(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate601(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate602(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1485(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1486(.a(gate76inter0), .b(s_134), .O(gate76inter1));
  and2  gate1487(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1488(.a(s_134), .O(gate76inter3));
  inv1  gate1489(.a(s_135), .O(gate76inter4));
  nand2 gate1490(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1491(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1492(.a(G13), .O(gate76inter7));
  inv1  gate1493(.a(G317), .O(gate76inter8));
  nand2 gate1494(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1495(.a(s_135), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1496(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1497(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1498(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1051(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1052(.a(gate85inter0), .b(s_72), .O(gate85inter1));
  and2  gate1053(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1054(.a(s_72), .O(gate85inter3));
  inv1  gate1055(.a(s_73), .O(gate85inter4));
  nand2 gate1056(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1057(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1058(.a(G4), .O(gate85inter7));
  inv1  gate1059(.a(G332), .O(gate85inter8));
  nand2 gate1060(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1061(.a(s_73), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1062(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1063(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1064(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1723(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1724(.a(gate90inter0), .b(s_168), .O(gate90inter1));
  and2  gate1725(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1726(.a(s_168), .O(gate90inter3));
  inv1  gate1727(.a(s_169), .O(gate90inter4));
  nand2 gate1728(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1729(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1730(.a(G21), .O(gate90inter7));
  inv1  gate1731(.a(G338), .O(gate90inter8));
  nand2 gate1732(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1733(.a(s_169), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1734(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1735(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1736(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1751(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1752(.a(gate92inter0), .b(s_172), .O(gate92inter1));
  and2  gate1753(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1754(.a(s_172), .O(gate92inter3));
  inv1  gate1755(.a(s_173), .O(gate92inter4));
  nand2 gate1756(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1757(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1758(.a(G29), .O(gate92inter7));
  inv1  gate1759(.a(G341), .O(gate92inter8));
  nand2 gate1760(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1761(.a(s_173), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1762(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1763(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1764(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1457(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1458(.a(gate93inter0), .b(s_130), .O(gate93inter1));
  and2  gate1459(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1460(.a(s_130), .O(gate93inter3));
  inv1  gate1461(.a(s_131), .O(gate93inter4));
  nand2 gate1462(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1463(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1464(.a(G18), .O(gate93inter7));
  inv1  gate1465(.a(G344), .O(gate93inter8));
  nand2 gate1466(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1467(.a(s_131), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1468(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1469(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1470(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1037(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1038(.a(gate97inter0), .b(s_70), .O(gate97inter1));
  and2  gate1039(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1040(.a(s_70), .O(gate97inter3));
  inv1  gate1041(.a(s_71), .O(gate97inter4));
  nand2 gate1042(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1043(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1044(.a(G19), .O(gate97inter7));
  inv1  gate1045(.a(G350), .O(gate97inter8));
  nand2 gate1046(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1047(.a(s_71), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1048(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1049(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1050(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1653(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1654(.a(gate101inter0), .b(s_158), .O(gate101inter1));
  and2  gate1655(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1656(.a(s_158), .O(gate101inter3));
  inv1  gate1657(.a(s_159), .O(gate101inter4));
  nand2 gate1658(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1659(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1660(.a(G20), .O(gate101inter7));
  inv1  gate1661(.a(G356), .O(gate101inter8));
  nand2 gate1662(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1663(.a(s_159), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1664(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1665(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1666(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1737(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1738(.a(gate104inter0), .b(s_170), .O(gate104inter1));
  and2  gate1739(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1740(.a(s_170), .O(gate104inter3));
  inv1  gate1741(.a(s_171), .O(gate104inter4));
  nand2 gate1742(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1743(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1744(.a(G32), .O(gate104inter7));
  inv1  gate1745(.a(G359), .O(gate104inter8));
  nand2 gate1746(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1747(.a(s_171), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1748(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1749(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1750(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1317(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1318(.a(gate106inter0), .b(s_110), .O(gate106inter1));
  and2  gate1319(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1320(.a(s_110), .O(gate106inter3));
  inv1  gate1321(.a(s_111), .O(gate106inter4));
  nand2 gate1322(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1323(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1324(.a(G364), .O(gate106inter7));
  inv1  gate1325(.a(G365), .O(gate106inter8));
  nand2 gate1326(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1327(.a(s_111), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1328(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1329(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1330(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1177(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1178(.a(gate109inter0), .b(s_90), .O(gate109inter1));
  and2  gate1179(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1180(.a(s_90), .O(gate109inter3));
  inv1  gate1181(.a(s_91), .O(gate109inter4));
  nand2 gate1182(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1183(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1184(.a(G370), .O(gate109inter7));
  inv1  gate1185(.a(G371), .O(gate109inter8));
  nand2 gate1186(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1187(.a(s_91), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1188(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1189(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1190(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate757(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate758(.a(gate116inter0), .b(s_30), .O(gate116inter1));
  and2  gate759(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate760(.a(s_30), .O(gate116inter3));
  inv1  gate761(.a(s_31), .O(gate116inter4));
  nand2 gate762(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate763(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate764(.a(G384), .O(gate116inter7));
  inv1  gate765(.a(G385), .O(gate116inter8));
  nand2 gate766(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate767(.a(s_31), .b(gate116inter3), .O(gate116inter10));
  nor2  gate768(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate769(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate770(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1373(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1374(.a(gate117inter0), .b(s_118), .O(gate117inter1));
  and2  gate1375(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1376(.a(s_118), .O(gate117inter3));
  inv1  gate1377(.a(s_119), .O(gate117inter4));
  nand2 gate1378(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1379(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1380(.a(G386), .O(gate117inter7));
  inv1  gate1381(.a(G387), .O(gate117inter8));
  nand2 gate1382(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1383(.a(s_119), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1384(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1385(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1386(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate953(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate954(.a(gate123inter0), .b(s_58), .O(gate123inter1));
  and2  gate955(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate956(.a(s_58), .O(gate123inter3));
  inv1  gate957(.a(s_59), .O(gate123inter4));
  nand2 gate958(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate959(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate960(.a(G398), .O(gate123inter7));
  inv1  gate961(.a(G399), .O(gate123inter8));
  nand2 gate962(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate963(.a(s_59), .b(gate123inter3), .O(gate123inter10));
  nor2  gate964(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate965(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate966(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1107(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1108(.a(gate125inter0), .b(s_80), .O(gate125inter1));
  and2  gate1109(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1110(.a(s_80), .O(gate125inter3));
  inv1  gate1111(.a(s_81), .O(gate125inter4));
  nand2 gate1112(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1113(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1114(.a(G402), .O(gate125inter7));
  inv1  gate1115(.a(G403), .O(gate125inter8));
  nand2 gate1116(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1117(.a(s_81), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1118(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1119(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1120(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1065(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1066(.a(gate126inter0), .b(s_74), .O(gate126inter1));
  and2  gate1067(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1068(.a(s_74), .O(gate126inter3));
  inv1  gate1069(.a(s_75), .O(gate126inter4));
  nand2 gate1070(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1071(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1072(.a(G404), .O(gate126inter7));
  inv1  gate1073(.a(G405), .O(gate126inter8));
  nand2 gate1074(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1075(.a(s_75), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1076(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1077(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1078(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1499(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1500(.a(gate128inter0), .b(s_136), .O(gate128inter1));
  and2  gate1501(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1502(.a(s_136), .O(gate128inter3));
  inv1  gate1503(.a(s_137), .O(gate128inter4));
  nand2 gate1504(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1505(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1506(.a(G408), .O(gate128inter7));
  inv1  gate1507(.a(G409), .O(gate128inter8));
  nand2 gate1508(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1509(.a(s_137), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1510(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1511(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1512(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1639(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1640(.a(gate129inter0), .b(s_156), .O(gate129inter1));
  and2  gate1641(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1642(.a(s_156), .O(gate129inter3));
  inv1  gate1643(.a(s_157), .O(gate129inter4));
  nand2 gate1644(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1645(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1646(.a(G410), .O(gate129inter7));
  inv1  gate1647(.a(G411), .O(gate129inter8));
  nand2 gate1648(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1649(.a(s_157), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1650(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1651(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1652(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate715(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate716(.a(gate131inter0), .b(s_24), .O(gate131inter1));
  and2  gate717(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate718(.a(s_24), .O(gate131inter3));
  inv1  gate719(.a(s_25), .O(gate131inter4));
  nand2 gate720(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate721(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate722(.a(G414), .O(gate131inter7));
  inv1  gate723(.a(G415), .O(gate131inter8));
  nand2 gate724(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate725(.a(s_25), .b(gate131inter3), .O(gate131inter10));
  nor2  gate726(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate727(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate728(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1429(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1430(.a(gate137inter0), .b(s_126), .O(gate137inter1));
  and2  gate1431(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1432(.a(s_126), .O(gate137inter3));
  inv1  gate1433(.a(s_127), .O(gate137inter4));
  nand2 gate1434(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1435(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1436(.a(G426), .O(gate137inter7));
  inv1  gate1437(.a(G429), .O(gate137inter8));
  nand2 gate1438(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1439(.a(s_127), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1440(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1441(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1442(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate925(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate926(.a(gate141inter0), .b(s_54), .O(gate141inter1));
  and2  gate927(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate928(.a(s_54), .O(gate141inter3));
  inv1  gate929(.a(s_55), .O(gate141inter4));
  nand2 gate930(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate931(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate932(.a(G450), .O(gate141inter7));
  inv1  gate933(.a(G453), .O(gate141inter8));
  nand2 gate934(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate935(.a(s_55), .b(gate141inter3), .O(gate141inter10));
  nor2  gate936(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate937(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate938(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate939(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate940(.a(gate146inter0), .b(s_56), .O(gate146inter1));
  and2  gate941(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate942(.a(s_56), .O(gate146inter3));
  inv1  gate943(.a(s_57), .O(gate146inter4));
  nand2 gate944(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate945(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate946(.a(G480), .O(gate146inter7));
  inv1  gate947(.a(G483), .O(gate146inter8));
  nand2 gate948(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate949(.a(s_57), .b(gate146inter3), .O(gate146inter10));
  nor2  gate950(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate951(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate952(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1863(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1864(.a(gate148inter0), .b(s_188), .O(gate148inter1));
  and2  gate1865(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1866(.a(s_188), .O(gate148inter3));
  inv1  gate1867(.a(s_189), .O(gate148inter4));
  nand2 gate1868(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1869(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1870(.a(G492), .O(gate148inter7));
  inv1  gate1871(.a(G495), .O(gate148inter8));
  nand2 gate1872(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1873(.a(s_189), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1874(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1875(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1876(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate869(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate870(.a(gate150inter0), .b(s_46), .O(gate150inter1));
  and2  gate871(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate872(.a(s_46), .O(gate150inter3));
  inv1  gate873(.a(s_47), .O(gate150inter4));
  nand2 gate874(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate875(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate876(.a(G504), .O(gate150inter7));
  inv1  gate877(.a(G507), .O(gate150inter8));
  nand2 gate878(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate879(.a(s_47), .b(gate150inter3), .O(gate150inter10));
  nor2  gate880(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate881(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate882(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1345(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1346(.a(gate151inter0), .b(s_114), .O(gate151inter1));
  and2  gate1347(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1348(.a(s_114), .O(gate151inter3));
  inv1  gate1349(.a(s_115), .O(gate151inter4));
  nand2 gate1350(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1351(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1352(.a(G510), .O(gate151inter7));
  inv1  gate1353(.a(G513), .O(gate151inter8));
  nand2 gate1354(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1355(.a(s_115), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1356(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1357(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1358(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1765(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1766(.a(gate166inter0), .b(s_174), .O(gate166inter1));
  and2  gate1767(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1768(.a(s_174), .O(gate166inter3));
  inv1  gate1769(.a(s_175), .O(gate166inter4));
  nand2 gate1770(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1771(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1772(.a(G465), .O(gate166inter7));
  inv1  gate1773(.a(G540), .O(gate166inter8));
  nand2 gate1774(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1775(.a(s_175), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1776(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1777(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1778(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1331(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1332(.a(gate178inter0), .b(s_112), .O(gate178inter1));
  and2  gate1333(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1334(.a(s_112), .O(gate178inter3));
  inv1  gate1335(.a(s_113), .O(gate178inter4));
  nand2 gate1336(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1337(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1338(.a(G501), .O(gate178inter7));
  inv1  gate1339(.a(G558), .O(gate178inter8));
  nand2 gate1340(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1341(.a(s_113), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1342(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1343(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1344(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate785(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate786(.a(gate181inter0), .b(s_34), .O(gate181inter1));
  and2  gate787(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate788(.a(s_34), .O(gate181inter3));
  inv1  gate789(.a(s_35), .O(gate181inter4));
  nand2 gate790(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate791(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate792(.a(G510), .O(gate181inter7));
  inv1  gate793(.a(G564), .O(gate181inter8));
  nand2 gate794(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate795(.a(s_35), .b(gate181inter3), .O(gate181inter10));
  nor2  gate796(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate797(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate798(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate687(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate688(.a(gate185inter0), .b(s_20), .O(gate185inter1));
  and2  gate689(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate690(.a(s_20), .O(gate185inter3));
  inv1  gate691(.a(s_21), .O(gate185inter4));
  nand2 gate692(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate693(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate694(.a(G570), .O(gate185inter7));
  inv1  gate695(.a(G571), .O(gate185inter8));
  nand2 gate696(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate697(.a(s_21), .b(gate185inter3), .O(gate185inter10));
  nor2  gate698(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate699(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate700(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1513(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1514(.a(gate186inter0), .b(s_138), .O(gate186inter1));
  and2  gate1515(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1516(.a(s_138), .O(gate186inter3));
  inv1  gate1517(.a(s_139), .O(gate186inter4));
  nand2 gate1518(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1519(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1520(.a(G572), .O(gate186inter7));
  inv1  gate1521(.a(G573), .O(gate186inter8));
  nand2 gate1522(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1523(.a(s_139), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1524(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1525(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1526(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1877(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1878(.a(gate191inter0), .b(s_190), .O(gate191inter1));
  and2  gate1879(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1880(.a(s_190), .O(gate191inter3));
  inv1  gate1881(.a(s_191), .O(gate191inter4));
  nand2 gate1882(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1883(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1884(.a(G582), .O(gate191inter7));
  inv1  gate1885(.a(G583), .O(gate191inter8));
  nand2 gate1886(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1887(.a(s_191), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1888(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1889(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1890(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1191(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1192(.a(gate193inter0), .b(s_92), .O(gate193inter1));
  and2  gate1193(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1194(.a(s_92), .O(gate193inter3));
  inv1  gate1195(.a(s_93), .O(gate193inter4));
  nand2 gate1196(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1197(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1198(.a(G586), .O(gate193inter7));
  inv1  gate1199(.a(G587), .O(gate193inter8));
  nand2 gate1200(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1201(.a(s_93), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1202(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1203(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1204(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1849(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1850(.a(gate197inter0), .b(s_186), .O(gate197inter1));
  and2  gate1851(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1852(.a(s_186), .O(gate197inter3));
  inv1  gate1853(.a(s_187), .O(gate197inter4));
  nand2 gate1854(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1855(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1856(.a(G594), .O(gate197inter7));
  inv1  gate1857(.a(G595), .O(gate197inter8));
  nand2 gate1858(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1859(.a(s_187), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1860(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1861(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1862(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1205(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1206(.a(gate203inter0), .b(s_94), .O(gate203inter1));
  and2  gate1207(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1208(.a(s_94), .O(gate203inter3));
  inv1  gate1209(.a(s_95), .O(gate203inter4));
  nand2 gate1210(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1211(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1212(.a(G602), .O(gate203inter7));
  inv1  gate1213(.a(G612), .O(gate203inter8));
  nand2 gate1214(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1215(.a(s_95), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1216(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1217(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1218(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate603(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate604(.a(gate219inter0), .b(s_8), .O(gate219inter1));
  and2  gate605(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate606(.a(s_8), .O(gate219inter3));
  inv1  gate607(.a(s_9), .O(gate219inter4));
  nand2 gate608(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate609(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate610(.a(G632), .O(gate219inter7));
  inv1  gate611(.a(G681), .O(gate219inter8));
  nand2 gate612(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate613(.a(s_9), .b(gate219inter3), .O(gate219inter10));
  nor2  gate614(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate615(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate616(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1471(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1472(.a(gate224inter0), .b(s_132), .O(gate224inter1));
  and2  gate1473(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1474(.a(s_132), .O(gate224inter3));
  inv1  gate1475(.a(s_133), .O(gate224inter4));
  nand2 gate1476(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1477(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1478(.a(G637), .O(gate224inter7));
  inv1  gate1479(.a(G687), .O(gate224inter8));
  nand2 gate1480(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1481(.a(s_133), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1482(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1483(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1484(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1387(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1388(.a(gate234inter0), .b(s_120), .O(gate234inter1));
  and2  gate1389(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1390(.a(s_120), .O(gate234inter3));
  inv1  gate1391(.a(s_121), .O(gate234inter4));
  nand2 gate1392(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1393(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1394(.a(G245), .O(gate234inter7));
  inv1  gate1395(.a(G721), .O(gate234inter8));
  nand2 gate1396(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1397(.a(s_121), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1398(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1399(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1400(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate561(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate562(.a(gate253inter0), .b(s_2), .O(gate253inter1));
  and2  gate563(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate564(.a(s_2), .O(gate253inter3));
  inv1  gate565(.a(s_3), .O(gate253inter4));
  nand2 gate566(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate567(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate568(.a(G260), .O(gate253inter7));
  inv1  gate569(.a(G748), .O(gate253inter8));
  nand2 gate570(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate571(.a(s_3), .b(gate253inter3), .O(gate253inter10));
  nor2  gate572(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate573(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate574(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1219(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1220(.a(gate265inter0), .b(s_96), .O(gate265inter1));
  and2  gate1221(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1222(.a(s_96), .O(gate265inter3));
  inv1  gate1223(.a(s_97), .O(gate265inter4));
  nand2 gate1224(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1225(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1226(.a(G642), .O(gate265inter7));
  inv1  gate1227(.a(G770), .O(gate265inter8));
  nand2 gate1228(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1229(.a(s_97), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1230(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1231(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1232(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1667(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1668(.a(gate268inter0), .b(s_160), .O(gate268inter1));
  and2  gate1669(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1670(.a(s_160), .O(gate268inter3));
  inv1  gate1671(.a(s_161), .O(gate268inter4));
  nand2 gate1672(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1673(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1674(.a(G651), .O(gate268inter7));
  inv1  gate1675(.a(G779), .O(gate268inter8));
  nand2 gate1676(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1677(.a(s_161), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1678(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1679(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1680(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate645(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate646(.a(gate271inter0), .b(s_14), .O(gate271inter1));
  and2  gate647(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate648(.a(s_14), .O(gate271inter3));
  inv1  gate649(.a(s_15), .O(gate271inter4));
  nand2 gate650(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate651(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate652(.a(G660), .O(gate271inter7));
  inv1  gate653(.a(G788), .O(gate271inter8));
  nand2 gate654(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate655(.a(s_15), .b(gate271inter3), .O(gate271inter10));
  nor2  gate656(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate657(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate658(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1135(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1136(.a(gate272inter0), .b(s_84), .O(gate272inter1));
  and2  gate1137(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1138(.a(s_84), .O(gate272inter3));
  inv1  gate1139(.a(s_85), .O(gate272inter4));
  nand2 gate1140(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1141(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1142(.a(G663), .O(gate272inter7));
  inv1  gate1143(.a(G791), .O(gate272inter8));
  nand2 gate1144(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1145(.a(s_85), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1146(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1147(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1148(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1303(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1304(.a(gate273inter0), .b(s_108), .O(gate273inter1));
  and2  gate1305(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1306(.a(s_108), .O(gate273inter3));
  inv1  gate1307(.a(s_109), .O(gate273inter4));
  nand2 gate1308(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1309(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1310(.a(G642), .O(gate273inter7));
  inv1  gate1311(.a(G794), .O(gate273inter8));
  nand2 gate1312(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1313(.a(s_109), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1314(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1315(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1316(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate995(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate996(.a(gate274inter0), .b(s_64), .O(gate274inter1));
  and2  gate997(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate998(.a(s_64), .O(gate274inter3));
  inv1  gate999(.a(s_65), .O(gate274inter4));
  nand2 gate1000(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1001(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1002(.a(G770), .O(gate274inter7));
  inv1  gate1003(.a(G794), .O(gate274inter8));
  nand2 gate1004(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1005(.a(s_65), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1006(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1007(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1008(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate813(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate814(.a(gate279inter0), .b(s_38), .O(gate279inter1));
  and2  gate815(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate816(.a(s_38), .O(gate279inter3));
  inv1  gate817(.a(s_39), .O(gate279inter4));
  nand2 gate818(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate819(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate820(.a(G651), .O(gate279inter7));
  inv1  gate821(.a(G803), .O(gate279inter8));
  nand2 gate822(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate823(.a(s_39), .b(gate279inter3), .O(gate279inter10));
  nor2  gate824(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate825(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate826(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1093(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1094(.a(gate288inter0), .b(s_78), .O(gate288inter1));
  and2  gate1095(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1096(.a(s_78), .O(gate288inter3));
  inv1  gate1097(.a(s_79), .O(gate288inter4));
  nand2 gate1098(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1099(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1100(.a(G791), .O(gate288inter7));
  inv1  gate1101(.a(G815), .O(gate288inter8));
  nand2 gate1102(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1103(.a(s_79), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1104(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1105(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1106(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1023(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1024(.a(gate290inter0), .b(s_68), .O(gate290inter1));
  and2  gate1025(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1026(.a(s_68), .O(gate290inter3));
  inv1  gate1027(.a(s_69), .O(gate290inter4));
  nand2 gate1028(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1029(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1030(.a(G820), .O(gate290inter7));
  inv1  gate1031(.a(G821), .O(gate290inter8));
  nand2 gate1032(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1033(.a(s_69), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1034(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1035(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1036(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate799(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate800(.a(gate294inter0), .b(s_36), .O(gate294inter1));
  and2  gate801(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate802(.a(s_36), .O(gate294inter3));
  inv1  gate803(.a(s_37), .O(gate294inter4));
  nand2 gate804(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate805(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate806(.a(G832), .O(gate294inter7));
  inv1  gate807(.a(G833), .O(gate294inter8));
  nand2 gate808(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate809(.a(s_37), .b(gate294inter3), .O(gate294inter10));
  nor2  gate810(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate811(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate812(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1443(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1444(.a(gate395inter0), .b(s_128), .O(gate395inter1));
  and2  gate1445(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1446(.a(s_128), .O(gate395inter3));
  inv1  gate1447(.a(s_129), .O(gate395inter4));
  nand2 gate1448(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1449(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1450(.a(G9), .O(gate395inter7));
  inv1  gate1451(.a(G1060), .O(gate395inter8));
  nand2 gate1452(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1453(.a(s_129), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1454(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1455(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1456(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate771(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate772(.a(gate401inter0), .b(s_32), .O(gate401inter1));
  and2  gate773(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate774(.a(s_32), .O(gate401inter3));
  inv1  gate775(.a(s_33), .O(gate401inter4));
  nand2 gate776(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate777(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate778(.a(G15), .O(gate401inter7));
  inv1  gate779(.a(G1078), .O(gate401inter8));
  nand2 gate780(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate781(.a(s_33), .b(gate401inter3), .O(gate401inter10));
  nor2  gate782(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate783(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate784(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate673(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate674(.a(gate407inter0), .b(s_18), .O(gate407inter1));
  and2  gate675(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate676(.a(s_18), .O(gate407inter3));
  inv1  gate677(.a(s_19), .O(gate407inter4));
  nand2 gate678(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate679(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate680(.a(G21), .O(gate407inter7));
  inv1  gate681(.a(G1096), .O(gate407inter8));
  nand2 gate682(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate683(.a(s_19), .b(gate407inter3), .O(gate407inter10));
  nor2  gate684(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate685(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate686(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate897(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate898(.a(gate418inter0), .b(s_50), .O(gate418inter1));
  and2  gate899(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate900(.a(s_50), .O(gate418inter3));
  inv1  gate901(.a(s_51), .O(gate418inter4));
  nand2 gate902(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate903(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate904(.a(G32), .O(gate418inter7));
  inv1  gate905(.a(G1129), .O(gate418inter8));
  nand2 gate906(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate907(.a(s_51), .b(gate418inter3), .O(gate418inter10));
  nor2  gate908(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate909(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate910(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1527(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1528(.a(gate425inter0), .b(s_140), .O(gate425inter1));
  and2  gate1529(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1530(.a(s_140), .O(gate425inter3));
  inv1  gate1531(.a(s_141), .O(gate425inter4));
  nand2 gate1532(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1533(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1534(.a(G4), .O(gate425inter7));
  inv1  gate1535(.a(G1141), .O(gate425inter8));
  nand2 gate1536(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1537(.a(s_141), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1538(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1539(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1540(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1079(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1080(.a(gate433inter0), .b(s_76), .O(gate433inter1));
  and2  gate1081(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1082(.a(s_76), .O(gate433inter3));
  inv1  gate1083(.a(s_77), .O(gate433inter4));
  nand2 gate1084(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1085(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1086(.a(G8), .O(gate433inter7));
  inv1  gate1087(.a(G1153), .O(gate433inter8));
  nand2 gate1088(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1089(.a(s_77), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1090(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1091(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1092(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate743(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate744(.a(gate435inter0), .b(s_28), .O(gate435inter1));
  and2  gate745(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate746(.a(s_28), .O(gate435inter3));
  inv1  gate747(.a(s_29), .O(gate435inter4));
  nand2 gate748(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate749(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate750(.a(G9), .O(gate435inter7));
  inv1  gate751(.a(G1156), .O(gate435inter8));
  nand2 gate752(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate753(.a(s_29), .b(gate435inter3), .O(gate435inter10));
  nor2  gate754(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate755(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate756(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate967(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate968(.a(gate440inter0), .b(s_60), .O(gate440inter1));
  and2  gate969(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate970(.a(s_60), .O(gate440inter3));
  inv1  gate971(.a(s_61), .O(gate440inter4));
  nand2 gate972(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate973(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate974(.a(G1066), .O(gate440inter7));
  inv1  gate975(.a(G1162), .O(gate440inter8));
  nand2 gate976(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate977(.a(s_61), .b(gate440inter3), .O(gate440inter10));
  nor2  gate978(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate979(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate980(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate729(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate730(.a(gate443inter0), .b(s_26), .O(gate443inter1));
  and2  gate731(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate732(.a(s_26), .O(gate443inter3));
  inv1  gate733(.a(s_27), .O(gate443inter4));
  nand2 gate734(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate735(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate736(.a(G13), .O(gate443inter7));
  inv1  gate737(.a(G1168), .O(gate443inter8));
  nand2 gate738(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate739(.a(s_27), .b(gate443inter3), .O(gate443inter10));
  nor2  gate740(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate741(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate742(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1709(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1710(.a(gate445inter0), .b(s_166), .O(gate445inter1));
  and2  gate1711(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1712(.a(s_166), .O(gate445inter3));
  inv1  gate1713(.a(s_167), .O(gate445inter4));
  nand2 gate1714(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1715(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1716(.a(G14), .O(gate445inter7));
  inv1  gate1717(.a(G1171), .O(gate445inter8));
  nand2 gate1718(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1719(.a(s_167), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1720(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1721(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1722(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate631(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate632(.a(gate455inter0), .b(s_12), .O(gate455inter1));
  and2  gate633(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate634(.a(s_12), .O(gate455inter3));
  inv1  gate635(.a(s_13), .O(gate455inter4));
  nand2 gate636(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate637(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate638(.a(G19), .O(gate455inter7));
  inv1  gate639(.a(G1186), .O(gate455inter8));
  nand2 gate640(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate641(.a(s_13), .b(gate455inter3), .O(gate455inter10));
  nor2  gate642(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate643(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate644(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1541(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1542(.a(gate462inter0), .b(s_142), .O(gate462inter1));
  and2  gate1543(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1544(.a(s_142), .O(gate462inter3));
  inv1  gate1545(.a(s_143), .O(gate462inter4));
  nand2 gate1546(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1547(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1548(.a(G1099), .O(gate462inter7));
  inv1  gate1549(.a(G1195), .O(gate462inter8));
  nand2 gate1550(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1551(.a(s_143), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1552(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1553(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1554(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1163(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1164(.a(gate464inter0), .b(s_88), .O(gate464inter1));
  and2  gate1165(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1166(.a(s_88), .O(gate464inter3));
  inv1  gate1167(.a(s_89), .O(gate464inter4));
  nand2 gate1168(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1169(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1170(.a(G1102), .O(gate464inter7));
  inv1  gate1171(.a(G1198), .O(gate464inter8));
  nand2 gate1172(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1173(.a(s_89), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1174(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1175(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1176(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1247(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1248(.a(gate466inter0), .b(s_100), .O(gate466inter1));
  and2  gate1249(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1250(.a(s_100), .O(gate466inter3));
  inv1  gate1251(.a(s_101), .O(gate466inter4));
  nand2 gate1252(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1253(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1254(.a(G1105), .O(gate466inter7));
  inv1  gate1255(.a(G1201), .O(gate466inter8));
  nand2 gate1256(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1257(.a(s_101), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1258(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1259(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1260(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate883(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate884(.a(gate467inter0), .b(s_48), .O(gate467inter1));
  and2  gate885(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate886(.a(s_48), .O(gate467inter3));
  inv1  gate887(.a(s_49), .O(gate467inter4));
  nand2 gate888(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate889(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate890(.a(G25), .O(gate467inter7));
  inv1  gate891(.a(G1204), .O(gate467inter8));
  nand2 gate892(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate893(.a(s_49), .b(gate467inter3), .O(gate467inter10));
  nor2  gate894(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate895(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate896(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1359(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1360(.a(gate470inter0), .b(s_116), .O(gate470inter1));
  and2  gate1361(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1362(.a(s_116), .O(gate470inter3));
  inv1  gate1363(.a(s_117), .O(gate470inter4));
  nand2 gate1364(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1365(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1366(.a(G1111), .O(gate470inter7));
  inv1  gate1367(.a(G1207), .O(gate470inter8));
  nand2 gate1368(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1369(.a(s_117), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1370(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1371(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1372(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1261(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1262(.a(gate476inter0), .b(s_102), .O(gate476inter1));
  and2  gate1263(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1264(.a(s_102), .O(gate476inter3));
  inv1  gate1265(.a(s_103), .O(gate476inter4));
  nand2 gate1266(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1267(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1268(.a(G1120), .O(gate476inter7));
  inv1  gate1269(.a(G1216), .O(gate476inter8));
  nand2 gate1270(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1271(.a(s_103), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1272(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1273(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1274(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1597(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1598(.a(gate478inter0), .b(s_150), .O(gate478inter1));
  and2  gate1599(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1600(.a(s_150), .O(gate478inter3));
  inv1  gate1601(.a(s_151), .O(gate478inter4));
  nand2 gate1602(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1603(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1604(.a(G1123), .O(gate478inter7));
  inv1  gate1605(.a(G1219), .O(gate478inter8));
  nand2 gate1606(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1607(.a(s_151), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1608(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1609(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1610(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1793(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1794(.a(gate482inter0), .b(s_178), .O(gate482inter1));
  and2  gate1795(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1796(.a(s_178), .O(gate482inter3));
  inv1  gate1797(.a(s_179), .O(gate482inter4));
  nand2 gate1798(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1799(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1800(.a(G1129), .O(gate482inter7));
  inv1  gate1801(.a(G1225), .O(gate482inter8));
  nand2 gate1802(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1803(.a(s_179), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1804(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1805(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1806(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate547(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate548(.a(gate483inter0), .b(s_0), .O(gate483inter1));
  and2  gate549(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate550(.a(s_0), .O(gate483inter3));
  inv1  gate551(.a(s_1), .O(gate483inter4));
  nand2 gate552(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate553(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate554(.a(G1228), .O(gate483inter7));
  inv1  gate555(.a(G1229), .O(gate483inter8));
  nand2 gate556(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate557(.a(s_1), .b(gate483inter3), .O(gate483inter10));
  nor2  gate558(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate559(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate560(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate575(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate576(.a(gate489inter0), .b(s_4), .O(gate489inter1));
  and2  gate577(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate578(.a(s_4), .O(gate489inter3));
  inv1  gate579(.a(s_5), .O(gate489inter4));
  nand2 gate580(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate581(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate582(.a(G1240), .O(gate489inter7));
  inv1  gate583(.a(G1241), .O(gate489inter8));
  nand2 gate584(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate585(.a(s_5), .b(gate489inter3), .O(gate489inter10));
  nor2  gate586(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate587(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate588(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1009(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1010(.a(gate490inter0), .b(s_66), .O(gate490inter1));
  and2  gate1011(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1012(.a(s_66), .O(gate490inter3));
  inv1  gate1013(.a(s_67), .O(gate490inter4));
  nand2 gate1014(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1015(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1016(.a(G1242), .O(gate490inter7));
  inv1  gate1017(.a(G1243), .O(gate490inter8));
  nand2 gate1018(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1019(.a(s_67), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1020(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1021(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1022(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1149(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1150(.a(gate494inter0), .b(s_86), .O(gate494inter1));
  and2  gate1151(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1152(.a(s_86), .O(gate494inter3));
  inv1  gate1153(.a(s_87), .O(gate494inter4));
  nand2 gate1154(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1155(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1156(.a(G1250), .O(gate494inter7));
  inv1  gate1157(.a(G1251), .O(gate494inter8));
  nand2 gate1158(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1159(.a(s_87), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1160(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1161(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1162(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1275(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1276(.a(gate495inter0), .b(s_104), .O(gate495inter1));
  and2  gate1277(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1278(.a(s_104), .O(gate495inter3));
  inv1  gate1279(.a(s_105), .O(gate495inter4));
  nand2 gate1280(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1281(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1282(.a(G1252), .O(gate495inter7));
  inv1  gate1283(.a(G1253), .O(gate495inter8));
  nand2 gate1284(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1285(.a(s_105), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1286(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1287(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1288(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate1583(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1584(.a(gate496inter0), .b(s_148), .O(gate496inter1));
  and2  gate1585(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1586(.a(s_148), .O(gate496inter3));
  inv1  gate1587(.a(s_149), .O(gate496inter4));
  nand2 gate1588(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1589(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1590(.a(G1254), .O(gate496inter7));
  inv1  gate1591(.a(G1255), .O(gate496inter8));
  nand2 gate1592(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1593(.a(s_149), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1594(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1595(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1596(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate617(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate618(.a(gate497inter0), .b(s_10), .O(gate497inter1));
  and2  gate619(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate620(.a(s_10), .O(gate497inter3));
  inv1  gate621(.a(s_11), .O(gate497inter4));
  nand2 gate622(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate623(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate624(.a(G1256), .O(gate497inter7));
  inv1  gate625(.a(G1257), .O(gate497inter8));
  nand2 gate626(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate627(.a(s_11), .b(gate497inter3), .O(gate497inter10));
  nor2  gate628(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate629(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate630(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1415(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1416(.a(gate511inter0), .b(s_124), .O(gate511inter1));
  and2  gate1417(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1418(.a(s_124), .O(gate511inter3));
  inv1  gate1419(.a(s_125), .O(gate511inter4));
  nand2 gate1420(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1421(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1422(.a(G1284), .O(gate511inter7));
  inv1  gate1423(.a(G1285), .O(gate511inter8));
  nand2 gate1424(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1425(.a(s_125), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1426(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1427(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1428(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate827(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate828(.a(gate512inter0), .b(s_40), .O(gate512inter1));
  and2  gate829(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate830(.a(s_40), .O(gate512inter3));
  inv1  gate831(.a(s_41), .O(gate512inter4));
  nand2 gate832(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate833(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate834(.a(G1286), .O(gate512inter7));
  inv1  gate835(.a(G1287), .O(gate512inter8));
  nand2 gate836(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate837(.a(s_41), .b(gate512inter3), .O(gate512inter10));
  nor2  gate838(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate839(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate840(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate855(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate856(.a(gate514inter0), .b(s_44), .O(gate514inter1));
  and2  gate857(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate858(.a(s_44), .O(gate514inter3));
  inv1  gate859(.a(s_45), .O(gate514inter4));
  nand2 gate860(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate861(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate862(.a(G1290), .O(gate514inter7));
  inv1  gate863(.a(G1291), .O(gate514inter8));
  nand2 gate864(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate865(.a(s_45), .b(gate514inter3), .O(gate514inter10));
  nor2  gate866(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate867(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate868(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule