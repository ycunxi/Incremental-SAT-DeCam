module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate511(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate512(.a(gate24inter0), .b(s_50), .O(gate24inter1));
  and2  gate513(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate514(.a(s_50), .O(gate24inter3));
  inv1  gate515(.a(s_51), .O(gate24inter4));
  nand2 gate516(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate517(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate518(.a(N130), .O(gate24inter7));
  inv1  gate519(.a(N43), .O(gate24inter8));
  nand2 gate520(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate521(.a(s_51), .b(gate24inter3), .O(gate24inter10));
  nor2  gate522(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate523(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate524(.a(gate24inter12), .b(gate24inter1), .O(N165));

  xor2  gate567(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate568(.a(gate25inter0), .b(s_58), .O(gate25inter1));
  and2  gate569(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate570(.a(s_58), .O(gate25inter3));
  inv1  gate571(.a(s_59), .O(gate25inter4));
  nand2 gate572(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate573(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate574(.a(N134), .O(gate25inter7));
  inv1  gate575(.a(N56), .O(gate25inter8));
  nand2 gate576(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate577(.a(s_59), .b(gate25inter3), .O(gate25inter10));
  nor2  gate578(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate579(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate580(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate441(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate442(.a(gate29inter0), .b(s_40), .O(gate29inter1));
  and2  gate443(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate444(.a(s_40), .O(gate29inter3));
  inv1  gate445(.a(s_41), .O(gate29inter4));
  nand2 gate446(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate447(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate448(.a(N150), .O(gate29inter7));
  inv1  gate449(.a(N108), .O(gate29inter8));
  nand2 gate450(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate451(.a(s_41), .b(gate29inter3), .O(gate29inter10));
  nor2  gate452(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate453(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate454(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );

  xor2  gate371(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate372(.a(gate31inter0), .b(s_30), .O(gate31inter1));
  and2  gate373(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate374(.a(s_30), .O(gate31inter3));
  inv1  gate375(.a(s_31), .O(gate31inter4));
  nand2 gate376(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate377(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate378(.a(N27), .O(gate31inter7));
  inv1  gate379(.a(N123), .O(gate31inter8));
  nand2 gate380(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate381(.a(s_31), .b(gate31inter3), .O(gate31inter10));
  nor2  gate382(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate383(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate384(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );

  xor2  gate189(.a(N127), .b(N40), .O(gate33inter0));
  nand2 gate190(.a(gate33inter0), .b(s_4), .O(gate33inter1));
  and2  gate191(.a(N127), .b(N40), .O(gate33inter2));
  inv1  gate192(.a(s_4), .O(gate33inter3));
  inv1  gate193(.a(s_5), .O(gate33inter4));
  nand2 gate194(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate195(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate196(.a(N40), .O(gate33inter7));
  inv1  gate197(.a(N127), .O(gate33inter8));
  nand2 gate198(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate199(.a(s_5), .b(gate33inter3), .O(gate33inter10));
  nor2  gate200(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate201(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate202(.a(gate33inter12), .b(gate33inter1), .O(N186));

  xor2  gate455(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate456(.a(gate34inter0), .b(s_42), .O(gate34inter1));
  and2  gate457(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate458(.a(s_42), .O(gate34inter3));
  inv1  gate459(.a(s_43), .O(gate34inter4));
  nand2 gate460(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate461(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate462(.a(N47), .O(gate34inter7));
  inv1  gate463(.a(N131), .O(gate34inter8));
  nand2 gate464(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate465(.a(s_43), .b(gate34inter3), .O(gate34inter10));
  nor2  gate466(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate467(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate468(.a(gate34inter12), .b(gate34inter1), .O(N187));
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate217(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate218(.a(gate37inter0), .b(s_8), .O(gate37inter1));
  and2  gate219(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate220(.a(s_8), .O(gate37inter3));
  inv1  gate221(.a(s_9), .O(gate37inter4));
  nand2 gate222(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate223(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate224(.a(N66), .O(gate37inter7));
  inv1  gate225(.a(N135), .O(gate37inter8));
  nand2 gate226(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate227(.a(s_9), .b(gate37inter3), .O(gate37inter10));
  nor2  gate228(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate229(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate230(.a(gate37inter12), .b(gate37inter1), .O(N190));

  xor2  gate273(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate274(.a(gate38inter0), .b(s_16), .O(gate38inter1));
  and2  gate275(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate276(.a(s_16), .O(gate38inter3));
  inv1  gate277(.a(s_17), .O(gate38inter4));
  nand2 gate278(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate279(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate280(.a(N73), .O(gate38inter7));
  inv1  gate281(.a(N139), .O(gate38inter8));
  nand2 gate282(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate283(.a(s_17), .b(gate38inter3), .O(gate38inter10));
  nor2  gate284(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate285(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate286(.a(gate38inter12), .b(gate38inter1), .O(N191));
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );

  xor2  gate231(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate232(.a(gate42inter0), .b(s_10), .O(gate42inter1));
  and2  gate233(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate234(.a(s_10), .O(gate42inter3));
  inv1  gate235(.a(s_11), .O(gate42inter4));
  nand2 gate236(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate237(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate238(.a(N99), .O(gate42inter7));
  inv1  gate239(.a(N147), .O(gate42inter8));
  nand2 gate240(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate241(.a(s_11), .b(gate42inter3), .O(gate42inter10));
  nor2  gate242(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate243(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate244(.a(gate42inter12), .b(gate42inter1), .O(N195));

  xor2  gate427(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate428(.a(gate43inter0), .b(s_38), .O(gate43inter1));
  and2  gate429(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate430(.a(s_38), .O(gate43inter3));
  inv1  gate431(.a(s_39), .O(gate43inter4));
  nand2 gate432(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate433(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate434(.a(N105), .O(gate43inter7));
  inv1  gate435(.a(N147), .O(gate43inter8));
  nand2 gate436(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate437(.a(s_39), .b(gate43inter3), .O(gate43inter10));
  nor2  gate438(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate439(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate440(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate301(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate302(.a(gate50inter0), .b(s_20), .O(gate50inter1));
  and2  gate303(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate304(.a(s_20), .O(gate50inter3));
  inv1  gate305(.a(s_21), .O(gate50inter4));
  nand2 gate306(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate307(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate308(.a(N203), .O(gate50inter7));
  inv1  gate309(.a(N154), .O(gate50inter8));
  nand2 gate310(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate311(.a(s_21), .b(gate50inter3), .O(gate50inter10));
  nor2  gate312(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate313(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate314(.a(gate50inter12), .b(gate50inter1), .O(N224));

  xor2  gate343(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate344(.a(gate51inter0), .b(s_26), .O(gate51inter1));
  and2  gate345(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate346(.a(s_26), .O(gate51inter3));
  inv1  gate347(.a(s_27), .O(gate51inter4));
  nand2 gate348(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate349(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate350(.a(N203), .O(gate51inter7));
  inv1  gate351(.a(N159), .O(gate51inter8));
  nand2 gate352(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate353(.a(s_27), .b(gate51inter3), .O(gate51inter10));
  nor2  gate354(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate355(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate356(.a(gate51inter12), .b(gate51inter1), .O(N227));

  xor2  gate315(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate316(.a(gate52inter0), .b(s_22), .O(gate52inter1));
  and2  gate317(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate318(.a(s_22), .O(gate52inter3));
  inv1  gate319(.a(s_23), .O(gate52inter4));
  nand2 gate320(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate321(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate322(.a(N203), .O(gate52inter7));
  inv1  gate323(.a(N162), .O(gate52inter8));
  nand2 gate324(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate325(.a(s_23), .b(gate52inter3), .O(gate52inter10));
  nor2  gate326(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate327(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate328(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );

  xor2  gate413(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate414(.a(gate55inter0), .b(s_36), .O(gate55inter1));
  and2  gate415(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate416(.a(s_36), .O(gate55inter3));
  inv1  gate417(.a(s_37), .O(gate55inter4));
  nand2 gate418(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate419(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate420(.a(N203), .O(gate55inter7));
  inv1  gate421(.a(N171), .O(gate55inter8));
  nand2 gate422(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate423(.a(s_37), .b(gate55inter3), .O(gate55inter10));
  nor2  gate424(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate425(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate426(.a(gate55inter12), .b(gate55inter1), .O(N239));

  xor2  gate483(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate484(.a(gate56inter0), .b(s_46), .O(gate56inter1));
  and2  gate485(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate486(.a(s_46), .O(gate56inter3));
  inv1  gate487(.a(s_47), .O(gate56inter4));
  nand2 gate488(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate489(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate490(.a(N1), .O(gate56inter7));
  inv1  gate491(.a(N213), .O(gate56inter8));
  nand2 gate492(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate493(.a(s_47), .b(gate56inter3), .O(gate56inter10));
  nor2  gate494(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate495(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate496(.a(gate56inter12), .b(gate56inter1), .O(N242));
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );

  xor2  gate287(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate288(.a(gate67inter0), .b(s_18), .O(gate67inter1));
  and2  gate289(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate290(.a(s_18), .O(gate67inter3));
  inv1  gate291(.a(s_19), .O(gate67inter4));
  nand2 gate292(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate293(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate294(.a(N213), .O(gate67inter7));
  inv1  gate295(.a(N102), .O(gate67inter8));
  nand2 gate296(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate297(.a(s_19), .b(gate67inter3), .O(gate67inter10));
  nor2  gate298(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate299(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate300(.a(gate67inter12), .b(gate67inter1), .O(N259));
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate553(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate554(.a(gate72inter0), .b(s_56), .O(gate72inter1));
  and2  gate555(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate556(.a(s_56), .O(gate72inter3));
  inv1  gate557(.a(s_57), .O(gate72inter4));
  nand2 gate558(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate559(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate560(.a(N233), .O(gate72inter7));
  inv1  gate561(.a(N187), .O(gate72inter8));
  nand2 gate562(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate563(.a(s_57), .b(gate72inter3), .O(gate72inter10));
  nor2  gate564(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate565(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate566(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate357(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate358(.a(gate75inter0), .b(s_28), .O(gate75inter1));
  and2  gate359(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate360(.a(s_28), .O(gate75inter3));
  inv1  gate361(.a(s_29), .O(gate75inter4));
  nand2 gate362(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate363(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate364(.a(N243), .O(gate75inter7));
  inv1  gate365(.a(N193), .O(gate75inter8));
  nand2 gate366(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate367(.a(s_29), .b(gate75inter3), .O(gate75inter10));
  nor2  gate368(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate369(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate370(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );

  xor2  gate399(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate400(.a(gate79inter0), .b(s_34), .O(gate79inter1));
  and2  gate401(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate402(.a(s_34), .O(gate79inter3));
  inv1  gate403(.a(s_35), .O(gate79inter4));
  nand2 gate404(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate405(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate406(.a(N230), .O(gate79inter7));
  inv1  gate407(.a(N186), .O(gate79inter8));
  nand2 gate408(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate409(.a(s_35), .b(gate79inter3), .O(gate79inter10));
  nor2  gate410(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate411(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate412(.a(gate79inter12), .b(gate79inter1), .O(N289));
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );

  xor2  gate259(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate260(.a(gate82inter0), .b(s_14), .O(gate82inter1));
  and2  gate261(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate262(.a(s_14), .O(gate82inter3));
  inv1  gate263(.a(s_15), .O(gate82inter4));
  nand2 gate264(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate265(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate266(.a(N239), .O(gate82inter7));
  inv1  gate267(.a(N192), .O(gate82inter8));
  nand2 gate268(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate269(.a(s_15), .b(gate82inter3), .O(gate82inter10));
  nor2  gate270(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate271(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate272(.a(gate82inter12), .b(gate82inter1), .O(N292));
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate469(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate470(.a(gate103inter0), .b(s_44), .O(gate103inter1));
  and2  gate471(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate472(.a(s_44), .O(gate103inter3));
  inv1  gate473(.a(s_45), .O(gate103inter4));
  nand2 gate474(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate475(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate476(.a(N8), .O(gate103inter7));
  inv1  gate477(.a(N319), .O(gate103inter8));
  nand2 gate478(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate479(.a(s_45), .b(gate103inter3), .O(gate103inter10));
  nor2  gate480(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate481(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate482(.a(gate103inter12), .b(gate103inter1), .O(N334));

  xor2  gate245(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate246(.a(gate104inter0), .b(s_12), .O(gate104inter1));
  and2  gate247(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate248(.a(s_12), .O(gate104inter3));
  inv1  gate249(.a(s_13), .O(gate104inter4));
  nand2 gate250(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate251(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate252(.a(N309), .O(gate104inter7));
  inv1  gate253(.a(N273), .O(gate104inter8));
  nand2 gate254(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate255(.a(s_13), .b(gate104inter3), .O(gate104inter10));
  nor2  gate256(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate257(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate258(.a(gate104inter12), .b(gate104inter1), .O(N335));

  xor2  gate525(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate526(.a(gate105inter0), .b(s_52), .O(gate105inter1));
  and2  gate527(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate528(.a(s_52), .O(gate105inter3));
  inv1  gate529(.a(s_53), .O(gate105inter4));
  nand2 gate530(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate531(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate532(.a(N319), .O(gate105inter7));
  inv1  gate533(.a(N21), .O(gate105inter8));
  nand2 gate534(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate535(.a(s_53), .b(gate105inter3), .O(gate105inter10));
  nor2  gate536(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate537(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate538(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate385(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate386(.a(gate110inter0), .b(s_32), .O(gate110inter1));
  and2  gate387(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate388(.a(s_32), .O(gate110inter3));
  inv1  gate389(.a(s_33), .O(gate110inter4));
  nand2 gate390(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate391(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate392(.a(N309), .O(gate110inter7));
  inv1  gate393(.a(N282), .O(gate110inter8));
  nand2 gate394(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate395(.a(s_33), .b(gate110inter3), .O(gate110inter10));
  nor2  gate396(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate397(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate398(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );

  xor2  gate497(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate498(.a(gate112inter0), .b(s_48), .O(gate112inter1));
  and2  gate499(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate500(.a(s_48), .O(gate112inter3));
  inv1  gate501(.a(s_49), .O(gate112inter4));
  nand2 gate502(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate503(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate504(.a(N309), .O(gate112inter7));
  inv1  gate505(.a(N285), .O(gate112inter8));
  nand2 gate506(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate507(.a(s_49), .b(gate112inter3), .O(gate112inter10));
  nor2  gate508(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate509(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate510(.a(gate112inter12), .b(gate112inter1), .O(N343));

  xor2  gate539(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate540(.a(gate113inter0), .b(s_54), .O(gate113inter1));
  and2  gate541(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate542(.a(s_54), .O(gate113inter3));
  inv1  gate543(.a(s_55), .O(gate113inter4));
  nand2 gate544(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate545(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate546(.a(N319), .O(gate113inter7));
  inv1  gate547(.a(N73), .O(gate113inter8));
  nand2 gate548(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate549(.a(s_55), .b(gate113inter3), .O(gate113inter10));
  nor2  gate550(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate551(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate552(.a(gate113inter12), .b(gate113inter1), .O(N344));

  xor2  gate581(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate582(.a(gate114inter0), .b(s_60), .O(gate114inter1));
  and2  gate583(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate584(.a(s_60), .O(gate114inter3));
  inv1  gate585(.a(s_61), .O(gate114inter4));
  nand2 gate586(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate587(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate588(.a(N319), .O(gate114inter7));
  inv1  gate589(.a(N86), .O(gate114inter8));
  nand2 gate590(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate591(.a(s_61), .b(gate114inter3), .O(gate114inter10));
  nor2  gate592(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate593(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate594(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate175(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate176(.a(gate119inter0), .b(s_2), .O(gate119inter1));
  and2  gate177(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate178(.a(s_2), .O(gate119inter3));
  inv1  gate179(.a(s_3), .O(gate119inter4));
  nand2 gate180(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate181(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate182(.a(N332), .O(gate119inter7));
  inv1  gate183(.a(N302), .O(gate119inter8));
  nand2 gate184(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate185(.a(s_3), .b(gate119inter3), .O(gate119inter10));
  nor2  gate186(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate187(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate188(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );

  xor2  gate161(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate162(.a(gate122inter0), .b(s_0), .O(gate122inter1));
  and2  gate163(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate164(.a(s_0), .O(gate122inter3));
  inv1  gate165(.a(s_1), .O(gate122inter4));
  nand2 gate166(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate167(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate168(.a(N337), .O(gate122inter7));
  inv1  gate169(.a(N305), .O(gate122inter8));
  nand2 gate170(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate171(.a(s_1), .b(gate122inter3), .O(gate122inter10));
  nor2  gate172(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate173(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate174(.a(gate122inter12), .b(gate122inter1), .O(N353));
nand2 gate123( .a(N339), .b(N306), .O(N354) );

  xor2  gate203(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate204(.a(gate124inter0), .b(s_6), .O(gate124inter1));
  and2  gate205(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate206(.a(s_6), .O(gate124inter3));
  inv1  gate207(.a(s_7), .O(gate124inter4));
  nand2 gate208(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate209(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate210(.a(N341), .O(gate124inter7));
  inv1  gate211(.a(N307), .O(gate124inter8));
  nand2 gate212(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate213(.a(s_7), .b(gate124inter3), .O(gate124inter10));
  nor2  gate214(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate215(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate216(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate329(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate330(.a(gate131inter0), .b(s_24), .O(gate131inter1));
  and2  gate331(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate332(.a(s_24), .O(gate131inter3));
  inv1  gate333(.a(s_25), .O(gate131inter4));
  nand2 gate334(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate335(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate336(.a(N360), .O(gate131inter7));
  inv1  gate337(.a(N40), .O(gate131inter8));
  nand2 gate338(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate339(.a(s_25), .b(gate131inter3), .O(gate131inter10));
  nor2  gate340(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate341(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate342(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule