module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );

  xor2  gate301(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate302(.a(gate2inter0), .b(s_14), .O(gate2inter1));
  and2  gate303(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate304(.a(s_14), .O(gate2inter3));
  inv1  gate305(.a(s_15), .O(gate2inter4));
  nand2 gate306(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate307(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate308(.a(N9), .O(gate2inter7));
  inv1  gate309(.a(N13), .O(gate2inter8));
  nand2 gate310(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate311(.a(s_15), .b(gate2inter3), .O(gate2inter10));
  nor2  gate312(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate313(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate314(.a(gate2inter12), .b(gate2inter1), .O(N251));

  xor2  gate357(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate358(.a(gate3inter0), .b(s_22), .O(gate3inter1));
  and2  gate359(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate360(.a(s_22), .O(gate3inter3));
  inv1  gate361(.a(s_23), .O(gate3inter4));
  nand2 gate362(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate363(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate364(.a(N17), .O(gate3inter7));
  inv1  gate365(.a(N21), .O(gate3inter8));
  nand2 gate366(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate367(.a(s_23), .b(gate3inter3), .O(gate3inter10));
  nor2  gate368(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate369(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate370(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );

  xor2  gate203(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate204(.a(gate5inter0), .b(s_0), .O(gate5inter1));
  and2  gate205(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate206(.a(s_0), .O(gate5inter3));
  inv1  gate207(.a(s_1), .O(gate5inter4));
  nand2 gate208(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate209(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate210(.a(N33), .O(gate5inter7));
  inv1  gate211(.a(N37), .O(gate5inter8));
  nand2 gate212(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate213(.a(s_1), .b(gate5inter3), .O(gate5inter10));
  nor2  gate214(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate215(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate216(.a(gate5inter12), .b(gate5inter1), .O(N254));

  xor2  gate231(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate232(.a(gate6inter0), .b(s_4), .O(gate6inter1));
  and2  gate233(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate234(.a(s_4), .O(gate6inter3));
  inv1  gate235(.a(s_5), .O(gate6inter4));
  nand2 gate236(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate237(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate238(.a(N41), .O(gate6inter7));
  inv1  gate239(.a(N45), .O(gate6inter8));
  nand2 gate240(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate241(.a(s_5), .b(gate6inter3), .O(gate6inter10));
  nor2  gate242(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate243(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate244(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );

  xor2  gate441(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate442(.a(gate10inter0), .b(s_34), .O(gate10inter1));
  and2  gate443(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate444(.a(s_34), .O(gate10inter3));
  inv1  gate445(.a(s_35), .O(gate10inter4));
  nand2 gate446(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate447(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate448(.a(N73), .O(gate10inter7));
  inv1  gate449(.a(N77), .O(gate10inter8));
  nand2 gate450(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate451(.a(s_35), .b(gate10inter3), .O(gate10inter10));
  nor2  gate452(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate453(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate454(.a(gate10inter12), .b(gate10inter1), .O(N259));
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );

  xor2  gate287(.a(N109), .b(N105), .O(gate14inter0));
  nand2 gate288(.a(gate14inter0), .b(s_12), .O(gate14inter1));
  and2  gate289(.a(N109), .b(N105), .O(gate14inter2));
  inv1  gate290(.a(s_12), .O(gate14inter3));
  inv1  gate291(.a(s_13), .O(gate14inter4));
  nand2 gate292(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate293(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate294(.a(N105), .O(gate14inter7));
  inv1  gate295(.a(N109), .O(gate14inter8));
  nand2 gate296(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate297(.a(s_13), .b(gate14inter3), .O(gate14inter10));
  nor2  gate298(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate299(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate300(.a(gate14inter12), .b(gate14inter1), .O(N263));
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );

  xor2  gate497(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate498(.a(gate26inter0), .b(s_42), .O(gate26inter1));
  and2  gate499(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate500(.a(s_42), .O(gate26inter3));
  inv1  gate501(.a(s_43), .O(gate26inter4));
  nand2 gate502(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate503(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate504(.a(N33), .O(gate26inter7));
  inv1  gate505(.a(N49), .O(gate26inter8));
  nand2 gate506(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate507(.a(s_43), .b(gate26inter3), .O(gate26inter10));
  nor2  gate508(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate509(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate510(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );

  xor2  gate217(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate218(.a(gate33inter0), .b(s_2), .O(gate33inter1));
  and2  gate219(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate220(.a(s_2), .O(gate33inter3));
  inv1  gate221(.a(s_3), .O(gate33inter4));
  nand2 gate222(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate223(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate224(.a(N65), .O(gate33inter7));
  inv1  gate225(.a(N81), .O(gate33inter8));
  nand2 gate226(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate227(.a(s_3), .b(gate33inter3), .O(gate33inter10));
  nor2  gate228(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate229(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate230(.a(gate33inter12), .b(gate33inter1), .O(N282));
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );

  xor2  gate539(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate540(.a(gate37inter0), .b(s_48), .O(gate37inter1));
  and2  gate541(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate542(.a(s_48), .O(gate37inter3));
  inv1  gate543(.a(s_49), .O(gate37inter4));
  nand2 gate544(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate545(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate546(.a(N73), .O(gate37inter7));
  inv1  gate547(.a(N89), .O(gate37inter8));
  nand2 gate548(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate549(.a(s_49), .b(gate37inter3), .O(gate37inter10));
  nor2  gate550(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate551(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate552(.a(gate37inter12), .b(gate37inter1), .O(N286));

  xor2  gate469(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate470(.a(gate38inter0), .b(s_38), .O(gate38inter1));
  and2  gate471(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate472(.a(s_38), .O(gate38inter3));
  inv1  gate473(.a(s_39), .O(gate38inter4));
  nand2 gate474(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate475(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate476(.a(N105), .O(gate38inter7));
  inv1  gate477(.a(N121), .O(gate38inter8));
  nand2 gate478(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate479(.a(s_39), .b(gate38inter3), .O(gate38inter10));
  nor2  gate480(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate481(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate482(.a(gate38inter12), .b(gate38inter1), .O(N287));
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate483(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate484(.a(gate47inter0), .b(s_40), .O(gate47inter1));
  and2  gate485(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate486(.a(s_40), .O(gate47inter3));
  inv1  gate487(.a(s_41), .O(gate47inter4));
  nand2 gate488(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate489(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate490(.a(N262), .O(gate47inter7));
  inv1  gate491(.a(N263), .O(gate47inter8));
  nand2 gate492(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate493(.a(s_41), .b(gate47inter3), .O(gate47inter10));
  nor2  gate494(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate495(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate496(.a(gate47inter12), .b(gate47inter1), .O(N308));

  xor2  gate343(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate344(.a(gate48inter0), .b(s_20), .O(gate48inter1));
  and2  gate345(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate346(.a(s_20), .O(gate48inter3));
  inv1  gate347(.a(s_21), .O(gate48inter4));
  nand2 gate348(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate349(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate350(.a(N264), .O(gate48inter7));
  inv1  gate351(.a(N265), .O(gate48inter8));
  nand2 gate352(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate353(.a(s_21), .b(gate48inter3), .O(gate48inter10));
  nor2  gate354(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate355(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate356(.a(gate48inter12), .b(gate48inter1), .O(N311));
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );

  xor2  gate399(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate400(.a(gate51inter0), .b(s_28), .O(gate51inter1));
  and2  gate401(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate402(.a(s_28), .O(gate51inter3));
  inv1  gate403(.a(s_29), .O(gate51inter4));
  nand2 gate404(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate405(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate406(.a(N278), .O(gate51inter7));
  inv1  gate407(.a(N279), .O(gate51inter8));
  nand2 gate408(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate409(.a(s_29), .b(gate51inter3), .O(gate51inter10));
  nor2  gate410(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate411(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate412(.a(gate51inter12), .b(gate51inter1), .O(N316));
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate385(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate386(.a(gate55inter0), .b(s_26), .O(gate55inter1));
  and2  gate387(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate388(.a(s_26), .O(gate55inter3));
  inv1  gate389(.a(s_27), .O(gate55inter4));
  nand2 gate390(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate391(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate392(.a(N286), .O(gate55inter7));
  inv1  gate393(.a(N287), .O(gate55inter8));
  nand2 gate394(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate395(.a(s_27), .b(gate55inter3), .O(gate55inter10));
  nor2  gate396(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate397(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate398(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate511(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate512(.a(gate62inter0), .b(s_44), .O(gate62inter1));
  and2  gate513(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate514(.a(s_44), .O(gate62inter3));
  inv1  gate515(.a(s_45), .O(gate62inter4));
  nand2 gate516(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate517(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate518(.a(N308), .O(gate62inter7));
  inv1  gate519(.a(N311), .O(gate62inter8));
  nand2 gate520(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate521(.a(s_45), .b(gate62inter3), .O(gate62inter10));
  nor2  gate522(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate523(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate524(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );

  xor2  gate455(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate456(.a(gate67inter0), .b(s_36), .O(gate67inter1));
  and2  gate457(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate458(.a(s_36), .O(gate67inter3));
  inv1  gate459(.a(s_37), .O(gate67inter4));
  nand2 gate460(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate461(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate462(.a(N268), .O(gate67inter7));
  inv1  gate463(.a(N344), .O(gate67inter8));
  nand2 gate464(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate465(.a(s_37), .b(gate67inter3), .O(gate67inter10));
  nor2  gate466(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate467(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate468(.a(gate67inter12), .b(gate67inter1), .O(N348));
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate273(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate274(.a(gate70inter0), .b(s_10), .O(gate70inter1));
  and2  gate275(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate276(.a(s_10), .O(gate70inter3));
  inv1  gate277(.a(s_11), .O(gate70inter4));
  nand2 gate278(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate279(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate280(.a(N271), .O(gate70inter7));
  inv1  gate281(.a(N339), .O(gate70inter8));
  nand2 gate282(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate283(.a(s_11), .b(gate70inter3), .O(gate70inter10));
  nor2  gate284(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate285(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate286(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );

  xor2  gate371(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate372(.a(gate77inter0), .b(s_24), .O(gate77inter1));
  and2  gate373(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate374(.a(s_24), .O(gate77inter3));
  inv1  gate375(.a(s_25), .O(gate77inter4));
  nand2 gate376(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate377(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate378(.a(N318), .O(gate77inter7));
  inv1  gate379(.a(N350), .O(gate77inter8));
  nand2 gate380(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate381(.a(s_25), .b(gate77inter3), .O(gate77inter10));
  nor2  gate382(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate383(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate384(.a(gate77inter12), .b(gate77inter1), .O(N406));
xor2 gate78( .a(N319), .b(N351), .O(N419) );

  xor2  gate259(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate260(.a(gate79inter0), .b(s_8), .O(gate79inter1));
  and2  gate261(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate262(.a(s_8), .O(gate79inter3));
  inv1  gate263(.a(s_9), .O(gate79inter4));
  nand2 gate264(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate265(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate266(.a(N320), .O(gate79inter7));
  inv1  gate267(.a(N352), .O(gate79inter8));
  nand2 gate268(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate269(.a(s_9), .b(gate79inter3), .O(gate79inter10));
  nor2  gate270(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate271(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate272(.a(gate79inter12), .b(gate79inter1), .O(N432));
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate315(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate316(.a(gate177inter0), .b(s_16), .O(gate177inter1));
  and2  gate317(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate318(.a(s_16), .O(gate177inter3));
  inv1  gate319(.a(s_17), .O(gate177inter4));
  nand2 gate320(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate321(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate322(.a(N25), .O(gate177inter7));
  inv1  gate323(.a(N698), .O(gate177inter8));
  nand2 gate324(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate325(.a(s_17), .b(gate177inter3), .O(gate177inter10));
  nor2  gate326(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate327(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate328(.a(gate177inter12), .b(gate177inter1), .O(N730));
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );

  xor2  gate329(.a(N701), .b(N37), .O(gate180inter0));
  nand2 gate330(.a(gate180inter0), .b(s_18), .O(gate180inter1));
  and2  gate331(.a(N701), .b(N37), .O(gate180inter2));
  inv1  gate332(.a(s_18), .O(gate180inter3));
  inv1  gate333(.a(s_19), .O(gate180inter4));
  nand2 gate334(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate335(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate336(.a(N37), .O(gate180inter7));
  inv1  gate337(.a(N701), .O(gate180inter8));
  nand2 gate338(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate339(.a(s_19), .b(gate180inter3), .O(gate180inter10));
  nor2  gate340(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate341(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate342(.a(gate180inter12), .b(gate180inter1), .O(N733));
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );

  xor2  gate553(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate554(.a(gate187inter0), .b(s_50), .O(gate187inter1));
  and2  gate555(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate556(.a(s_50), .O(gate187inter3));
  inv1  gate557(.a(s_51), .O(gate187inter4));
  nand2 gate558(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate559(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate560(.a(N65), .O(gate187inter7));
  inv1  gate561(.a(N708), .O(gate187inter8));
  nand2 gate562(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate563(.a(s_51), .b(gate187inter3), .O(gate187inter10));
  nor2  gate564(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate565(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate566(.a(gate187inter12), .b(gate187inter1), .O(N740));
xor2 gate188( .a(N69), .b(N709), .O(N741) );

  xor2  gate427(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate428(.a(gate189inter0), .b(s_32), .O(gate189inter1));
  and2  gate429(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate430(.a(s_32), .O(gate189inter3));
  inv1  gate431(.a(s_33), .O(gate189inter4));
  nand2 gate432(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate433(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate434(.a(N73), .O(gate189inter7));
  inv1  gate435(.a(N710), .O(gate189inter8));
  nand2 gate436(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate437(.a(s_33), .b(gate189inter3), .O(gate189inter10));
  nor2  gate438(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate439(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate440(.a(gate189inter12), .b(gate189inter1), .O(N742));
xor2 gate190( .a(N77), .b(N711), .O(N743) );

  xor2  gate525(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate526(.a(gate191inter0), .b(s_46), .O(gate191inter1));
  and2  gate527(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate528(.a(s_46), .O(gate191inter3));
  inv1  gate529(.a(s_47), .O(gate191inter4));
  nand2 gate530(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate531(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate532(.a(N81), .O(gate191inter7));
  inv1  gate533(.a(N712), .O(gate191inter8));
  nand2 gate534(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate535(.a(s_47), .b(gate191inter3), .O(gate191inter10));
  nor2  gate536(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate537(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate538(.a(gate191inter12), .b(gate191inter1), .O(N744));

  xor2  gate245(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate246(.a(gate192inter0), .b(s_6), .O(gate192inter1));
  and2  gate247(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate248(.a(s_6), .O(gate192inter3));
  inv1  gate249(.a(s_7), .O(gate192inter4));
  nand2 gate250(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate251(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate252(.a(N85), .O(gate192inter7));
  inv1  gate253(.a(N713), .O(gate192inter8));
  nand2 gate254(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate255(.a(s_7), .b(gate192inter3), .O(gate192inter10));
  nor2  gate256(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate257(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate258(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate413(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate414(.a(gate201inter0), .b(s_30), .O(gate201inter1));
  and2  gate415(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate416(.a(s_30), .O(gate201inter3));
  inv1  gate417(.a(s_31), .O(gate201inter4));
  nand2 gate418(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate419(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate420(.a(N121), .O(gate201inter7));
  inv1  gate421(.a(N722), .O(gate201inter8));
  nand2 gate422(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate423(.a(s_31), .b(gate201inter3), .O(gate201inter10));
  nor2  gate424(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate425(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate426(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule