module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12, gate679inter0, gate679inter1, gate679inter2, gate679inter3, gate679inter4, gate679inter5, gate679inter6, gate679inter7, gate679inter8, gate679inter9, gate679inter10, gate679inter11, gate679inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate552inter0, gate552inter1, gate552inter2, gate552inter3, gate552inter4, gate552inter5, gate552inter6, gate552inter7, gate552inter8, gate552inter9, gate552inter10, gate552inter11, gate552inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate541inter0, gate541inter1, gate541inter2, gate541inter3, gate541inter4, gate541inter5, gate541inter6, gate541inter7, gate541inter8, gate541inter9, gate541inter10, gate541inter11, gate541inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate351inter0, gate351inter1, gate351inter2, gate351inter3, gate351inter4, gate351inter5, gate351inter6, gate351inter7, gate351inter8, gate351inter9, gate351inter10, gate351inter11, gate351inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate843inter0, gate843inter1, gate843inter2, gate843inter3, gate843inter4, gate843inter5, gate843inter6, gate843inter7, gate843inter8, gate843inter9, gate843inter10, gate843inter11, gate843inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate760inter0, gate760inter1, gate760inter2, gate760inter3, gate760inter4, gate760inter5, gate760inter6, gate760inter7, gate760inter8, gate760inter9, gate760inter10, gate760inter11, gate760inter12, gate563inter0, gate563inter1, gate563inter2, gate563inter3, gate563inter4, gate563inter5, gate563inter6, gate563inter7, gate563inter8, gate563inter9, gate563inter10, gate563inter11, gate563inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate576inter0, gate576inter1, gate576inter2, gate576inter3, gate576inter4, gate576inter5, gate576inter6, gate576inter7, gate576inter8, gate576inter9, gate576inter10, gate576inter11, gate576inter12, gate858inter0, gate858inter1, gate858inter2, gate858inter3, gate858inter4, gate858inter5, gate858inter6, gate858inter7, gate858inter8, gate858inter9, gate858inter10, gate858inter11, gate858inter12, gate675inter0, gate675inter1, gate675inter2, gate675inter3, gate675inter4, gate675inter5, gate675inter6, gate675inter7, gate675inter8, gate675inter9, gate675inter10, gate675inter11, gate675inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate325inter0, gate325inter1, gate325inter2, gate325inter3, gate325inter4, gate325inter5, gate325inter6, gate325inter7, gate325inter8, gate325inter9, gate325inter10, gate325inter11, gate325inter12, gate517inter0, gate517inter1, gate517inter2, gate517inter3, gate517inter4, gate517inter5, gate517inter6, gate517inter7, gate517inter8, gate517inter9, gate517inter10, gate517inter11, gate517inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate318inter0, gate318inter1, gate318inter2, gate318inter3, gate318inter4, gate318inter5, gate318inter6, gate318inter7, gate318inter8, gate318inter9, gate318inter10, gate318inter11, gate318inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate861inter0, gate861inter1, gate861inter2, gate861inter3, gate861inter4, gate861inter5, gate861inter6, gate861inter7, gate861inter8, gate861inter9, gate861inter10, gate861inter11, gate861inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate649inter0, gate649inter1, gate649inter2, gate649inter3, gate649inter4, gate649inter5, gate649inter6, gate649inter7, gate649inter8, gate649inter9, gate649inter10, gate649inter11, gate649inter12, gate374inter0, gate374inter1, gate374inter2, gate374inter3, gate374inter4, gate374inter5, gate374inter6, gate374inter7, gate374inter8, gate374inter9, gate374inter10, gate374inter11, gate374inter12, gate807inter0, gate807inter1, gate807inter2, gate807inter3, gate807inter4, gate807inter5, gate807inter6, gate807inter7, gate807inter8, gate807inter9, gate807inter10, gate807inter11, gate807inter12, gate816inter0, gate816inter1, gate816inter2, gate816inter3, gate816inter4, gate816inter5, gate816inter6, gate816inter7, gate816inter8, gate816inter9, gate816inter10, gate816inter11, gate816inter12, gate775inter0, gate775inter1, gate775inter2, gate775inter3, gate775inter4, gate775inter5, gate775inter6, gate775inter7, gate775inter8, gate775inter9, gate775inter10, gate775inter11, gate775inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate616inter0, gate616inter1, gate616inter2, gate616inter3, gate616inter4, gate616inter5, gate616inter6, gate616inter7, gate616inter8, gate616inter9, gate616inter10, gate616inter11, gate616inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate817inter0, gate817inter1, gate817inter2, gate817inter3, gate817inter4, gate817inter5, gate817inter6, gate817inter7, gate817inter8, gate817inter9, gate817inter10, gate817inter11, gate817inter12, gate623inter0, gate623inter1, gate623inter2, gate623inter3, gate623inter4, gate623inter5, gate623inter6, gate623inter7, gate623inter8, gate623inter9, gate623inter10, gate623inter11, gate623inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate794inter0, gate794inter1, gate794inter2, gate794inter3, gate794inter4, gate794inter5, gate794inter6, gate794inter7, gate794inter8, gate794inter9, gate794inter10, gate794inter11, gate794inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate780inter0, gate780inter1, gate780inter2, gate780inter3, gate780inter4, gate780inter5, gate780inter6, gate780inter7, gate780inter8, gate780inter9, gate780inter10, gate780inter11, gate780inter12, gate789inter0, gate789inter1, gate789inter2, gate789inter3, gate789inter4, gate789inter5, gate789inter6, gate789inter7, gate789inter8, gate789inter9, gate789inter10, gate789inter11, gate789inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate350inter0, gate350inter1, gate350inter2, gate350inter3, gate350inter4, gate350inter5, gate350inter6, gate350inter7, gate350inter8, gate350inter9, gate350inter10, gate350inter11, gate350inter12, gate600inter0, gate600inter1, gate600inter2, gate600inter3, gate600inter4, gate600inter5, gate600inter6, gate600inter7, gate600inter8, gate600inter9, gate600inter10, gate600inter11, gate600inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate340inter0, gate340inter1, gate340inter2, gate340inter3, gate340inter4, gate340inter5, gate340inter6, gate340inter7, gate340inter8, gate340inter9, gate340inter10, gate340inter11, gate340inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate361inter0, gate361inter1, gate361inter2, gate361inter3, gate361inter4, gate361inter5, gate361inter6, gate361inter7, gate361inter8, gate361inter9, gate361inter10, gate361inter11, gate361inter12, gate665inter0, gate665inter1, gate665inter2, gate665inter3, gate665inter4, gate665inter5, gate665inter6, gate665inter7, gate665inter8, gate665inter9, gate665inter10, gate665inter11, gate665inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate324inter0, gate324inter1, gate324inter2, gate324inter3, gate324inter4, gate324inter5, gate324inter6, gate324inter7, gate324inter8, gate324inter9, gate324inter10, gate324inter11, gate324inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate570inter0, gate570inter1, gate570inter2, gate570inter3, gate570inter4, gate570inter5, gate570inter6, gate570inter7, gate570inter8, gate570inter9, gate570inter10, gate570inter11, gate570inter12, gate621inter0, gate621inter1, gate621inter2, gate621inter3, gate621inter4, gate621inter5, gate621inter6, gate621inter7, gate621inter8, gate621inter9, gate621inter10, gate621inter11, gate621inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate663inter0, gate663inter1, gate663inter2, gate663inter3, gate663inter4, gate663inter5, gate663inter6, gate663inter7, gate663inter8, gate663inter9, gate663inter10, gate663inter11, gate663inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate767inter0, gate767inter1, gate767inter2, gate767inter3, gate767inter4, gate767inter5, gate767inter6, gate767inter7, gate767inter8, gate767inter9, gate767inter10, gate767inter11, gate767inter12, gate639inter0, gate639inter1, gate639inter2, gate639inter3, gate639inter4, gate639inter5, gate639inter6, gate639inter7, gate639inter8, gate639inter9, gate639inter10, gate639inter11, gate639inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate686inter0, gate686inter1, gate686inter2, gate686inter3, gate686inter4, gate686inter5, gate686inter6, gate686inter7, gate686inter8, gate686inter9, gate686inter10, gate686inter11, gate686inter12, gate624inter0, gate624inter1, gate624inter2, gate624inter3, gate624inter4, gate624inter5, gate624inter6, gate624inter7, gate624inter8, gate624inter9, gate624inter10, gate624inter11, gate624inter12, gate572inter0, gate572inter1, gate572inter2, gate572inter3, gate572inter4, gate572inter5, gate572inter6, gate572inter7, gate572inter8, gate572inter9, gate572inter10, gate572inter11, gate572inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate804inter0, gate804inter1, gate804inter2, gate804inter3, gate804inter4, gate804inter5, gate804inter6, gate804inter7, gate804inter8, gate804inter9, gate804inter10, gate804inter11, gate804inter12, gate835inter0, gate835inter1, gate835inter2, gate835inter3, gate835inter4, gate835inter5, gate835inter6, gate835inter7, gate835inter8, gate835inter9, gate835inter10, gate835inter11, gate835inter12, gate681inter0, gate681inter1, gate681inter2, gate681inter3, gate681inter4, gate681inter5, gate681inter6, gate681inter7, gate681inter8, gate681inter9, gate681inter10, gate681inter11, gate681inter12, gate329inter0, gate329inter1, gate329inter2, gate329inter3, gate329inter4, gate329inter5, gate329inter6, gate329inter7, gate329inter8, gate329inter9, gate329inter10, gate329inter11, gate329inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate368inter0, gate368inter1, gate368inter2, gate368inter3, gate368inter4, gate368inter5, gate368inter6, gate368inter7, gate368inter8, gate368inter9, gate368inter10, gate368inter11, gate368inter12, gate864inter0, gate864inter1, gate864inter2, gate864inter3, gate864inter4, gate864inter5, gate864inter6, gate864inter7, gate864inter8, gate864inter9, gate864inter10, gate864inter11, gate864inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate766inter0, gate766inter1, gate766inter2, gate766inter3, gate766inter4, gate766inter5, gate766inter6, gate766inter7, gate766inter8, gate766inter9, gate766inter10, gate766inter11, gate766inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate863inter0, gate863inter1, gate863inter2, gate863inter3, gate863inter4, gate863inter5, gate863inter6, gate863inter7, gate863inter8, gate863inter9, gate863inter10, gate863inter11, gate863inter12, gate669inter0, gate669inter1, gate669inter2, gate669inter3, gate669inter4, gate669inter5, gate669inter6, gate669inter7, gate669inter8, gate669inter9, gate669inter10, gate669inter11, gate669inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate676inter0, gate676inter1, gate676inter2, gate676inter3, gate676inter4, gate676inter5, gate676inter6, gate676inter7, gate676inter8, gate676inter9, gate676inter10, gate676inter11, gate676inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate841inter0, gate841inter1, gate841inter2, gate841inter3, gate841inter4, gate841inter5, gate841inter6, gate841inter7, gate841inter8, gate841inter9, gate841inter10, gate841inter11, gate841inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate534inter0, gate534inter1, gate534inter2, gate534inter3, gate534inter4, gate534inter5, gate534inter6, gate534inter7, gate534inter8, gate534inter9, gate534inter10, gate534inter11, gate534inter12, gate516inter0, gate516inter1, gate516inter2, gate516inter3, gate516inter4, gate516inter5, gate516inter6, gate516inter7, gate516inter8, gate516inter9, gate516inter10, gate516inter11, gate516inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate851inter0, gate851inter1, gate851inter2, gate851inter3, gate851inter4, gate851inter5, gate851inter6, gate851inter7, gate851inter8, gate851inter9, gate851inter10, gate851inter11, gate851inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate304inter0, gate304inter1, gate304inter2, gate304inter3, gate304inter4, gate304inter5, gate304inter6, gate304inter7, gate304inter8, gate304inter9, gate304inter10, gate304inter11, gate304inter12, gate683inter0, gate683inter1, gate683inter2, gate683inter3, gate683inter4, gate683inter5, gate683inter6, gate683inter7, gate683inter8, gate683inter9, gate683inter10, gate683inter11, gate683inter12, gate637inter0, gate637inter1, gate637inter2, gate637inter3, gate637inter4, gate637inter5, gate637inter6, gate637inter7, gate637inter8, gate637inter9, gate637inter10, gate637inter11, gate637inter12, gate800inter0, gate800inter1, gate800inter2, gate800inter3, gate800inter4, gate800inter5, gate800inter6, gate800inter7, gate800inter8, gate800inter9, gate800inter10, gate800inter11, gate800inter12, gate750inter0, gate750inter1, gate750inter2, gate750inter3, gate750inter4, gate750inter5, gate750inter6, gate750inter7, gate750inter8, gate750inter9, gate750inter10, gate750inter11, gate750inter12, gate786inter0, gate786inter1, gate786inter2, gate786inter3, gate786inter4, gate786inter5, gate786inter6, gate786inter7, gate786inter8, gate786inter9, gate786inter10, gate786inter11, gate786inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate528inter0, gate528inter1, gate528inter2, gate528inter3, gate528inter4, gate528inter5, gate528inter6, gate528inter7, gate528inter8, gate528inter9, gate528inter10, gate528inter11, gate528inter12, gate536inter0, gate536inter1, gate536inter2, gate536inter3, gate536inter4, gate536inter5, gate536inter6, gate536inter7, gate536inter8, gate536inter9, gate536inter10, gate536inter11, gate536inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate526inter0, gate526inter1, gate526inter2, gate526inter3, gate526inter4, gate526inter5, gate526inter6, gate526inter7, gate526inter8, gate526inter9, gate526inter10, gate526inter11, gate526inter12, gate820inter0, gate820inter1, gate820inter2, gate820inter3, gate820inter4, gate820inter5, gate820inter6, gate820inter7, gate820inter8, gate820inter9, gate820inter10, gate820inter11, gate820inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate650inter0, gate650inter1, gate650inter2, gate650inter3, gate650inter4, gate650inter5, gate650inter6, gate650inter7, gate650inter8, gate650inter9, gate650inter10, gate650inter11, gate650inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate550inter0, gate550inter1, gate550inter2, gate550inter3, gate550inter4, gate550inter5, gate550inter6, gate550inter7, gate550inter8, gate550inter9, gate550inter10, gate550inter11, gate550inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate837inter0, gate837inter1, gate837inter2, gate837inter3, gate837inter4, gate837inter5, gate837inter6, gate837inter7, gate837inter8, gate837inter9, gate837inter10, gate837inter11, gate837inter12, gate822inter0, gate822inter1, gate822inter2, gate822inter3, gate822inter4, gate822inter5, gate822inter6, gate822inter7, gate822inter8, gate822inter9, gate822inter10, gate822inter11, gate822inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate636inter0, gate636inter1, gate636inter2, gate636inter3, gate636inter4, gate636inter5, gate636inter6, gate636inter7, gate636inter8, gate636inter9, gate636inter10, gate636inter11, gate636inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12, gate796inter0, gate796inter1, gate796inter2, gate796inter3, gate796inter4, gate796inter5, gate796inter6, gate796inter7, gate796inter8, gate796inter9, gate796inter10, gate796inter11, gate796inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate812inter0, gate812inter1, gate812inter2, gate812inter3, gate812inter4, gate812inter5, gate812inter6, gate812inter7, gate812inter8, gate812inter9, gate812inter10, gate812inter11, gate812inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate353inter0, gate353inter1, gate353inter2, gate353inter3, gate353inter4, gate353inter5, gate353inter6, gate353inter7, gate353inter8, gate353inter9, gate353inter10, gate353inter11, gate353inter12, gate852inter0, gate852inter1, gate852inter2, gate852inter3, gate852inter4, gate852inter5, gate852inter6, gate852inter7, gate852inter8, gate852inter9, gate852inter10, gate852inter11, gate852inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate801inter0, gate801inter1, gate801inter2, gate801inter3, gate801inter4, gate801inter5, gate801inter6, gate801inter7, gate801inter8, gate801inter9, gate801inter10, gate801inter11, gate801inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate673inter0, gate673inter1, gate673inter2, gate673inter3, gate673inter4, gate673inter5, gate673inter6, gate673inter7, gate673inter8, gate673inter9, gate673inter10, gate673inter11, gate673inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate357inter0, gate357inter1, gate357inter2, gate357inter3, gate357inter4, gate357inter5, gate357inter6, gate357inter7, gate357inter8, gate357inter9, gate357inter10, gate357inter11, gate357inter12, gate378inter0, gate378inter1, gate378inter2, gate378inter3, gate378inter4, gate378inter5, gate378inter6, gate378inter7, gate378inter8, gate378inter9, gate378inter10, gate378inter11, gate378inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate828inter0, gate828inter1, gate828inter2, gate828inter3, gate828inter4, gate828inter5, gate828inter6, gate828inter7, gate828inter8, gate828inter9, gate828inter10, gate828inter11, gate828inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate850inter0, gate850inter1, gate850inter2, gate850inter3, gate850inter4, gate850inter5, gate850inter6, gate850inter7, gate850inter8, gate850inter9, gate850inter10, gate850inter11, gate850inter12, gate765inter0, gate765inter1, gate765inter2, gate765inter3, gate765inter4, gate765inter5, gate765inter6, gate765inter7, gate765inter8, gate765inter9, gate765inter10, gate765inter11, gate765inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );

  xor2  gate1511(.a(N91), .b(N66), .O(gate18inter0));
  nand2 gate1512(.a(gate18inter0), .b(s_90), .O(gate18inter1));
  and2  gate1513(.a(N91), .b(N66), .O(gate18inter2));
  inv1  gate1514(.a(s_90), .O(gate18inter3));
  inv1  gate1515(.a(s_91), .O(gate18inter4));
  nand2 gate1516(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1517(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1518(.a(N66), .O(gate18inter7));
  inv1  gate1519(.a(N91), .O(gate18inter8));
  nand2 gate1520(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1521(.a(s_91), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1522(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1523(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1524(.a(gate18inter12), .b(gate18inter1), .O(N252));
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );

  xor2  gate1329(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate1330(.a(gate77inter0), .b(s_64), .O(gate77inter1));
  and2  gate1331(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate1332(.a(s_64), .O(gate77inter3));
  inv1  gate1333(.a(s_65), .O(gate77inter4));
  nand2 gate1334(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1335(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1336(.a(N306), .O(gate77inter7));
  inv1  gate1337(.a(N331), .O(gate77inter8));
  nand2 gate1338(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1339(.a(s_65), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1340(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1341(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1342(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );

  xor2  gate2253(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate2254(.a(gate79inter0), .b(s_196), .O(gate79inter1));
  and2  gate2255(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate2256(.a(s_196), .O(gate79inter3));
  inv1  gate2257(.a(s_197), .O(gate79inter4));
  nand2 gate2258(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2259(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2260(.a(N306), .O(gate79inter7));
  inv1  gate2261(.a(N331), .O(gate79inter8));
  nand2 gate2262(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2263(.a(s_197), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2264(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2265(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2266(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );

  xor2  gate1413(.a(N280), .b(N326), .O(gate97inter0));
  nand2 gate1414(.a(gate97inter0), .b(s_76), .O(gate97inter1));
  and2  gate1415(.a(N280), .b(N326), .O(gate97inter2));
  inv1  gate1416(.a(s_76), .O(gate97inter3));
  inv1  gate1417(.a(s_77), .O(gate97inter4));
  nand2 gate1418(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1419(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1420(.a(N326), .O(gate97inter7));
  inv1  gate1421(.a(N280), .O(gate97inter8));
  nand2 gate1422(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1423(.a(s_77), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1424(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1425(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1426(.a(gate97inter12), .b(gate97inter1), .O(N602));

  xor2  gate951(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate952(.a(gate98inter0), .b(s_10), .O(gate98inter1));
  and2  gate953(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate954(.a(s_10), .O(gate98inter3));
  inv1  gate955(.a(s_11), .O(gate98inter4));
  nand2 gate956(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate957(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate958(.a(N260), .O(gate98inter7));
  inv1  gate959(.a(N72), .O(gate98inter8));
  nand2 gate960(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate961(.a(s_11), .b(gate98inter3), .O(gate98inter10));
  nor2  gate962(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate963(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate964(.a(gate98inter12), .b(gate98inter1), .O(N603));

  xor2  gate3303(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate3304(.a(gate99inter0), .b(s_346), .O(gate99inter1));
  and2  gate3305(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate3306(.a(s_346), .O(gate99inter3));
  inv1  gate3307(.a(s_347), .O(gate99inter4));
  nand2 gate3308(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate3309(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate3310(.a(N260), .O(gate99inter7));
  inv1  gate3311(.a(N300), .O(gate99inter8));
  nand2 gate3312(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate3313(.a(s_347), .b(gate99inter3), .O(gate99inter10));
  nor2  gate3314(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate3315(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate3316(.a(gate99inter12), .b(gate99inter1), .O(N608));
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );

  xor2  gate2169(.a(N612), .b(N53), .O(gate160inter0));
  nand2 gate2170(.a(gate160inter0), .b(s_184), .O(gate160inter1));
  and2  gate2171(.a(N612), .b(N53), .O(gate160inter2));
  inv1  gate2172(.a(s_184), .O(gate160inter3));
  inv1  gate2173(.a(s_185), .O(gate160inter4));
  nand2 gate2174(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2175(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2176(.a(N53), .O(gate160inter7));
  inv1  gate2177(.a(N612), .O(gate160inter8));
  nand2 gate2178(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2179(.a(s_185), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2180(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2181(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2182(.a(gate160inter12), .b(gate160inter1), .O(N899));

  xor2  gate2323(.a(N608), .b(N60), .O(gate161inter0));
  nand2 gate2324(.a(gate161inter0), .b(s_206), .O(gate161inter1));
  and2  gate2325(.a(N608), .b(N60), .O(gate161inter2));
  inv1  gate2326(.a(s_206), .O(gate161inter3));
  inv1  gate2327(.a(s_207), .O(gate161inter4));
  nand2 gate2328(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2329(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2330(.a(N60), .O(gate161inter7));
  inv1  gate2331(.a(N608), .O(gate161inter8));
  nand2 gate2332(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2333(.a(s_207), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2334(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2335(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2336(.a(gate161inter12), .b(gate161inter1), .O(N903));
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );

  xor2  gate3219(.a(N889), .b(N616), .O(gate234inter0));
  nand2 gate3220(.a(gate234inter0), .b(s_334), .O(gate234inter1));
  and2  gate3221(.a(N889), .b(N616), .O(gate234inter2));
  inv1  gate3222(.a(s_334), .O(gate234inter3));
  inv1  gate3223(.a(s_335), .O(gate234inter4));
  nand2 gate3224(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate3225(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate3226(.a(N616), .O(gate234inter7));
  inv1  gate3227(.a(N889), .O(gate234inter8));
  nand2 gate3228(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate3229(.a(s_335), .b(gate234inter3), .O(gate234inter10));
  nor2  gate3230(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate3231(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate3232(.a(gate234inter12), .b(gate234inter1), .O(N1055));

  xor2  gate1203(.a(N890), .b(N625), .O(gate235inter0));
  nand2 gate1204(.a(gate235inter0), .b(s_46), .O(gate235inter1));
  and2  gate1205(.a(N890), .b(N625), .O(gate235inter2));
  inv1  gate1206(.a(s_46), .O(gate235inter3));
  inv1  gate1207(.a(s_47), .O(gate235inter4));
  nand2 gate1208(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1209(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1210(.a(N625), .O(gate235inter7));
  inv1  gate1211(.a(N890), .O(gate235inter8));
  nand2 gate1212(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1213(.a(s_47), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1214(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1215(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1216(.a(gate235inter12), .b(gate235inter1), .O(N1063));

  xor2  gate1273(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate1274(.a(gate236inter0), .b(s_56), .O(gate236inter1));
  and2  gate1275(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate1276(.a(s_56), .O(gate236inter3));
  inv1  gate1277(.a(s_57), .O(gate236inter4));
  nand2 gate1278(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1279(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1280(.a(N622), .O(gate236inter7));
  inv1  gate1281(.a(N891), .O(gate236inter8));
  nand2 gate1282(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1283(.a(s_57), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1284(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1285(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1286(.a(gate236inter12), .b(gate236inter1), .O(N1064));
nand2 gate237( .a(N655), .b(N895), .O(N1067) );

  xor2  gate2099(.a(N896), .b(N652), .O(gate238inter0));
  nand2 gate2100(.a(gate238inter0), .b(s_174), .O(gate238inter1));
  and2  gate2101(.a(N896), .b(N652), .O(gate238inter2));
  inv1  gate2102(.a(s_174), .O(gate238inter3));
  inv1  gate2103(.a(s_175), .O(gate238inter4));
  nand2 gate2104(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2105(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2106(.a(N652), .O(gate238inter7));
  inv1  gate2107(.a(N896), .O(gate238inter8));
  nand2 gate2108(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2109(.a(s_175), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2110(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2111(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2112(.a(gate238inter12), .b(gate238inter1), .O(N1068));
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );

  xor2  gate1595(.a(N991), .b(N727), .O(gate241inter0));
  nand2 gate1596(.a(gate241inter0), .b(s_102), .O(gate241inter1));
  and2  gate1597(.a(N991), .b(N727), .O(gate241inter2));
  inv1  gate1598(.a(s_102), .O(gate241inter3));
  inv1  gate1599(.a(s_103), .O(gate241inter4));
  nand2 gate1600(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1601(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1602(.a(N727), .O(gate241inter7));
  inv1  gate1603(.a(N991), .O(gate241inter8));
  nand2 gate1604(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1605(.a(s_103), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1606(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1607(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1608(.a(gate241inter12), .b(gate241inter1), .O(N1121));

  xor2  gate3443(.a(N992), .b(N724), .O(gate242inter0));
  nand2 gate3444(.a(gate242inter0), .b(s_366), .O(gate242inter1));
  and2  gate3445(.a(N992), .b(N724), .O(gate242inter2));
  inv1  gate3446(.a(s_366), .O(gate242inter3));
  inv1  gate3447(.a(s_367), .O(gate242inter4));
  nand2 gate3448(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate3449(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate3450(.a(N724), .O(gate242inter7));
  inv1  gate3451(.a(N992), .O(gate242inter8));
  nand2 gate3452(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate3453(.a(s_367), .b(gate242inter3), .O(gate242inter10));
  nor2  gate3454(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate3455(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate3456(.a(gate242inter12), .b(gate242inter1), .O(N1122));

  xor2  gate3177(.a(N1002), .b(N739), .O(gate243inter0));
  nand2 gate3178(.a(gate243inter0), .b(s_328), .O(gate243inter1));
  and2  gate3179(.a(N1002), .b(N739), .O(gate243inter2));
  inv1  gate3180(.a(s_328), .O(gate243inter3));
  inv1  gate3181(.a(s_329), .O(gate243inter4));
  nand2 gate3182(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate3183(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate3184(.a(N739), .O(gate243inter7));
  inv1  gate3185(.a(N1002), .O(gate243inter8));
  nand2 gate3186(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate3187(.a(s_329), .b(gate243inter3), .O(gate243inter10));
  nor2  gate3188(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate3189(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate3190(.a(gate243inter12), .b(gate243inter1), .O(N1128));
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );

  xor2  gate1063(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate1064(.a(gate245inter0), .b(s_26), .O(gate245inter1));
  and2  gate1065(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate1066(.a(s_26), .O(gate245inter3));
  inv1  gate1067(.a(s_27), .O(gate245inter4));
  nand2 gate1068(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1069(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1070(.a(N745), .O(gate245inter7));
  inv1  gate1071(.a(N1005), .O(gate245inter8));
  nand2 gate1072(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1073(.a(s_27), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1074(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1075(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1076(.a(gate245inter12), .b(gate245inter1), .O(N1130));

  xor2  gate3415(.a(N1006), .b(N742), .O(gate246inter0));
  nand2 gate3416(.a(gate246inter0), .b(s_362), .O(gate246inter1));
  and2  gate3417(.a(N1006), .b(N742), .O(gate246inter2));
  inv1  gate3418(.a(s_362), .O(gate246inter3));
  inv1  gate3419(.a(s_363), .O(gate246inter4));
  nand2 gate3420(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate3421(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate3422(.a(N742), .O(gate246inter7));
  inv1  gate3423(.a(N1006), .O(gate246inter8));
  nand2 gate3424(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate3425(.a(s_363), .b(gate246inter3), .O(gate246inter10));
  nor2  gate3426(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate3427(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate3428(.a(gate246inter12), .b(gate246inter1), .O(N1131));

  xor2  gate3023(.a(N1008), .b(N751), .O(gate247inter0));
  nand2 gate3024(.a(gate247inter0), .b(s_306), .O(gate247inter1));
  and2  gate3025(.a(N1008), .b(N751), .O(gate247inter2));
  inv1  gate3026(.a(s_306), .O(gate247inter3));
  inv1  gate3027(.a(s_307), .O(gate247inter4));
  nand2 gate3028(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate3029(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate3030(.a(N751), .O(gate247inter7));
  inv1  gate3031(.a(N1008), .O(gate247inter8));
  nand2 gate3032(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate3033(.a(s_307), .b(gate247inter3), .O(gate247inter10));
  nor2  gate3034(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate3035(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate3036(.a(gate247inter12), .b(gate247inter1), .O(N1132));
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );

  xor2  gate2295(.a(N892), .b(N985), .O(gate261inter0));
  nand2 gate2296(.a(gate261inter0), .b(s_202), .O(gate261inter1));
  and2  gate2297(.a(N892), .b(N985), .O(gate261inter2));
  inv1  gate2298(.a(s_202), .O(gate261inter3));
  inv1  gate2299(.a(s_203), .O(gate261inter4));
  nand2 gate2300(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2301(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2302(.a(N985), .O(gate261inter7));
  inv1  gate2303(.a(N892), .O(gate261inter8));
  nand2 gate2304(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2305(.a(s_203), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2306(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2307(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2308(.a(gate261inter12), .b(gate261inter1), .O(N1160));
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate895(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate896(.a(gate275inter0), .b(s_2), .O(gate275inter1));
  and2  gate897(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate898(.a(s_2), .O(gate275inter3));
  inv1  gate899(.a(s_3), .O(gate275inter4));
  nand2 gate900(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate901(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate902(.a(N1016), .O(gate275inter7));
  inv1  gate903(.a(N946), .O(gate275inter8));
  nand2 gate904(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate905(.a(s_3), .b(gate275inter3), .O(gate275inter10));
  nor2  gate906(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate907(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate908(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );

  xor2  gate1077(.a(N954), .b(N1022), .O(gate279inter0));
  nand2 gate1078(.a(gate279inter0), .b(s_28), .O(gate279inter1));
  and2  gate1079(.a(N954), .b(N1022), .O(gate279inter2));
  inv1  gate1080(.a(s_28), .O(gate279inter3));
  inv1  gate1081(.a(s_29), .O(gate279inter4));
  nand2 gate1082(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1083(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1084(.a(N1022), .O(gate279inter7));
  inv1  gate1085(.a(N954), .O(gate279inter8));
  nand2 gate1086(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1087(.a(s_29), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1088(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1089(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1090(.a(gate279inter12), .b(gate279inter1), .O(N1214));
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );

  xor2  gate2211(.a(N972), .b(N1037), .O(gate289inter0));
  nand2 gate2212(.a(gate289inter0), .b(s_190), .O(gate289inter1));
  and2  gate2213(.a(N972), .b(N1037), .O(gate289inter2));
  inv1  gate2214(.a(s_190), .O(gate289inter3));
  inv1  gate2215(.a(s_191), .O(gate289inter4));
  nand2 gate2216(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2217(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2218(.a(N1037), .O(gate289inter7));
  inv1  gate2219(.a(N972), .O(gate289inter8));
  nand2 gate2220(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2221(.a(s_191), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2222(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2223(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2224(.a(gate289inter12), .b(gate289inter1), .O(N1224));
inv1 gate290( .a(N1040), .O(N1225) );

  xor2  gate1371(.a(N976), .b(N1040), .O(gate291inter0));
  nand2 gate1372(.a(gate291inter0), .b(s_70), .O(gate291inter1));
  and2  gate1373(.a(N976), .b(N1040), .O(gate291inter2));
  inv1  gate1374(.a(s_70), .O(gate291inter3));
  inv1  gate1375(.a(s_71), .O(gate291inter4));
  nand2 gate1376(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1377(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1378(.a(N1040), .O(gate291inter7));
  inv1  gate1379(.a(N976), .O(gate291inter8));
  nand2 gate1380(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1381(.a(s_71), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1382(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1383(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1384(.a(gate291inter12), .b(gate291inter1), .O(N1226));
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );

  xor2  gate1525(.a(N980), .b(N1043), .O(gate294inter0));
  nand2 gate1526(.a(gate294inter0), .b(s_92), .O(gate294inter1));
  and2  gate1527(.a(N980), .b(N1043), .O(gate294inter2));
  inv1  gate1528(.a(s_92), .O(gate294inter3));
  inv1  gate1529(.a(s_93), .O(gate294inter4));
  nand2 gate1530(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1531(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1532(.a(N1043), .O(gate294inter7));
  inv1  gate1533(.a(N980), .O(gate294inter8));
  nand2 gate1534(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1535(.a(s_93), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1536(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1537(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1538(.a(gate294inter12), .b(gate294inter1), .O(N1229));
inv1 gate295( .a(N981), .O(N1230) );

  xor2  gate2071(.a(N984), .b(N981), .O(gate296inter0));
  nand2 gate2072(.a(gate296inter0), .b(s_170), .O(gate296inter1));
  and2  gate2073(.a(N984), .b(N981), .O(gate296inter2));
  inv1  gate2074(.a(s_170), .O(gate296inter3));
  inv1  gate2075(.a(s_171), .O(gate296inter4));
  nand2 gate2076(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2077(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2078(.a(N981), .O(gate296inter7));
  inv1  gate2079(.a(N984), .O(gate296inter8));
  nand2 gate2080(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2081(.a(s_171), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2082(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2083(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2084(.a(gate296inter12), .b(gate296inter1), .O(N1231));
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );

  xor2  gate1707(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate1708(.a(gate298inter0), .b(s_118), .O(gate298inter1));
  and2  gate1709(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate1710(.a(s_118), .O(gate298inter3));
  inv1  gate1711(.a(s_119), .O(gate298inter4));
  nand2 gate1712(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate1713(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate1714(.a(N1121), .O(gate298inter7));
  inv1  gate1715(.a(N1122), .O(gate298inter8));
  nand2 gate1716(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate1717(.a(s_119), .b(gate298inter3), .O(gate298inter10));
  nor2  gate1718(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate1719(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate1720(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );

  xor2  gate1861(.a(N997), .b(N1046), .O(gate300inter0));
  nand2 gate1862(.a(gate300inter0), .b(s_140), .O(gate300inter1));
  and2  gate1863(.a(N997), .b(N1046), .O(gate300inter2));
  inv1  gate1864(.a(s_140), .O(gate300inter3));
  inv1  gate1865(.a(s_141), .O(gate300inter4));
  nand2 gate1866(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate1867(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate1868(.a(N1046), .O(gate300inter7));
  inv1  gate1869(.a(N997), .O(gate300inter8));
  nand2 gate1870(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate1871(.a(s_141), .b(gate300inter3), .O(gate300inter10));
  nor2  gate1872(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate1873(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate1874(.a(gate300inter12), .b(gate300inter1), .O(N1239));
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );

  xor2  gate2757(.a(N1129), .b(N1128), .O(gate304inter0));
  nand2 gate2758(.a(gate304inter0), .b(s_268), .O(gate304inter1));
  and2  gate2759(.a(N1129), .b(N1128), .O(gate304inter2));
  inv1  gate2760(.a(s_268), .O(gate304inter3));
  inv1  gate2761(.a(s_269), .O(gate304inter4));
  nand2 gate2762(.a(gate304inter4), .b(gate304inter3), .O(gate304inter5));
  nor2  gate2763(.a(gate304inter5), .b(gate304inter2), .O(gate304inter6));
  inv1  gate2764(.a(N1128), .O(gate304inter7));
  inv1  gate2765(.a(N1129), .O(gate304inter8));
  nand2 gate2766(.a(gate304inter8), .b(gate304inter7), .O(gate304inter9));
  nand2 gate2767(.a(s_269), .b(gate304inter3), .O(gate304inter10));
  nor2  gate2768(.a(gate304inter10), .b(gate304inter9), .O(gate304inter11));
  nor2  gate2769(.a(gate304inter11), .b(gate304inter6), .O(gate304inter12));
  nand2 gate2770(.a(gate304inter12), .b(gate304inter1), .O(N1243));
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate2883(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate2884(.a(gate312inter0), .b(s_286), .O(gate312inter1));
  and2  gate2885(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate2886(.a(s_286), .O(gate312inter3));
  inv1  gate2887(.a(s_287), .O(gate312inter4));
  nand2 gate2888(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate2889(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate2890(.a(N631), .O(gate312inter7));
  inv1  gate2891(.a(N1159), .O(gate312inter8));
  nand2 gate2892(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate2893(.a(s_287), .b(gate312inter3), .O(gate312inter10));
  nor2  gate2894(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate2895(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate2896(.a(gate312inter12), .b(gate312inter1), .O(N1267));

  xor2  gate2421(.a(N1205), .b(N688), .O(gate313inter0));
  nand2 gate2422(.a(gate313inter0), .b(s_220), .O(gate313inter1));
  and2  gate2423(.a(N1205), .b(N688), .O(gate313inter2));
  inv1  gate2424(.a(s_220), .O(gate313inter3));
  inv1  gate2425(.a(s_221), .O(gate313inter4));
  nand2 gate2426(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate2427(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate2428(.a(N688), .O(gate313inter7));
  inv1  gate2429(.a(N1205), .O(gate313inter8));
  nand2 gate2430(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate2431(.a(s_221), .b(gate313inter3), .O(gate313inter10));
  nor2  gate2432(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate2433(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate2434(.a(gate313inter12), .b(gate313inter1), .O(N1309));
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );

  xor2  gate1357(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate1358(.a(gate316inter0), .b(s_68), .O(gate316inter1));
  and2  gate1359(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate1360(.a(s_68), .O(gate316inter3));
  inv1  gate1361(.a(s_69), .O(gate316inter4));
  nand2 gate1362(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate1363(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate1364(.a(N697), .O(gate316inter7));
  inv1  gate1365(.a(N1211), .O(gate316inter8));
  nand2 gate1366(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate1367(.a(s_69), .b(gate316inter3), .O(gate316inter10));
  nor2  gate1368(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate1369(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate1370(.a(gate316inter12), .b(gate316inter1), .O(N1312));

  xor2  gate993(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate994(.a(gate317inter0), .b(s_16), .O(gate317inter1));
  and2  gate995(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate996(.a(s_16), .O(gate317inter3));
  inv1  gate997(.a(s_17), .O(gate317inter4));
  nand2 gate998(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate999(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate1000(.a(N700), .O(gate317inter7));
  inv1  gate1001(.a(N1213), .O(gate317inter8));
  nand2 gate1002(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate1003(.a(s_17), .b(gate317inter3), .O(gate317inter10));
  nor2  gate1004(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate1005(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate1006(.a(gate317inter12), .b(gate317inter1), .O(N1313));

  xor2  gate1427(.a(N1215), .b(N703), .O(gate318inter0));
  nand2 gate1428(.a(gate318inter0), .b(s_78), .O(gate318inter1));
  and2  gate1429(.a(N1215), .b(N703), .O(gate318inter2));
  inv1  gate1430(.a(s_78), .O(gate318inter3));
  inv1  gate1431(.a(s_79), .O(gate318inter4));
  nand2 gate1432(.a(gate318inter4), .b(gate318inter3), .O(gate318inter5));
  nor2  gate1433(.a(gate318inter5), .b(gate318inter2), .O(gate318inter6));
  inv1  gate1434(.a(N703), .O(gate318inter7));
  inv1  gate1435(.a(N1215), .O(gate318inter8));
  nand2 gate1436(.a(gate318inter8), .b(gate318inter7), .O(gate318inter9));
  nand2 gate1437(.a(s_79), .b(gate318inter3), .O(gate318inter10));
  nor2  gate1438(.a(gate318inter10), .b(gate318inter9), .O(gate318inter11));
  nor2  gate1439(.a(gate318inter11), .b(gate318inter6), .O(gate318inter12));
  nand2 gate1440(.a(gate318inter12), .b(gate318inter1), .O(N1314));
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );

  xor2  gate2155(.a(N1230), .b(N628), .O(gate324inter0));
  nand2 gate2156(.a(gate324inter0), .b(s_182), .O(gate324inter1));
  and2  gate2157(.a(N1230), .b(N628), .O(gate324inter2));
  inv1  gate2158(.a(s_182), .O(gate324inter3));
  inv1  gate2159(.a(s_183), .O(gate324inter4));
  nand2 gate2160(.a(gate324inter4), .b(gate324inter3), .O(gate324inter5));
  nor2  gate2161(.a(gate324inter5), .b(gate324inter2), .O(gate324inter6));
  inv1  gate2162(.a(N628), .O(gate324inter7));
  inv1  gate2163(.a(N1230), .O(gate324inter8));
  nand2 gate2164(.a(gate324inter8), .b(gate324inter7), .O(gate324inter9));
  nand2 gate2165(.a(s_183), .b(gate324inter3), .O(gate324inter10));
  nor2  gate2166(.a(gate324inter10), .b(gate324inter9), .O(gate324inter11));
  nor2  gate2167(.a(gate324inter11), .b(gate324inter6), .O(gate324inter12));
  nand2 gate2168(.a(gate324inter12), .b(gate324inter1), .O(N1322));

  xor2  gate1287(.a(N1238), .b(N730), .O(gate325inter0));
  nand2 gate1288(.a(gate325inter0), .b(s_58), .O(gate325inter1));
  and2  gate1289(.a(N1238), .b(N730), .O(gate325inter2));
  inv1  gate1290(.a(s_58), .O(gate325inter3));
  inv1  gate1291(.a(s_59), .O(gate325inter4));
  nand2 gate1292(.a(gate325inter4), .b(gate325inter3), .O(gate325inter5));
  nor2  gate1293(.a(gate325inter5), .b(gate325inter2), .O(gate325inter6));
  inv1  gate1294(.a(N730), .O(gate325inter7));
  inv1  gate1295(.a(N1238), .O(gate325inter8));
  nand2 gate1296(.a(gate325inter8), .b(gate325inter7), .O(gate325inter9));
  nand2 gate1297(.a(s_59), .b(gate325inter3), .O(gate325inter10));
  nor2  gate1298(.a(gate325inter10), .b(gate325inter9), .O(gate325inter11));
  nor2  gate1299(.a(gate325inter11), .b(gate325inter6), .O(gate325inter12));
  nand2 gate1300(.a(gate325inter12), .b(gate325inter1), .O(N1327));

  xor2  gate1217(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate1218(.a(gate326inter0), .b(s_48), .O(gate326inter1));
  and2  gate1219(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate1220(.a(s_48), .O(gate326inter3));
  inv1  gate1221(.a(s_49), .O(gate326inter4));
  nand2 gate1222(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate1223(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate1224(.a(N733), .O(gate326inter7));
  inv1  gate1225(.a(N1241), .O(gate326inter8));
  nand2 gate1226(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate1227(.a(s_49), .b(gate326inter3), .O(gate326inter10));
  nor2  gate1228(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate1229(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate1230(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );

  xor2  gate2477(.a(N894), .b(N1249), .O(gate329inter0));
  nand2 gate2478(.a(gate329inter0), .b(s_228), .O(gate329inter1));
  and2  gate2479(.a(N894), .b(N1249), .O(gate329inter2));
  inv1  gate2480(.a(s_228), .O(gate329inter3));
  inv1  gate2481(.a(s_229), .O(gate329inter4));
  nand2 gate2482(.a(gate329inter4), .b(gate329inter3), .O(gate329inter5));
  nor2  gate2483(.a(gate329inter5), .b(gate329inter2), .O(gate329inter6));
  inv1  gate2484(.a(N1249), .O(gate329inter7));
  inv1  gate2485(.a(N894), .O(gate329inter8));
  nand2 gate2486(.a(gate329inter8), .b(gate329inter7), .O(gate329inter9));
  nand2 gate2487(.a(s_229), .b(gate329inter3), .O(gate329inter10));
  nor2  gate2488(.a(gate329inter10), .b(gate329inter9), .O(gate329inter11));
  nor2  gate2489(.a(gate329inter11), .b(gate329inter6), .O(gate329inter12));
  nand2 gate2490(.a(gate329inter12), .b(gate329inter1), .O(N1345));
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );

  xor2  gate2967(.a(N1206), .b(N1309), .O(gate335inter0));
  nand2 gate2968(.a(gate335inter0), .b(s_298), .O(gate335inter1));
  and2  gate2969(.a(N1206), .b(N1309), .O(gate335inter2));
  inv1  gate2970(.a(s_298), .O(gate335inter3));
  inv1  gate2971(.a(s_299), .O(gate335inter4));
  nand2 gate2972(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate2973(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate2974(.a(N1309), .O(gate335inter7));
  inv1  gate2975(.a(N1206), .O(gate335inter8));
  nand2 gate2976(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate2977(.a(s_299), .b(gate335inter3), .O(gate335inter10));
  nor2  gate2978(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate2979(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate2980(.a(gate335inter12), .b(gate335inter1), .O(N1352));
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );

  xor2  gate2001(.a(N1216), .b(N1314), .O(gate340inter0));
  nand2 gate2002(.a(gate340inter0), .b(s_160), .O(gate340inter1));
  and2  gate2003(.a(N1216), .b(N1314), .O(gate340inter2));
  inv1  gate2004(.a(s_160), .O(gate340inter3));
  inv1  gate2005(.a(s_161), .O(gate340inter4));
  nand2 gate2006(.a(gate340inter4), .b(gate340inter3), .O(gate340inter5));
  nor2  gate2007(.a(gate340inter5), .b(gate340inter2), .O(gate340inter6));
  inv1  gate2008(.a(N1314), .O(gate340inter7));
  inv1  gate2009(.a(N1216), .O(gate340inter8));
  nand2 gate2010(.a(gate340inter8), .b(gate340inter7), .O(gate340inter9));
  nand2 gate2011(.a(s_161), .b(gate340inter3), .O(gate340inter10));
  nor2  gate2012(.a(gate340inter10), .b(gate340inter9), .O(gate340inter11));
  nor2  gate2013(.a(gate340inter11), .b(gate340inter6), .O(gate340inter12));
  nand2 gate2014(.a(gate340inter12), .b(gate340inter1), .O(N1367));
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );

  xor2  gate1987(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate1988(.a(gate342inter0), .b(s_158), .O(gate342inter1));
  and2  gate1989(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate1990(.a(s_158), .O(gate342inter3));
  inv1  gate1991(.a(s_159), .O(gate342inter4));
  nand2 gate1992(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate1993(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate1994(.a(N1316), .O(gate342inter7));
  inv1  gate1995(.a(N1224), .O(gate342inter8));
  nand2 gate1996(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate1997(.a(s_159), .b(gate342inter3), .O(gate342inter10));
  nor2  gate1998(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate1999(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate2000(.a(gate342inter12), .b(gate342inter1), .O(N1373));
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );

  xor2  gate3037(.a(N1229), .b(N1318), .O(gate344inter0));
  nand2 gate3038(.a(gate344inter0), .b(s_308), .O(gate344inter1));
  and2  gate3039(.a(N1229), .b(N1318), .O(gate344inter2));
  inv1  gate3040(.a(s_308), .O(gate344inter3));
  inv1  gate3041(.a(s_309), .O(gate344inter4));
  nand2 gate3042(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate3043(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate3044(.a(N1318), .O(gate344inter7));
  inv1  gate3045(.a(N1229), .O(gate344inter8));
  nand2 gate3046(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate3047(.a(s_309), .b(gate344inter3), .O(gate344inter10));
  nor2  gate3048(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate3049(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate3050(.a(gate344inter12), .b(gate344inter1), .O(N1379));
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate1441(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate1442(.a(gate347inter0), .b(s_80), .O(gate347inter1));
  and2  gate1443(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate1444(.a(s_80), .O(gate347inter3));
  inv1  gate1445(.a(s_81), .O(gate347inter4));
  nand2 gate1446(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate1447(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate1448(.a(N1232), .O(gate347inter7));
  inv1  gate1449(.a(N990), .O(gate347inter8));
  nand2 gate1450(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate1451(.a(s_81), .b(gate347inter3), .O(gate347inter10));
  nor2  gate1452(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate1453(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate1454(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );

  xor2  gate1875(.a(N1239), .b(N1327), .O(gate350inter0));
  nand2 gate1876(.a(gate350inter0), .b(s_142), .O(gate350inter1));
  and2  gate1877(.a(N1239), .b(N1327), .O(gate350inter2));
  inv1  gate1878(.a(s_142), .O(gate350inter3));
  inv1  gate1879(.a(s_143), .O(gate350inter4));
  nand2 gate1880(.a(gate350inter4), .b(gate350inter3), .O(gate350inter5));
  nor2  gate1881(.a(gate350inter5), .b(gate350inter2), .O(gate350inter6));
  inv1  gate1882(.a(N1327), .O(gate350inter7));
  inv1  gate1883(.a(N1239), .O(gate350inter8));
  nand2 gate1884(.a(gate350inter8), .b(gate350inter7), .O(gate350inter9));
  nand2 gate1885(.a(s_143), .b(gate350inter3), .O(gate350inter10));
  nor2  gate1886(.a(gate350inter10), .b(gate350inter9), .O(gate350inter11));
  nor2  gate1887(.a(gate350inter11), .b(gate350inter6), .O(gate350inter12));
  nand2 gate1888(.a(gate350inter12), .b(gate350inter1), .O(N1390));

  xor2  gate1035(.a(N1242), .b(N1328), .O(gate351inter0));
  nand2 gate1036(.a(gate351inter0), .b(s_22), .O(gate351inter1));
  and2  gate1037(.a(N1242), .b(N1328), .O(gate351inter2));
  inv1  gate1038(.a(s_22), .O(gate351inter3));
  inv1  gate1039(.a(s_23), .O(gate351inter4));
  nand2 gate1040(.a(gate351inter4), .b(gate351inter3), .O(gate351inter5));
  nor2  gate1041(.a(gate351inter5), .b(gate351inter2), .O(gate351inter6));
  inv1  gate1042(.a(N1328), .O(gate351inter7));
  inv1  gate1043(.a(N1242), .O(gate351inter8));
  nand2 gate1044(.a(gate351inter8), .b(gate351inter7), .O(gate351inter9));
  nand2 gate1045(.a(s_23), .b(gate351inter3), .O(gate351inter10));
  nor2  gate1046(.a(gate351inter10), .b(gate351inter9), .O(gate351inter11));
  nor2  gate1047(.a(gate351inter11), .b(gate351inter6), .O(gate351inter12));
  nand2 gate1048(.a(gate351inter12), .b(gate351inter1), .O(N1393));
inv1 gate352( .a(N1243), .O(N1396) );

  xor2  gate3233(.a(N1004), .b(N1243), .O(gate353inter0));
  nand2 gate3234(.a(gate353inter0), .b(s_336), .O(gate353inter1));
  and2  gate3235(.a(N1004), .b(N1243), .O(gate353inter2));
  inv1  gate3236(.a(s_336), .O(gate353inter3));
  inv1  gate3237(.a(s_337), .O(gate353inter4));
  nand2 gate3238(.a(gate353inter4), .b(gate353inter3), .O(gate353inter5));
  nor2  gate3239(.a(gate353inter5), .b(gate353inter2), .O(gate353inter6));
  inv1  gate3240(.a(N1243), .O(gate353inter7));
  inv1  gate3241(.a(N1004), .O(gate353inter8));
  nand2 gate3242(.a(gate353inter8), .b(gate353inter7), .O(gate353inter9));
  nand2 gate3243(.a(s_337), .b(gate353inter3), .O(gate353inter10));
  nor2  gate3244(.a(gate353inter10), .b(gate353inter9), .O(gate353inter11));
  nor2  gate3245(.a(gate353inter11), .b(gate353inter6), .O(gate353inter12));
  nand2 gate3246(.a(gate353inter12), .b(gate353inter1), .O(N1397));
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );

  xor2  gate3387(.a(N1346), .b(N649), .O(gate357inter0));
  nand2 gate3388(.a(gate357inter0), .b(s_358), .O(gate357inter1));
  and2  gate3389(.a(N1346), .b(N649), .O(gate357inter2));
  inv1  gate3390(.a(s_358), .O(gate357inter3));
  inv1  gate3391(.a(s_359), .O(gate357inter4));
  nand2 gate3392(.a(gate357inter4), .b(gate357inter3), .O(gate357inter5));
  nor2  gate3393(.a(gate357inter5), .b(gate357inter2), .O(gate357inter6));
  inv1  gate3394(.a(N649), .O(gate357inter7));
  inv1  gate3395(.a(N1346), .O(gate357inter8));
  nand2 gate3396(.a(gate357inter8), .b(gate357inter7), .O(gate357inter9));
  nand2 gate3397(.a(s_359), .b(gate357inter3), .O(gate357inter10));
  nor2  gate3398(.a(gate357inter10), .b(gate357inter9), .O(gate357inter11));
  nor2  gate3399(.a(gate357inter11), .b(gate357inter6), .O(gate357inter12));
  nand2 gate3400(.a(gate357inter12), .b(gate357inter1), .O(N1412));
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );

  xor2  gate2043(.a(N1386), .b(N634), .O(gate361inter0));
  nand2 gate2044(.a(gate361inter0), .b(s_166), .O(gate361inter1));
  and2  gate2045(.a(N1386), .b(N634), .O(gate361inter2));
  inv1  gate2046(.a(s_166), .O(gate361inter3));
  inv1  gate2047(.a(s_167), .O(gate361inter4));
  nand2 gate2048(.a(gate361inter4), .b(gate361inter3), .O(gate361inter5));
  nor2  gate2049(.a(gate361inter5), .b(gate361inter2), .O(gate361inter6));
  inv1  gate2050(.a(N634), .O(gate361inter7));
  inv1  gate2051(.a(N1386), .O(gate361inter8));
  nand2 gate2052(.a(gate361inter8), .b(gate361inter7), .O(gate361inter9));
  nand2 gate2053(.a(s_167), .b(gate361inter3), .O(gate361inter10));
  nor2  gate2054(.a(gate361inter10), .b(gate361inter9), .O(gate361inter11));
  nor2  gate2055(.a(gate361inter11), .b(gate361inter6), .O(gate361inter12));
  nand2 gate2056(.a(gate361inter12), .b(gate361inter1), .O(N1433));

  xor2  gate2113(.a(N1388), .b(N637), .O(gate362inter0));
  nand2 gate2114(.a(gate362inter0), .b(s_176), .O(gate362inter1));
  and2  gate2115(.a(N1388), .b(N637), .O(gate362inter2));
  inv1  gate2116(.a(s_176), .O(gate362inter3));
  inv1  gate2117(.a(s_177), .O(gate362inter4));
  nand2 gate2118(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate2119(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate2120(.a(N637), .O(gate362inter7));
  inv1  gate2121(.a(N1388), .O(gate362inter8));
  nand2 gate2122(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate2123(.a(s_177), .b(gate362inter3), .O(gate362inter10));
  nor2  gate2124(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate2125(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate2126(.a(gate362inter12), .b(gate362inter1), .O(N1434));
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );

  xor2  gate3317(.a(N1398), .b(N646), .O(gate364inter0));
  nand2 gate3318(.a(gate364inter0), .b(s_348), .O(gate364inter1));
  and2  gate3319(.a(N1398), .b(N646), .O(gate364inter2));
  inv1  gate3320(.a(s_348), .O(gate364inter3));
  inv1  gate3321(.a(s_349), .O(gate364inter4));
  nand2 gate3322(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate3323(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate3324(.a(N646), .O(gate364inter7));
  inv1  gate3325(.a(N1398), .O(gate364inter8));
  nand2 gate3326(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate3327(.a(s_349), .b(gate364inter3), .O(gate364inter10));
  nor2  gate3328(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate3329(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate3330(.a(gate364inter12), .b(gate364inter1), .O(N1439));
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );

  xor2  gate2505(.a(N1149), .b(N1352), .O(gate368inter0));
  nand2 gate2506(.a(gate368inter0), .b(s_232), .O(gate368inter1));
  and2  gate2507(.a(N1149), .b(N1352), .O(gate368inter2));
  inv1  gate2508(.a(s_232), .O(gate368inter3));
  inv1  gate2509(.a(s_233), .O(gate368inter4));
  nand2 gate2510(.a(gate368inter4), .b(gate368inter3), .O(gate368inter5));
  nor2  gate2511(.a(gate368inter5), .b(gate368inter2), .O(gate368inter6));
  inv1  gate2512(.a(N1352), .O(gate368inter7));
  inv1  gate2513(.a(N1149), .O(gate368inter8));
  nand2 gate2514(.a(gate368inter8), .b(gate368inter7), .O(gate368inter9));
  nand2 gate2515(.a(s_233), .b(gate368inter3), .O(gate368inter10));
  nor2  gate2516(.a(gate368inter10), .b(gate368inter9), .O(gate368inter11));
  nor2  gate2517(.a(gate368inter11), .b(gate368inter6), .O(gate368inter12));
  nand2 gate2518(.a(gate368inter12), .b(gate368inter1), .O(N1445));
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );

  xor2  gate1623(.a(N1153), .b(N1367), .O(gate374inter0));
  nand2 gate1624(.a(gate374inter0), .b(s_106), .O(gate374inter1));
  and2  gate1625(.a(N1153), .b(N1367), .O(gate374inter2));
  inv1  gate1626(.a(s_106), .O(gate374inter3));
  inv1  gate1627(.a(s_107), .O(gate374inter4));
  nand2 gate1628(.a(gate374inter4), .b(gate374inter3), .O(gate374inter5));
  nor2  gate1629(.a(gate374inter5), .b(gate374inter2), .O(gate374inter6));
  inv1  gate1630(.a(N1367), .O(gate374inter7));
  inv1  gate1631(.a(N1153), .O(gate374inter8));
  nand2 gate1632(.a(gate374inter8), .b(gate374inter7), .O(gate374inter9));
  nand2 gate1633(.a(s_107), .b(gate374inter3), .O(gate374inter10));
  nor2  gate1634(.a(gate374inter10), .b(gate374inter9), .O(gate374inter11));
  nor2  gate1635(.a(gate374inter11), .b(gate374inter6), .O(gate374inter12));
  nand2 gate1636(.a(gate374inter12), .b(gate374inter1), .O(N1453));
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate3191(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate3192(.a(gate376inter0), .b(s_330), .O(gate376inter1));
  and2  gate3193(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate3194(.a(s_330), .O(gate376inter3));
  inv1  gate3195(.a(s_331), .O(gate376inter4));
  nand2 gate3196(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate3197(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate3198(.a(N1364), .O(gate376inter7));
  inv1  gate3199(.a(N1154), .O(gate376inter8));
  nand2 gate3200(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate3201(.a(s_331), .b(gate376inter3), .O(gate376inter10));
  nor2  gate3202(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate3203(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate3204(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );

  xor2  gate3401(.a(N1156), .b(N1373), .O(gate378inter0));
  nand2 gate3402(.a(gate378inter0), .b(s_360), .O(gate378inter1));
  and2  gate3403(.a(N1156), .b(N1373), .O(gate378inter2));
  inv1  gate3404(.a(s_360), .O(gate378inter3));
  inv1  gate3405(.a(s_361), .O(gate378inter4));
  nand2 gate3406(.a(gate378inter4), .b(gate378inter3), .O(gate378inter5));
  nor2  gate3407(.a(gate378inter5), .b(gate378inter2), .O(gate378inter6));
  inv1  gate3408(.a(N1373), .O(gate378inter7));
  inv1  gate3409(.a(N1156), .O(gate378inter8));
  nand2 gate3410(.a(gate378inter8), .b(gate378inter7), .O(gate378inter9));
  nand2 gate3411(.a(s_361), .b(gate378inter3), .O(gate378inter10));
  nor2  gate3412(.a(gate378inter10), .b(gate378inter9), .O(gate378inter11));
  nor2  gate3413(.a(gate378inter11), .b(gate378inter6), .O(gate378inter12));
  nand2 gate3414(.a(gate378inter12), .b(gate378inter1), .O(N1457));
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate1553(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate1554(.a(gate383inter0), .b(s_96), .O(gate383inter1));
  and2  gate1555(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate1556(.a(s_96), .O(gate383inter3));
  inv1  gate1557(.a(s_97), .O(gate383inter4));
  nand2 gate1558(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate1559(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate1560(.a(N1393), .O(gate383inter7));
  inv1  gate1561(.a(N1161), .O(gate383inter8));
  nand2 gate1562(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate1563(.a(s_97), .b(gate383inter3), .O(gate383inter10));
  nor2  gate1564(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate1565(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate1566(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );

  xor2  gate1343(.a(N1222), .b(N1370), .O(gate387inter0));
  nand2 gate1344(.a(gate387inter0), .b(s_66), .O(gate387inter1));
  and2  gate1345(.a(N1222), .b(N1370), .O(gate387inter2));
  inv1  gate1346(.a(s_66), .O(gate387inter3));
  inv1  gate1347(.a(s_67), .O(gate387inter4));
  nand2 gate1348(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1349(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1350(.a(N1370), .O(gate387inter7));
  inv1  gate1351(.a(N1222), .O(gate387inter8));
  nand2 gate1352(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1353(.a(s_67), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1354(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1355(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1356(.a(gate387inter12), .b(gate387inter1), .O(N1469));
inv1 gate388( .a(N1376), .O(N1470) );

  xor2  gate1469(.a(N1227), .b(N1376), .O(gate389inter0));
  nand2 gate1470(.a(gate389inter0), .b(s_84), .O(gate389inter1));
  and2  gate1471(.a(N1227), .b(N1376), .O(gate389inter2));
  inv1  gate1472(.a(s_84), .O(gate389inter3));
  inv1  gate1473(.a(s_85), .O(gate389inter4));
  nand2 gate1474(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1475(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1476(.a(N1376), .O(gate389inter7));
  inv1  gate1477(.a(N1227), .O(gate389inter8));
  nand2 gate1478(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1479(.a(s_85), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1480(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1481(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1482(.a(gate389inter12), .b(gate389inter1), .O(N1471));

  xor2  gate3093(.a(N1433), .b(N1387), .O(gate390inter0));
  nand2 gate3094(.a(gate390inter0), .b(s_316), .O(gate390inter1));
  and2  gate3095(.a(N1433), .b(N1387), .O(gate390inter2));
  inv1  gate3096(.a(s_316), .O(gate390inter3));
  inv1  gate3097(.a(s_317), .O(gate390inter4));
  nand2 gate3098(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate3099(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate3100(.a(N1387), .O(gate390inter7));
  inv1  gate3101(.a(N1433), .O(gate390inter8));
  nand2 gate3102(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate3103(.a(s_317), .b(gate390inter3), .O(gate390inter10));
  nor2  gate3104(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate3105(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate3106(.a(gate390inter12), .b(gate390inter1), .O(N1472));
inv1 gate391( .a(N1390), .O(N1475) );

  xor2  gate1147(.a(N1240), .b(N1390), .O(gate392inter0));
  nand2 gate1148(.a(gate392inter0), .b(s_38), .O(gate392inter1));
  and2  gate1149(.a(N1240), .b(N1390), .O(gate392inter2));
  inv1  gate1150(.a(s_38), .O(gate392inter3));
  inv1  gate1151(.a(s_39), .O(gate392inter4));
  nand2 gate1152(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1153(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1154(.a(N1390), .O(gate392inter7));
  inv1  gate1155(.a(N1240), .O(gate392inter8));
  nand2 gate1156(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1157(.a(s_39), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1158(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1159(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1160(.a(gate392inter12), .b(gate392inter1), .O(N1476));

  xor2  gate2645(.a(N1434), .b(N1389), .O(gate393inter0));
  nand2 gate2646(.a(gate393inter0), .b(s_252), .O(gate393inter1));
  and2  gate2647(.a(N1434), .b(N1389), .O(gate393inter2));
  inv1  gate2648(.a(s_252), .O(gate393inter3));
  inv1  gate2649(.a(s_253), .O(gate393inter4));
  nand2 gate2650(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2651(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2652(.a(N1389), .O(gate393inter7));
  inv1  gate2653(.a(N1434), .O(gate393inter8));
  nand2 gate2654(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2655(.a(s_253), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2656(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2657(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2658(.a(gate393inter12), .b(gate393inter1), .O(N1478));
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );

  xor2  gate3345(.a(N1444), .b(N939), .O(gate396inter0));
  nand2 gate3346(.a(gate396inter0), .b(s_352), .O(gate396inter1));
  and2  gate3347(.a(N1444), .b(N939), .O(gate396inter2));
  inv1  gate3348(.a(s_352), .O(gate396inter3));
  inv1  gate3349(.a(s_353), .O(gate396inter4));
  nand2 gate3350(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate3351(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate3352(.a(N939), .O(gate396inter7));
  inv1  gate3353(.a(N1444), .O(gate396inter8));
  nand2 gate3354(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate3355(.a(s_353), .b(gate396inter3), .O(gate396inter10));
  nor2  gate3356(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate3357(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate3358(.a(gate396inter12), .b(gate396inter1), .O(N1487));
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );

  xor2  gate1805(.a(N1448), .b(N943), .O(gate398inter0));
  nand2 gate1806(.a(gate398inter0), .b(s_132), .O(gate398inter1));
  and2  gate1807(.a(N1448), .b(N943), .O(gate398inter2));
  inv1  gate1808(.a(s_132), .O(gate398inter3));
  inv1  gate1809(.a(s_133), .O(gate398inter4));
  nand2 gate1810(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1811(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1812(.a(N943), .O(gate398inter7));
  inv1  gate1813(.a(N1448), .O(gate398inter8));
  nand2 gate1814(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1815(.a(s_133), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1816(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1817(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1818(.a(gate398inter12), .b(gate398inter1), .O(N1489));
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );

  xor2  gate2715(.a(N1452), .b(N947), .O(gate401inter0));
  nand2 gate2716(.a(gate401inter0), .b(s_262), .O(gate401inter1));
  and2  gate2717(.a(N1452), .b(N947), .O(gate401inter2));
  inv1  gate2718(.a(s_262), .O(gate401inter3));
  inv1  gate2719(.a(s_263), .O(gate401inter4));
  nand2 gate2720(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2721(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2722(.a(N947), .O(gate401inter7));
  inv1  gate2723(.a(N1452), .O(gate401inter8));
  nand2 gate2724(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2725(.a(s_263), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2726(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2727(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2728(.a(gate401inter12), .b(gate401inter1), .O(N1492));
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );

  xor2  gate1959(.a(N1456), .b(N951), .O(gate403inter0));
  nand2 gate1960(.a(gate403inter0), .b(s_154), .O(gate403inter1));
  and2  gate1961(.a(N1456), .b(N951), .O(gate403inter2));
  inv1  gate1962(.a(s_154), .O(gate403inter3));
  inv1  gate1963(.a(s_155), .O(gate403inter4));
  nand2 gate1964(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1965(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1966(.a(N951), .O(gate403inter7));
  inv1  gate1967(.a(N1456), .O(gate403inter8));
  nand2 gate1968(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1969(.a(s_155), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1970(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1971(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1972(.a(gate403inter12), .b(gate403inter1), .O(N1494));
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );

  xor2  gate1161(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate1162(.a(gate406inter0), .b(s_40), .O(gate406inter1));
  and2  gate1163(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate1164(.a(s_40), .O(gate406inter3));
  inv1  gate1165(.a(s_41), .O(gate406inter4));
  nand2 gate1166(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1167(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1168(.a(N998), .O(gate406inter7));
  inv1  gate1169(.a(N1463), .O(gate406inter8));
  nand2 gate1170(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1171(.a(s_41), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1172(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1173(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1174(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );

  xor2  gate3373(.a(N1487), .b(N1443), .O(gate412inter0));
  nand2 gate3374(.a(gate412inter0), .b(s_356), .O(gate412inter1));
  and2  gate3375(.a(N1487), .b(N1443), .O(gate412inter2));
  inv1  gate3376(.a(s_356), .O(gate412inter3));
  inv1  gate3377(.a(s_357), .O(gate412inter4));
  nand2 gate3378(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate3379(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate3380(.a(N1443), .O(gate412inter7));
  inv1  gate3381(.a(N1487), .O(gate412inter8));
  nand2 gate3382(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate3383(.a(s_357), .b(gate412inter3), .O(gate412inter10));
  nor2  gate3384(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate3385(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate3386(.a(gate412inter12), .b(gate412inter1), .O(N1513));

  xor2  gate2491(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate2492(.a(gate413inter0), .b(s_230), .O(gate413inter1));
  and2  gate2493(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate2494(.a(s_230), .O(gate413inter3));
  inv1  gate2495(.a(s_231), .O(gate413inter4));
  nand2 gate2496(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2497(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2498(.a(N1445), .O(gate413inter7));
  inv1  gate2499(.a(N1488), .O(gate413inter8));
  nand2 gate2500(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2501(.a(s_231), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2502(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2503(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2504(.a(gate413inter12), .b(gate413inter1), .O(N1514));
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );

  xor2  gate1119(.a(N1492), .b(N1451), .O(gate415inter0));
  nand2 gate1120(.a(gate415inter0), .b(s_34), .O(gate415inter1));
  and2  gate1121(.a(N1492), .b(N1451), .O(gate415inter2));
  inv1  gate1122(.a(s_34), .O(gate415inter3));
  inv1  gate1123(.a(s_35), .O(gate415inter4));
  nand2 gate1124(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1125(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1126(.a(N1451), .O(gate415inter7));
  inv1  gate1127(.a(N1492), .O(gate415inter8));
  nand2 gate1128(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1129(.a(s_35), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1130(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1131(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1132(.a(gate415inter12), .b(gate415inter1), .O(N1520));

  xor2  gate2239(.a(N1493), .b(N1453), .O(gate416inter0));
  nand2 gate2240(.a(gate416inter0), .b(s_194), .O(gate416inter1));
  and2  gate2241(.a(N1493), .b(N1453), .O(gate416inter2));
  inv1  gate2242(.a(s_194), .O(gate416inter3));
  inv1  gate2243(.a(s_195), .O(gate416inter4));
  nand2 gate2244(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2245(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2246(.a(N1453), .O(gate416inter7));
  inv1  gate2247(.a(N1493), .O(gate416inter8));
  nand2 gate2248(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2249(.a(s_195), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2250(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2251(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2252(.a(gate416inter12), .b(gate416inter1), .O(N1521));

  xor2  gate2533(.a(N1494), .b(N1455), .O(gate417inter0));
  nand2 gate2534(.a(gate417inter0), .b(s_236), .O(gate417inter1));
  and2  gate2535(.a(N1494), .b(N1455), .O(gate417inter2));
  inv1  gate2536(.a(s_236), .O(gate417inter3));
  inv1  gate2537(.a(s_237), .O(gate417inter4));
  nand2 gate2538(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2539(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2540(.a(N1455), .O(gate417inter7));
  inv1  gate2541(.a(N1494), .O(gate417inter8));
  nand2 gate2542(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2543(.a(s_237), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2544(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2545(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2546(.a(gate417inter12), .b(gate417inter1), .O(N1522));
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate1133(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate1134(.a(gate421inter0), .b(s_36), .O(gate421inter1));
  and2  gate1135(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate1136(.a(s_36), .O(gate421inter3));
  inv1  gate1137(.a(s_37), .O(gate421inter4));
  nand2 gate1138(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1139(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1140(.a(N1462), .O(gate421inter7));
  inv1  gate1141(.a(N1498), .O(gate421inter8));
  nand2 gate1142(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1143(.a(s_37), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1144(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1145(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1146(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );

  xor2  gate1945(.a(N1532), .b(N1481), .O(gate433inter0));
  nand2 gate1946(.a(gate433inter0), .b(s_152), .O(gate433inter1));
  and2  gate1947(.a(N1532), .b(N1481), .O(gate433inter2));
  inv1  gate1948(.a(s_152), .O(gate433inter3));
  inv1  gate1949(.a(s_153), .O(gate433inter4));
  nand2 gate1950(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1951(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1952(.a(N1481), .O(gate433inter7));
  inv1  gate1953(.a(N1532), .O(gate433inter8));
  nand2 gate1954(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1955(.a(s_153), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1956(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1957(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1958(.a(gate433inter12), .b(gate433inter1), .O(N1568));
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );

  xor2  gate2911(.a(N1568), .b(N1567), .O(gate442inter0));
  nand2 gate2912(.a(gate442inter0), .b(s_290), .O(gate442inter1));
  and2  gate2913(.a(N1568), .b(N1567), .O(gate442inter2));
  inv1  gate2914(.a(s_290), .O(gate442inter3));
  inv1  gate2915(.a(s_291), .O(gate442inter4));
  nand2 gate2916(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2917(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2918(.a(N1567), .O(gate442inter7));
  inv1  gate2919(.a(N1568), .O(gate442inter8));
  nand2 gate2920(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2921(.a(s_291), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2922(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2923(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2924(.a(gate442inter12), .b(gate442inter1), .O(N1596));
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );

  xor2  gate1021(.a(N893), .b(N1596), .O(gate462inter0));
  nand2 gate1022(.a(gate462inter0), .b(s_20), .O(gate462inter1));
  and2  gate1023(.a(N893), .b(N1596), .O(gate462inter2));
  inv1  gate1024(.a(s_20), .O(gate462inter3));
  inv1  gate1025(.a(s_21), .O(gate462inter4));
  nand2 gate1026(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1027(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1028(.a(N1596), .O(gate462inter7));
  inv1  gate1029(.a(N893), .O(gate462inter8));
  nand2 gate1030(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1031(.a(s_21), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1032(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1033(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1034(.a(gate462inter12), .b(gate462inter1), .O(N1671));
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );

  xor2  gate2029(.a(N1636), .b(N1594), .O(gate472inter0));
  nand2 gate2030(.a(gate472inter0), .b(s_164), .O(gate472inter1));
  and2  gate2031(.a(N1636), .b(N1594), .O(gate472inter2));
  inv1  gate2032(.a(s_164), .O(gate472inter3));
  inv1  gate2033(.a(s_165), .O(gate472inter4));
  nand2 gate2034(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2035(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2036(.a(N1594), .O(gate472inter7));
  inv1  gate2037(.a(N1636), .O(gate472inter8));
  nand2 gate2038(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2039(.a(s_165), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2040(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2041(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2042(.a(gate472inter12), .b(gate472inter1), .O(N1685));

  xor2  gate2337(.a(N1639), .b(N1510), .O(gate473inter0));
  nand2 gate2338(.a(gate473inter0), .b(s_208), .O(gate473inter1));
  and2  gate2339(.a(N1639), .b(N1510), .O(gate473inter2));
  inv1  gate2340(.a(s_208), .O(gate473inter3));
  inv1  gate2341(.a(s_209), .O(gate473inter4));
  nand2 gate2342(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2343(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2344(.a(N1510), .O(gate473inter7));
  inv1  gate2345(.a(N1639), .O(gate473inter8));
  nand2 gate2346(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2347(.a(s_209), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2348(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2349(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2350(.a(gate473inter12), .b(gate473inter1), .O(N1688));
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );

  xor2  gate2407(.a(N1672), .b(N643), .O(gate476inter0));
  nand2 gate2408(.a(gate476inter0), .b(s_218), .O(gate476inter1));
  and2  gate2409(.a(N1672), .b(N643), .O(gate476inter2));
  inv1  gate2410(.a(s_218), .O(gate476inter3));
  inv1  gate2411(.a(s_219), .O(gate476inter4));
  nand2 gate2412(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2413(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2414(.a(N643), .O(gate476inter7));
  inv1  gate2415(.a(N1672), .O(gate476inter8));
  nand2 gate2416(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2417(.a(s_219), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2418(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2419(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2420(.a(gate476inter12), .b(gate476inter1), .O(N1706));
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );

  xor2  gate1777(.a(N1677), .b(N1651), .O(gate480inter0));
  nand2 gate1778(.a(gate480inter0), .b(s_128), .O(gate480inter1));
  and2  gate1779(.a(N1677), .b(N1651), .O(gate480inter2));
  inv1  gate1780(.a(s_128), .O(gate480inter3));
  inv1  gate1781(.a(s_129), .O(gate480inter4));
  nand2 gate1782(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1783(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1784(.a(N1651), .O(gate480inter7));
  inv1  gate1785(.a(N1677), .O(gate480inter8));
  nand2 gate1786(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1787(.a(s_129), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1788(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1789(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1790(.a(gate480inter12), .b(gate480inter1), .O(N1710));
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );

  xor2  gate2085(.a(N1688), .b(N1638), .O(gate488inter0));
  nand2 gate2086(.a(gate488inter0), .b(s_172), .O(gate488inter1));
  and2  gate2087(.a(N1688), .b(N1638), .O(gate488inter2));
  inv1  gate2088(.a(s_172), .O(gate488inter3));
  inv1  gate2089(.a(s_173), .O(gate488inter4));
  nand2 gate2090(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2091(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2092(.a(N1638), .O(gate488inter7));
  inv1  gate2093(.a(N1688), .O(gate488inter8));
  nand2 gate2094(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2095(.a(s_173), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2096(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2097(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2098(.a(gate488inter12), .b(gate488inter1), .O(N1723));
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );

  xor2  gate2995(.a(N1528), .b(N1685), .O(gate494inter0));
  nand2 gate2996(.a(gate494inter0), .b(s_302), .O(gate494inter1));
  and2  gate2997(.a(N1528), .b(N1685), .O(gate494inter2));
  inv1  gate2998(.a(s_302), .O(gate494inter3));
  inv1  gate2999(.a(s_303), .O(gate494inter4));
  nand2 gate3000(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate3001(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate3002(.a(N1685), .O(gate494inter7));
  inv1  gate3003(.a(N1528), .O(gate494inter8));
  nand2 gate3004(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate3005(.a(s_303), .b(gate494inter3), .O(gate494inter10));
  nor2  gate3006(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate3007(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate3008(.a(gate494inter12), .b(gate494inter1), .O(N1740));
inv1 gate495( .a(N1685), .O(N1741) );

  xor2  gate1567(.a(N1706), .b(N1671), .O(gate496inter0));
  nand2 gate1568(.a(gate496inter0), .b(s_98), .O(gate496inter1));
  and2  gate1569(.a(N1706), .b(N1671), .O(gate496inter2));
  inv1  gate1570(.a(s_98), .O(gate496inter3));
  inv1  gate1571(.a(s_99), .O(gate496inter4));
  nand2 gate1572(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1573(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1574(.a(N1671), .O(gate496inter7));
  inv1  gate1575(.a(N1706), .O(gate496inter8));
  nand2 gate1576(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1577(.a(s_99), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1578(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1579(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1580(.a(gate496inter12), .b(gate496inter1), .O(N1742));

  xor2  gate2897(.a(N1709), .b(N1600), .O(gate497inter0));
  nand2 gate2898(.a(gate497inter0), .b(s_288), .O(gate497inter1));
  and2  gate2899(.a(N1709), .b(N1600), .O(gate497inter2));
  inv1  gate2900(.a(s_288), .O(gate497inter3));
  inv1  gate2901(.a(s_289), .O(gate497inter4));
  nand2 gate2902(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2903(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2904(.a(N1600), .O(gate497inter7));
  inv1  gate2905(.a(N1709), .O(gate497inter8));
  nand2 gate2906(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2907(.a(s_289), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2908(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2909(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2910(.a(gate497inter12), .b(gate497inter1), .O(N1746));

  xor2  gate3079(.a(N1711), .b(N1603), .O(gate498inter0));
  nand2 gate3080(.a(gate498inter0), .b(s_314), .O(gate498inter1));
  and2  gate3081(.a(N1711), .b(N1603), .O(gate498inter2));
  inv1  gate3082(.a(s_314), .O(gate498inter3));
  inv1  gate3083(.a(s_315), .O(gate498inter4));
  nand2 gate3084(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate3085(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate3086(.a(N1603), .O(gate498inter7));
  inv1  gate3087(.a(N1711), .O(gate498inter8));
  nand2 gate3088(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate3089(.a(s_315), .b(gate498inter3), .O(gate498inter10));
  nor2  gate3090(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate3091(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate3092(.a(gate498inter12), .b(gate498inter1), .O(N1747));
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );

  xor2  gate1917(.a(N1713), .b(N1680), .O(gate500inter0));
  nand2 gate1918(.a(gate500inter0), .b(s_148), .O(gate500inter1));
  and2  gate1919(.a(N1713), .b(N1680), .O(gate500inter2));
  inv1  gate1920(.a(s_148), .O(gate500inter3));
  inv1  gate1921(.a(s_149), .O(gate500inter4));
  nand2 gate1922(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1923(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1924(.a(N1680), .O(gate500inter7));
  inv1  gate1925(.a(N1713), .O(gate500inter8));
  nand2 gate1926(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1927(.a(s_149), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1928(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1929(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1930(.a(gate500inter12), .b(gate500inter1), .O(N1751));

  xor2  gate881(.a(N1721), .b(N1537), .O(gate501inter0));
  nand2 gate882(.a(gate501inter0), .b(s_0), .O(gate501inter1));
  and2  gate883(.a(N1721), .b(N1537), .O(gate501inter2));
  inv1  gate884(.a(s_0), .O(gate501inter3));
  inv1  gate885(.a(s_1), .O(gate501inter4));
  nand2 gate886(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate887(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate888(.a(N1537), .O(gate501inter7));
  inv1  gate889(.a(N1721), .O(gate501inter8));
  nand2 gate890(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate891(.a(s_1), .b(gate501inter3), .O(gate501inter10));
  nor2  gate892(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate893(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate894(.a(gate501inter12), .b(gate501inter1), .O(N1759));
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate3331(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate3332(.a(gate503inter0), .b(s_350), .O(gate503inter1));
  and2  gate3333(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate3334(.a(s_350), .O(gate503inter3));
  inv1  gate3335(.a(s_351), .O(gate503inter4));
  nand2 gate3336(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate3337(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate3338(.a(N1697), .O(gate503inter7));
  inv1  gate3339(.a(N1727), .O(gate503inter8));
  nand2 gate3340(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate3341(.a(s_351), .b(gate503inter3), .O(gate503inter10));
  nor2  gate3342(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate3343(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate3344(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );

  xor2  gate2547(.a(N1730), .b(N1701), .O(gate505inter0));
  nand2 gate2548(.a(gate505inter0), .b(s_238), .O(gate505inter1));
  and2  gate2549(.a(N1730), .b(N1701), .O(gate505inter2));
  inv1  gate2550(.a(s_238), .O(gate505inter3));
  inv1  gate2551(.a(s_239), .O(gate505inter4));
  nand2 gate2552(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2553(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2554(.a(N1701), .O(gate505inter7));
  inv1  gate2555(.a(N1730), .O(gate505inter8));
  nand2 gate2556(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2557(.a(s_239), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2558(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2559(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2560(.a(gate505inter12), .b(gate505inter1), .O(N1764));
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );

  xor2  gate2617(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate2618(.a(gate508inter0), .b(s_248), .O(gate508inter1));
  and2  gate2619(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate2620(.a(s_248), .O(gate508inter3));
  inv1  gate2621(.a(s_249), .O(gate508inter4));
  nand2 gate2622(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2623(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2624(.a(N1723), .O(gate508inter7));
  inv1  gate2625(.a(N1413), .O(gate508inter8));
  nand2 gate2626(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2627(.a(s_249), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2628(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2629(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2630(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );

  xor2  gate1497(.a(N1746), .b(N1708), .O(gate510inter0));
  nand2 gate1498(.a(gate510inter0), .b(s_88), .O(gate510inter1));
  and2  gate1499(.a(N1746), .b(N1708), .O(gate510inter2));
  inv1  gate1500(.a(s_88), .O(gate510inter3));
  inv1  gate1501(.a(s_89), .O(gate510inter4));
  nand2 gate1502(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1503(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1504(.a(N1708), .O(gate510inter7));
  inv1  gate1505(.a(N1746), .O(gate510inter8));
  nand2 gate1506(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1507(.a(s_89), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1508(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1509(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1510(.a(gate510inter12), .b(gate510inter1), .O(N1774));
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1931(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1932(.a(gate513inter0), .b(s_150), .O(gate513inter1));
  and2  gate1933(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1934(.a(s_150), .O(gate513inter3));
  inv1  gate1935(.a(s_151), .O(gate513inter4));
  nand2 gate1936(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1937(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1938(.a(N1731), .O(gate513inter7));
  inv1  gate1939(.a(N1682), .O(gate513inter8));
  nand2 gate1940(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1941(.a(s_151), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1942(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1943(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1944(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );

  xor2  gate2701(.a(N1683), .b(N1734), .O(gate516inter0));
  nand2 gate2702(.a(gate516inter0), .b(s_260), .O(gate516inter1));
  and2  gate2703(.a(N1683), .b(N1734), .O(gate516inter2));
  inv1  gate2704(.a(s_260), .O(gate516inter3));
  inv1  gate2705(.a(s_261), .O(gate516inter4));
  nand2 gate2706(.a(gate516inter4), .b(gate516inter3), .O(gate516inter5));
  nor2  gate2707(.a(gate516inter5), .b(gate516inter2), .O(gate516inter6));
  inv1  gate2708(.a(N1734), .O(gate516inter7));
  inv1  gate2709(.a(N1683), .O(gate516inter8));
  nand2 gate2710(.a(gate516inter8), .b(gate516inter7), .O(gate516inter9));
  nand2 gate2711(.a(s_261), .b(gate516inter3), .O(gate516inter10));
  nor2  gate2712(.a(gate516inter10), .b(gate516inter9), .O(gate516inter11));
  nor2  gate2713(.a(gate516inter11), .b(gate516inter6), .O(gate516inter12));
  nand2 gate2714(.a(gate516inter12), .b(gate516inter1), .O(N1787));

  xor2  gate1301(.a(N1759), .b(N1720), .O(gate517inter0));
  nand2 gate1302(.a(gate517inter0), .b(s_60), .O(gate517inter1));
  and2  gate1303(.a(N1759), .b(N1720), .O(gate517inter2));
  inv1  gate1304(.a(s_60), .O(gate517inter3));
  inv1  gate1305(.a(s_61), .O(gate517inter4));
  nand2 gate1306(.a(gate517inter4), .b(gate517inter3), .O(gate517inter5));
  nor2  gate1307(.a(gate517inter5), .b(gate517inter2), .O(gate517inter6));
  inv1  gate1308(.a(N1720), .O(gate517inter7));
  inv1  gate1309(.a(N1759), .O(gate517inter8));
  nand2 gate1310(.a(gate517inter8), .b(gate517inter7), .O(gate517inter9));
  nand2 gate1311(.a(s_61), .b(gate517inter3), .O(gate517inter10));
  nor2  gate1312(.a(gate517inter10), .b(gate517inter9), .O(gate517inter11));
  nor2  gate1313(.a(gate517inter11), .b(gate517inter6), .O(gate517inter12));
  nand2 gate1314(.a(gate517inter12), .b(gate517inter1), .O(N1788));
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );

  xor2  gate2575(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate2576(.a(gate520inter0), .b(s_242), .O(gate520inter1));
  and2  gate2577(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate2578(.a(s_242), .O(gate520inter3));
  inv1  gate2579(.a(s_243), .O(gate520inter4));
  nand2 gate2580(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate2581(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate2582(.a(N1751), .O(gate520inter7));
  inv1  gate2583(.a(N1155), .O(gate520inter8));
  nand2 gate2584(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate2585(.a(s_243), .b(gate520inter3), .O(gate520inter10));
  nor2  gate2586(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate2587(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate2588(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate3121(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate3122(.a(gate522inter0), .b(s_320), .O(gate522inter1));
  and2  gate3123(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate3124(.a(s_320), .O(gate522inter3));
  inv1  gate3125(.a(s_321), .O(gate522inter4));
  nand2 gate3126(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate3127(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate3128(.a(N1740), .O(gate522inter7));
  inv1  gate3129(.a(N1769), .O(gate522inter8));
  nand2 gate3130(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate3131(.a(s_321), .b(gate522inter3), .O(gate522inter10));
  nor2  gate3132(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate3133(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate3134(.a(gate522inter12), .b(gate522inter1), .O(N1798));
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );

  xor2  gate2925(.a(N1218), .b(N1748), .O(gate526inter0));
  nand2 gate2926(.a(gate526inter0), .b(s_292), .O(gate526inter1));
  and2  gate2927(.a(N1218), .b(N1748), .O(gate526inter2));
  inv1  gate2928(.a(s_292), .O(gate526inter3));
  inv1  gate2929(.a(s_293), .O(gate526inter4));
  nand2 gate2930(.a(gate526inter4), .b(gate526inter3), .O(gate526inter5));
  nor2  gate2931(.a(gate526inter5), .b(gate526inter2), .O(gate526inter6));
  inv1  gate2932(.a(N1748), .O(gate526inter7));
  inv1  gate2933(.a(N1218), .O(gate526inter8));
  nand2 gate2934(.a(gate526inter8), .b(gate526inter7), .O(gate526inter9));
  nand2 gate2935(.a(s_293), .b(gate526inter3), .O(gate526inter10));
  nor2  gate2936(.a(gate526inter10), .b(gate526inter9), .O(gate526inter11));
  nor2  gate2937(.a(gate526inter11), .b(gate526inter6), .O(gate526inter12));
  nand2 gate2938(.a(gate526inter12), .b(gate526inter1), .O(N1808));
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );

  xor2  gate2855(.a(N1786), .b(N1615), .O(gate528inter0));
  nand2 gate2856(.a(gate528inter0), .b(s_282), .O(gate528inter1));
  and2  gate2857(.a(N1786), .b(N1615), .O(gate528inter2));
  inv1  gate2858(.a(s_282), .O(gate528inter3));
  inv1  gate2859(.a(s_283), .O(gate528inter4));
  nand2 gate2860(.a(gate528inter4), .b(gate528inter3), .O(gate528inter5));
  nor2  gate2861(.a(gate528inter5), .b(gate528inter2), .O(gate528inter6));
  inv1  gate2862(.a(N1615), .O(gate528inter7));
  inv1  gate2863(.a(N1786), .O(gate528inter8));
  nand2 gate2864(.a(gate528inter8), .b(gate528inter7), .O(gate528inter9));
  nand2 gate2865(.a(s_283), .b(gate528inter3), .O(gate528inter10));
  nor2  gate2866(.a(gate528inter10), .b(gate528inter9), .O(gate528inter11));
  nor2  gate2867(.a(gate528inter11), .b(gate528inter6), .O(gate528inter12));
  nand2 gate2868(.a(gate528inter12), .b(gate528inter1), .O(N1810));

  xor2  gate3135(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate3136(.a(gate529inter0), .b(s_322), .O(gate529inter1));
  and2  gate3137(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate3138(.a(s_322), .O(gate529inter3));
  inv1  gate3139(.a(s_323), .O(gate529inter4));
  nand2 gate3140(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate3141(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate3142(.a(N1791), .O(gate529inter7));
  inv1  gate3143(.a(N1762), .O(gate529inter8));
  nand2 gate3144(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate3145(.a(s_323), .b(gate529inter3), .O(gate529inter10));
  nor2  gate3146(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate3147(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate3148(.a(gate529inter12), .b(gate529inter1), .O(N1812));
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate1847(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate1848(.a(gate532inter0), .b(s_138), .O(gate532inter1));
  and2  gate1849(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate1850(.a(s_138), .O(gate532inter3));
  inv1  gate1851(.a(s_139), .O(gate532inter4));
  nand2 gate1852(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate1853(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate1854(.a(N1777), .O(gate532inter7));
  inv1  gate1855(.a(N1490), .O(gate532inter8));
  nand2 gate1856(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate1857(.a(s_139), .b(gate532inter3), .O(gate532inter10));
  nor2  gate1858(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate1859(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate1860(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );

  xor2  gate2687(.a(N1491), .b(N1774), .O(gate534inter0));
  nand2 gate2688(.a(gate534inter0), .b(s_258), .O(gate534inter1));
  and2  gate2689(.a(N1491), .b(N1774), .O(gate534inter2));
  inv1  gate2690(.a(s_258), .O(gate534inter3));
  inv1  gate2691(.a(s_259), .O(gate534inter4));
  nand2 gate2692(.a(gate534inter4), .b(gate534inter3), .O(gate534inter5));
  nor2  gate2693(.a(gate534inter5), .b(gate534inter2), .O(gate534inter6));
  inv1  gate2694(.a(N1774), .O(gate534inter7));
  inv1  gate2695(.a(N1491), .O(gate534inter8));
  nand2 gate2696(.a(gate534inter8), .b(gate534inter7), .O(gate534inter9));
  nand2 gate2697(.a(s_259), .b(gate534inter3), .O(gate534inter10));
  nor2  gate2698(.a(gate534inter10), .b(gate534inter9), .O(gate534inter11));
  nor2  gate2699(.a(gate534inter11), .b(gate534inter6), .O(gate534inter12));
  nand2 gate2700(.a(gate534inter12), .b(gate534inter1), .O(N1823));
inv1 gate535( .a(N1774), .O(N1824) );

  xor2  gate2869(.a(N1796), .b(N962), .O(gate536inter0));
  nand2 gate2870(.a(gate536inter0), .b(s_284), .O(gate536inter1));
  and2  gate2871(.a(N1796), .b(N962), .O(gate536inter2));
  inv1  gate2872(.a(s_284), .O(gate536inter3));
  inv1  gate2873(.a(s_285), .O(gate536inter4));
  nand2 gate2874(.a(gate536inter4), .b(gate536inter3), .O(gate536inter5));
  nor2  gate2875(.a(gate536inter5), .b(gate536inter2), .O(gate536inter6));
  inv1  gate2876(.a(N962), .O(gate536inter7));
  inv1  gate2877(.a(N1796), .O(gate536inter8));
  nand2 gate2878(.a(gate536inter8), .b(gate536inter7), .O(gate536inter9));
  nand2 gate2879(.a(s_285), .b(gate536inter3), .O(gate536inter10));
  nor2  gate2880(.a(gate536inter10), .b(gate536inter9), .O(gate536inter11));
  nor2  gate2881(.a(gate536inter11), .b(gate536inter6), .O(gate536inter12));
  nand2 gate2882(.a(gate536inter12), .b(gate536inter1), .O(N1825));
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );

  xor2  gate1007(.a(N1784), .b(N1809), .O(gate541inter0));
  nand2 gate1008(.a(gate541inter0), .b(s_18), .O(gate541inter1));
  and2  gate1009(.a(N1784), .b(N1809), .O(gate541inter2));
  inv1  gate1010(.a(s_18), .O(gate541inter3));
  inv1  gate1011(.a(s_19), .O(gate541inter4));
  nand2 gate1012(.a(gate541inter4), .b(gate541inter3), .O(gate541inter5));
  nor2  gate1013(.a(gate541inter5), .b(gate541inter2), .O(gate541inter6));
  inv1  gate1014(.a(N1809), .O(gate541inter7));
  inv1  gate1015(.a(N1784), .O(gate541inter8));
  nand2 gate1016(.a(gate541inter8), .b(gate541inter7), .O(gate541inter9));
  nand2 gate1017(.a(s_19), .b(gate541inter3), .O(gate541inter10));
  nor2  gate1018(.a(gate541inter10), .b(gate541inter9), .O(gate541inter11));
  nor2  gate1019(.a(gate541inter11), .b(gate541inter6), .O(gate541inter12));
  nand2 gate1020(.a(gate541inter12), .b(gate541inter1), .O(N1838));
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );

  xor2  gate2141(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate2142(.a(gate546inter0), .b(s_180), .O(gate546inter1));
  and2  gate2143(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate2144(.a(s_180), .O(gate546inter3));
  inv1  gate2145(.a(s_181), .O(gate546inter4));
  nand2 gate2146(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate2147(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate2148(.a(N1319), .O(gate546inter7));
  inv1  gate2149(.a(N1827), .O(gate546inter8));
  nand2 gate2150(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate2151(.a(s_181), .b(gate546inter3), .O(gate546inter10));
  nor2  gate2152(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate2153(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate2154(.a(gate546inter12), .b(gate546inter1), .O(N1852));

  xor2  gate1539(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate1540(.a(gate547inter0), .b(s_94), .O(gate547inter1));
  and2  gate1541(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate1542(.a(s_94), .O(gate547inter3));
  inv1  gate1543(.a(s_95), .O(gate547inter4));
  nand2 gate1544(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate1545(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate1546(.a(N1815), .O(gate547inter7));
  inv1  gate1547(.a(N1707), .O(gate547inter8));
  nand2 gate1548(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate1549(.a(s_95), .b(gate547inter3), .O(gate547inter10));
  nor2  gate1550(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate1551(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate1552(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );

  xor2  gate3009(.a(N290), .b(N1798), .O(gate550inter0));
  nand2 gate3010(.a(gate550inter0), .b(s_304), .O(gate550inter1));
  and2  gate3011(.a(N290), .b(N1798), .O(gate550inter2));
  inv1  gate3012(.a(s_304), .O(gate550inter3));
  inv1  gate3013(.a(s_305), .O(gate550inter4));
  nand2 gate3014(.a(gate550inter4), .b(gate550inter3), .O(gate550inter5));
  nor2  gate3015(.a(gate550inter5), .b(gate550inter2), .O(gate550inter6));
  inv1  gate3016(.a(N1798), .O(gate550inter7));
  inv1  gate3017(.a(N290), .O(gate550inter8));
  nand2 gate3018(.a(gate550inter8), .b(gate550inter7), .O(gate550inter9));
  nand2 gate3019(.a(s_305), .b(gate550inter3), .O(gate550inter10));
  nor2  gate3020(.a(gate550inter10), .b(gate550inter9), .O(gate550inter11));
  nor2  gate3021(.a(gate550inter11), .b(gate550inter6), .O(gate550inter12));
  nand2 gate3022(.a(gate550inter12), .b(gate550inter1), .O(N1858));
inv1 gate551( .a(N1812), .O(N1864) );

  xor2  gate965(.a(N1728), .b(N1812), .O(gate552inter0));
  nand2 gate966(.a(gate552inter0), .b(s_12), .O(gate552inter1));
  and2  gate967(.a(N1728), .b(N1812), .O(gate552inter2));
  inv1  gate968(.a(s_12), .O(gate552inter3));
  inv1  gate969(.a(s_13), .O(gate552inter4));
  nand2 gate970(.a(gate552inter4), .b(gate552inter3), .O(gate552inter5));
  nor2  gate971(.a(gate552inter5), .b(gate552inter2), .O(gate552inter6));
  inv1  gate972(.a(N1812), .O(gate552inter7));
  inv1  gate973(.a(N1728), .O(gate552inter8));
  nand2 gate974(.a(gate552inter8), .b(gate552inter7), .O(gate552inter9));
  nand2 gate975(.a(s_13), .b(gate552inter3), .O(gate552inter10));
  nor2  gate976(.a(gate552inter10), .b(gate552inter9), .O(gate552inter11));
  nor2  gate977(.a(gate552inter11), .b(gate552inter6), .O(gate552inter12));
  nand2 gate978(.a(gate552inter12), .b(gate552inter1), .O(N1865));
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );

  xor2  gate1483(.a(N1849), .b(N1823), .O(gate558inter0));
  nand2 gate1484(.a(gate558inter0), .b(s_86), .O(gate558inter1));
  and2  gate1485(.a(N1849), .b(N1823), .O(gate558inter2));
  inv1  gate1486(.a(s_86), .O(gate558inter3));
  inv1  gate1487(.a(s_87), .O(gate558inter4));
  nand2 gate1488(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate1489(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate1490(.a(N1823), .O(gate558inter7));
  inv1  gate1491(.a(N1849), .O(gate558inter8));
  nand2 gate1492(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate1493(.a(s_87), .b(gate558inter3), .O(gate558inter10));
  nor2  gate1494(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate1495(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate1496(.a(gate558inter12), .b(gate558inter1), .O(N1879));

  xor2  gate3149(.a(N1768), .b(N1841), .O(gate559inter0));
  nand2 gate3150(.a(gate559inter0), .b(s_324), .O(gate559inter1));
  and2  gate3151(.a(N1768), .b(N1841), .O(gate559inter2));
  inv1  gate3152(.a(s_324), .O(gate559inter3));
  inv1  gate3153(.a(s_325), .O(gate559inter4));
  nand2 gate3154(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate3155(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate3156(.a(N1841), .O(gate559inter7));
  inv1  gate3157(.a(N1768), .O(gate559inter8));
  nand2 gate3158(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate3159(.a(s_325), .b(gate559inter3), .O(gate559inter10));
  nor2  gate3160(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate3161(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate3162(.a(gate559inter12), .b(gate559inter1), .O(N1882));
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );

  xor2  gate1189(.a(N290), .b(N1830), .O(gate563inter0));
  nand2 gate1190(.a(gate563inter0), .b(s_44), .O(gate563inter1));
  and2  gate1191(.a(N290), .b(N1830), .O(gate563inter2));
  inv1  gate1192(.a(s_44), .O(gate563inter3));
  inv1  gate1193(.a(s_45), .O(gate563inter4));
  nand2 gate1194(.a(gate563inter4), .b(gate563inter3), .O(gate563inter5));
  nor2  gate1195(.a(gate563inter5), .b(gate563inter2), .O(gate563inter6));
  inv1  gate1196(.a(N1830), .O(gate563inter7));
  inv1  gate1197(.a(N290), .O(gate563inter8));
  nand2 gate1198(.a(gate563inter8), .b(gate563inter7), .O(gate563inter9));
  nand2 gate1199(.a(s_45), .b(gate563inter3), .O(gate563inter10));
  nor2  gate1200(.a(gate563inter10), .b(gate563inter9), .O(gate563inter11));
  nor2  gate1201(.a(gate563inter11), .b(gate563inter6), .O(gate563inter12));
  nand2 gate1202(.a(gate563inter12), .b(gate563inter1), .O(N1889));
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );

  xor2  gate2015(.a(N1864), .b(N1640), .O(gate566inter0));
  nand2 gate2016(.a(gate566inter0), .b(s_162), .O(gate566inter1));
  and2  gate2017(.a(N1864), .b(N1640), .O(gate566inter2));
  inv1  gate2018(.a(s_162), .O(gate566inter3));
  inv1  gate2019(.a(s_163), .O(gate566inter4));
  nand2 gate2020(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate2021(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate2022(.a(N1640), .O(gate566inter7));
  inv1  gate2023(.a(N1864), .O(gate566inter8));
  nand2 gate2024(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate2025(.a(s_163), .b(gate566inter3), .O(gate566inter10));
  nor2  gate2026(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate2027(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate2028(.a(gate566inter12), .b(gate566inter1), .O(N1897));
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );

  xor2  gate2183(.a(N1883), .b(N1717), .O(gate570inter0));
  nand2 gate2184(.a(gate570inter0), .b(s_186), .O(gate570inter1));
  and2  gate2185(.a(N1883), .b(N1717), .O(gate570inter2));
  inv1  gate2186(.a(s_186), .O(gate570inter3));
  inv1  gate2187(.a(s_187), .O(gate570inter4));
  nand2 gate2188(.a(gate570inter4), .b(gate570inter3), .O(gate570inter5));
  nor2  gate2189(.a(gate570inter5), .b(gate570inter2), .O(gate570inter6));
  inv1  gate2190(.a(N1717), .O(gate570inter7));
  inv1  gate2191(.a(N1883), .O(gate570inter8));
  nand2 gate2192(.a(gate570inter8), .b(gate570inter7), .O(gate570inter9));
  nand2 gate2193(.a(s_187), .b(gate570inter3), .O(gate570inter10));
  nor2  gate2194(.a(gate570inter10), .b(gate570inter9), .O(gate570inter11));
  nor2  gate2195(.a(gate570inter11), .b(gate570inter6), .O(gate570inter12));
  nand2 gate2196(.a(gate570inter12), .b(gate570inter1), .O(N1911));
inv1 gate571( .a(N1884), .O(N1912) );

  xor2  gate2393(.a(N1885), .b(N1855), .O(gate572inter0));
  nand2 gate2394(.a(gate572inter0), .b(s_216), .O(gate572inter1));
  and2  gate2395(.a(N1885), .b(N1855), .O(gate572inter2));
  inv1  gate2396(.a(s_216), .O(gate572inter3));
  inv1  gate2397(.a(s_217), .O(gate572inter4));
  nand2 gate2398(.a(gate572inter4), .b(gate572inter3), .O(gate572inter5));
  nor2  gate2399(.a(gate572inter5), .b(gate572inter2), .O(gate572inter6));
  inv1  gate2400(.a(N1855), .O(gate572inter7));
  inv1  gate2401(.a(N1885), .O(gate572inter8));
  nand2 gate2402(.a(gate572inter8), .b(gate572inter7), .O(gate572inter9));
  nand2 gate2403(.a(s_217), .b(gate572inter3), .O(gate572inter10));
  nor2  gate2404(.a(gate572inter10), .b(gate572inter9), .O(gate572inter11));
  nor2  gate2405(.a(gate572inter11), .b(gate572inter6), .O(gate572inter12));
  nand2 gate2406(.a(gate572inter12), .b(gate572inter1), .O(N1913));
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );

  xor2  gate1231(.a(N920), .b(N1869), .O(gate576inter0));
  nand2 gate1232(.a(gate576inter0), .b(s_50), .O(gate576inter1));
  and2  gate1233(.a(N920), .b(N1869), .O(gate576inter2));
  inv1  gate1234(.a(s_50), .O(gate576inter3));
  inv1  gate1235(.a(s_51), .O(gate576inter4));
  nand2 gate1236(.a(gate576inter4), .b(gate576inter3), .O(gate576inter5));
  nor2  gate1237(.a(gate576inter5), .b(gate576inter2), .O(gate576inter6));
  inv1  gate1238(.a(N1869), .O(gate576inter7));
  inv1  gate1239(.a(N920), .O(gate576inter8));
  nand2 gate1240(.a(gate576inter8), .b(gate576inter7), .O(gate576inter9));
  nand2 gate1241(.a(s_51), .b(gate576inter3), .O(gate576inter10));
  nor2  gate1242(.a(gate576inter10), .b(gate576inter9), .O(gate576inter11));
  nor2  gate1243(.a(gate576inter11), .b(gate576inter6), .O(gate576inter12));
  nand2 gate1244(.a(gate576inter12), .b(gate576inter1), .O(N1921));
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate2841(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate2842(.a(gate579inter0), .b(s_280), .O(gate579inter1));
  and2  gate2843(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate2844(.a(s_280), .O(gate579inter3));
  inv1  gate2845(.a(s_281), .O(gate579inter4));
  nand2 gate2846(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate2847(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate2848(.a(N1714), .O(gate579inter7));
  inv1  gate2849(.a(N1895), .O(gate579inter8));
  nand2 gate2850(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate2851(.a(s_281), .b(gate579inter3), .O(gate579inter10));
  nor2  gate2852(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate2853(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate2854(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate2309(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate2310(.a(gate596inter0), .b(s_204), .O(gate596inter1));
  and2  gate2311(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate2312(.a(s_204), .O(gate596inter3));
  inv1  gate2313(.a(s_205), .O(gate596inter4));
  nand2 gate2314(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate2315(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate2316(.a(N1930), .O(gate596inter7));
  inv1  gate2317(.a(N917), .O(gate596inter8));
  nand2 gate2318(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate2319(.a(s_205), .b(gate596inter3), .O(gate596inter10));
  nor2  gate2320(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate2321(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate2322(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );

  xor2  gate2743(.a(N918), .b(N1927), .O(gate598inter0));
  nand2 gate2744(.a(gate598inter0), .b(s_266), .O(gate598inter1));
  and2  gate2745(.a(N918), .b(N1927), .O(gate598inter2));
  inv1  gate2746(.a(s_266), .O(gate598inter3));
  inv1  gate2747(.a(s_267), .O(gate598inter4));
  nand2 gate2748(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate2749(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate2750(.a(N1927), .O(gate598inter7));
  inv1  gate2751(.a(N918), .O(gate598inter8));
  nand2 gate2752(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate2753(.a(s_267), .b(gate598inter3), .O(gate598inter10));
  nor2  gate2754(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate2755(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate2756(.a(gate598inter12), .b(gate598inter1), .O(N1977));
inv1 gate599( .a(N1927), .O(N1978) );

  xor2  gate1889(.a(N1941), .b(N1919), .O(gate600inter0));
  nand2 gate1890(.a(gate600inter0), .b(s_144), .O(gate600inter1));
  and2  gate1891(.a(N1941), .b(N1919), .O(gate600inter2));
  inv1  gate1892(.a(s_144), .O(gate600inter3));
  inv1  gate1893(.a(s_145), .O(gate600inter4));
  nand2 gate1894(.a(gate600inter4), .b(gate600inter3), .O(gate600inter5));
  nor2  gate1895(.a(gate600inter5), .b(gate600inter2), .O(gate600inter6));
  inv1  gate1896(.a(N1919), .O(gate600inter7));
  inv1  gate1897(.a(N1941), .O(gate600inter8));
  nand2 gate1898(.a(gate600inter8), .b(gate600inter7), .O(gate600inter9));
  nand2 gate1899(.a(s_145), .b(gate600inter3), .O(gate600inter10));
  nor2  gate1900(.a(gate600inter10), .b(gate600inter9), .O(gate600inter11));
  nor2  gate1901(.a(gate600inter11), .b(gate600inter6), .O(gate600inter12));
  nand2 gate1902(.a(gate600inter12), .b(gate600inter1), .O(N1979));
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );

  xor2  gate1399(.a(N1351), .b(N1950), .O(gate610inter0));
  nand2 gate1400(.a(gate610inter0), .b(s_74), .O(gate610inter1));
  and2  gate1401(.a(N1351), .b(N1950), .O(gate610inter2));
  inv1  gate1402(.a(s_74), .O(gate610inter3));
  inv1  gate1403(.a(s_75), .O(gate610inter4));
  nand2 gate1404(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate1405(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate1406(.a(N1950), .O(gate610inter7));
  inv1  gate1407(.a(N1351), .O(gate610inter8));
  nand2 gate1408(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate1409(.a(s_75), .b(gate610inter3), .O(gate610inter10));
  nor2  gate1410(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate1411(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate1412(.a(gate610inter12), .b(gate610inter1), .O(N2006));
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate1385(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate1386(.a(gate612inter0), .b(s_72), .O(gate612inter1));
  and2  gate1387(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate1388(.a(s_72), .O(gate612inter3));
  inv1  gate1389(.a(s_73), .O(gate612inter4));
  nand2 gate1390(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate1391(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate1392(.a(N673), .O(gate612inter7));
  inv1  gate1393(.a(N1976), .O(gate612inter8));
  nand2 gate1394(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate1395(.a(s_73), .b(gate612inter3), .O(gate612inter10));
  nor2  gate1396(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate1397(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate1398(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );

  xor2  gate1693(.a(N1923), .b(N1958), .O(gate616inter0));
  nand2 gate1694(.a(gate616inter0), .b(s_116), .O(gate616inter1));
  and2  gate1695(.a(N1923), .b(N1958), .O(gate616inter2));
  inv1  gate1696(.a(s_116), .O(gate616inter3));
  inv1  gate1697(.a(s_117), .O(gate616inter4));
  nand2 gate1698(.a(gate616inter4), .b(gate616inter3), .O(gate616inter5));
  nor2  gate1699(.a(gate616inter5), .b(gate616inter2), .O(gate616inter6));
  inv1  gate1700(.a(N1958), .O(gate616inter7));
  inv1  gate1701(.a(N1923), .O(gate616inter8));
  nand2 gate1702(.a(gate616inter8), .b(gate616inter7), .O(gate616inter9));
  nand2 gate1703(.a(s_117), .b(gate616inter3), .O(gate616inter10));
  nor2  gate1704(.a(gate616inter10), .b(gate616inter9), .O(gate616inter11));
  nor2  gate1705(.a(gate616inter11), .b(gate616inter6), .O(gate616inter12));
  nand2 gate1706(.a(gate616inter12), .b(gate616inter1), .O(N2014));
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );

  xor2  gate2197(.a(N1999), .b(N1898), .O(gate621inter0));
  nand2 gate2198(.a(gate621inter0), .b(s_188), .O(gate621inter1));
  and2  gate2199(.a(N1999), .b(N1898), .O(gate621inter2));
  inv1  gate2200(.a(s_188), .O(gate621inter3));
  inv1  gate2201(.a(s_189), .O(gate621inter4));
  nand2 gate2202(.a(gate621inter4), .b(gate621inter3), .O(gate621inter5));
  nor2  gate2203(.a(gate621inter5), .b(gate621inter2), .O(gate621inter6));
  inv1  gate2204(.a(N1898), .O(gate621inter7));
  inv1  gate2205(.a(N1999), .O(gate621inter8));
  nand2 gate2206(.a(gate621inter8), .b(gate621inter7), .O(gate621inter9));
  nand2 gate2207(.a(s_189), .b(gate621inter3), .O(gate621inter10));
  nor2  gate2208(.a(gate621inter10), .b(gate621inter9), .O(gate621inter11));
  nor2  gate2209(.a(gate621inter11), .b(gate621inter6), .O(gate621inter12));
  nand2 gate2210(.a(gate621inter12), .b(gate621inter1), .O(N2020));
inv1 gate622( .a(N1987), .O(N2021) );

  xor2  gate1735(.a(N1591), .b(N1987), .O(gate623inter0));
  nand2 gate1736(.a(gate623inter0), .b(s_122), .O(gate623inter1));
  and2  gate1737(.a(N1591), .b(N1987), .O(gate623inter2));
  inv1  gate1738(.a(s_122), .O(gate623inter3));
  inv1  gate1739(.a(s_123), .O(gate623inter4));
  nand2 gate1740(.a(gate623inter4), .b(gate623inter3), .O(gate623inter5));
  nor2  gate1741(.a(gate623inter5), .b(gate623inter2), .O(gate623inter6));
  inv1  gate1742(.a(N1987), .O(gate623inter7));
  inv1  gate1743(.a(N1591), .O(gate623inter8));
  nand2 gate1744(.a(gate623inter8), .b(gate623inter7), .O(gate623inter9));
  nand2 gate1745(.a(s_123), .b(gate623inter3), .O(gate623inter10));
  nor2  gate1746(.a(gate623inter10), .b(gate623inter9), .O(gate623inter11));
  nor2  gate1747(.a(gate623inter11), .b(gate623inter6), .O(gate623inter12));
  nand2 gate1748(.a(gate623inter12), .b(gate623inter1), .O(N2022));

  xor2  gate2379(.a(N2002), .b(N1440), .O(gate624inter0));
  nand2 gate2380(.a(gate624inter0), .b(s_214), .O(gate624inter1));
  and2  gate2381(.a(N2002), .b(N1440), .O(gate624inter2));
  inv1  gate2382(.a(s_214), .O(gate624inter3));
  inv1  gate2383(.a(s_215), .O(gate624inter4));
  nand2 gate2384(.a(gate624inter4), .b(gate624inter3), .O(gate624inter5));
  nor2  gate2385(.a(gate624inter5), .b(gate624inter2), .O(gate624inter6));
  inv1  gate2386(.a(N1440), .O(gate624inter7));
  inv1  gate2387(.a(N2002), .O(gate624inter8));
  nand2 gate2388(.a(gate624inter8), .b(gate624inter7), .O(gate624inter9));
  nand2 gate2389(.a(s_215), .b(gate624inter3), .O(gate624inter10));
  nor2  gate2390(.a(gate624inter10), .b(gate624inter9), .O(gate624inter11));
  nor2  gate2391(.a(gate624inter11), .b(gate624inter6), .O(gate624inter12));
  nand2 gate2392(.a(gate624inter12), .b(gate624inter1), .O(N2023));
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate1749(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate1750(.a(gate633inter0), .b(s_124), .O(gate633inter1));
  and2  gate1751(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate1752(.a(s_124), .O(gate633inter3));
  inv1  gate1753(.a(s_125), .O(gate633inter4));
  nand2 gate1754(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate1755(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate1756(.a(N2020), .O(gate633inter7));
  inv1  gate1757(.a(N2000), .O(gate633inter8));
  nand2 gate1758(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate1759(.a(s_125), .b(gate633inter3), .O(gate633inter10));
  nor2  gate1760(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate1761(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate1762(.a(gate633inter12), .b(gate633inter1), .O(N2038));

  xor2  gate1791(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate1792(.a(gate634inter0), .b(s_130), .O(gate634inter1));
  and2  gate1793(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate1794(.a(s_130), .O(gate634inter3));
  inv1  gate1795(.a(s_131), .O(gate634inter4));
  nand2 gate1796(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate1797(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate1798(.a(N1534), .O(gate634inter7));
  inv1  gate1799(.a(N2021), .O(gate634inter8));
  nand2 gate1800(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate1801(.a(s_131), .b(gate634inter3), .O(gate634inter10));
  nor2  gate1802(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate1803(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate1804(.a(gate634inter12), .b(gate634inter1), .O(N2039));

  xor2  gate1455(.a(N2003), .b(N2023), .O(gate635inter0));
  nand2 gate1456(.a(gate635inter0), .b(s_82), .O(gate635inter1));
  and2  gate1457(.a(N2003), .b(N2023), .O(gate635inter2));
  inv1  gate1458(.a(s_82), .O(gate635inter3));
  inv1  gate1459(.a(s_83), .O(gate635inter4));
  nand2 gate1460(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate1461(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate1462(.a(N2023), .O(gate635inter7));
  inv1  gate1463(.a(N2003), .O(gate635inter8));
  nand2 gate1464(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate1465(.a(s_83), .b(gate635inter3), .O(gate635inter10));
  nor2  gate1466(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate1467(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate1468(.a(gate635inter12), .b(gate635inter1), .O(N2040));

  xor2  gate3107(.a(N2024), .b(N2004), .O(gate636inter0));
  nand2 gate3108(.a(gate636inter0), .b(s_318), .O(gate636inter1));
  and2  gate3109(.a(N2024), .b(N2004), .O(gate636inter2));
  inv1  gate3110(.a(s_318), .O(gate636inter3));
  inv1  gate3111(.a(s_319), .O(gate636inter4));
  nand2 gate3112(.a(gate636inter4), .b(gate636inter3), .O(gate636inter5));
  nor2  gate3113(.a(gate636inter5), .b(gate636inter2), .O(gate636inter6));
  inv1  gate3114(.a(N2004), .O(gate636inter7));
  inv1  gate3115(.a(N2024), .O(gate636inter8));
  nand2 gate3116(.a(gate636inter8), .b(gate636inter7), .O(gate636inter9));
  nand2 gate3117(.a(s_319), .b(gate636inter3), .O(gate636inter10));
  nor2  gate3118(.a(gate636inter10), .b(gate636inter9), .O(gate636inter11));
  nor2  gate3119(.a(gate636inter11), .b(gate636inter6), .O(gate636inter12));
  nand2 gate3120(.a(gate636inter12), .b(gate636inter1), .O(N2041));

  xor2  gate2785(.a(N2025), .b(N2006), .O(gate637inter0));
  nand2 gate2786(.a(gate637inter0), .b(s_272), .O(gate637inter1));
  and2  gate2787(.a(N2025), .b(N2006), .O(gate637inter2));
  inv1  gate2788(.a(s_272), .O(gate637inter3));
  inv1  gate2789(.a(s_273), .O(gate637inter4));
  nand2 gate2790(.a(gate637inter4), .b(gate637inter3), .O(gate637inter5));
  nor2  gate2791(.a(gate637inter5), .b(gate637inter2), .O(gate637inter6));
  inv1  gate2792(.a(N2006), .O(gate637inter7));
  inv1  gate2793(.a(N2025), .O(gate637inter8));
  nand2 gate2794(.a(gate637inter8), .b(gate637inter7), .O(gate637inter9));
  nand2 gate2795(.a(s_273), .b(gate637inter3), .O(gate637inter10));
  nor2  gate2796(.a(gate637inter10), .b(gate637inter9), .O(gate637inter11));
  nor2  gate2797(.a(gate637inter11), .b(gate637inter6), .O(gate637inter12));
  nand2 gate2798(.a(gate637inter12), .b(gate637inter1), .O(N2042));
inv1 gate638( .a(N2026), .O(N2047) );

  xor2  gate2281(.a(N2014), .b(N2036), .O(gate639inter0));
  nand2 gate2282(.a(gate639inter0), .b(s_200), .O(gate639inter1));
  and2  gate2283(.a(N2014), .b(N2036), .O(gate639inter2));
  inv1  gate2284(.a(s_200), .O(gate639inter3));
  inv1  gate2285(.a(s_201), .O(gate639inter4));
  nand2 gate2286(.a(gate639inter4), .b(gate639inter3), .O(gate639inter5));
  nor2  gate2287(.a(gate639inter5), .b(gate639inter2), .O(gate639inter6));
  inv1  gate2288(.a(N2036), .O(gate639inter7));
  inv1  gate2289(.a(N2014), .O(gate639inter8));
  nand2 gate2290(.a(gate639inter8), .b(gate639inter7), .O(gate639inter9));
  nand2 gate2291(.a(s_201), .b(gate639inter3), .O(gate639inter10));
  nor2  gate2292(.a(gate639inter10), .b(gate639inter9), .O(gate639inter11));
  nor2  gate2293(.a(gate639inter11), .b(gate639inter6), .O(gate639inter12));
  nand2 gate2294(.a(gate639inter12), .b(gate639inter1), .O(N2052));
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );

  xor2  gate1609(.a(N290), .b(N2060), .O(gate649inter0));
  nand2 gate1610(.a(gate649inter0), .b(s_104), .O(gate649inter1));
  and2  gate1611(.a(N290), .b(N2060), .O(gate649inter2));
  inv1  gate1612(.a(s_104), .O(gate649inter3));
  inv1  gate1613(.a(s_105), .O(gate649inter4));
  nand2 gate1614(.a(gate649inter4), .b(gate649inter3), .O(gate649inter5));
  nor2  gate1615(.a(gate649inter5), .b(gate649inter2), .O(gate649inter6));
  inv1  gate1616(.a(N2060), .O(gate649inter7));
  inv1  gate1617(.a(N290), .O(gate649inter8));
  nand2 gate1618(.a(gate649inter8), .b(gate649inter7), .O(gate649inter9));
  nand2 gate1619(.a(s_105), .b(gate649inter3), .O(gate649inter10));
  nor2  gate1620(.a(gate649inter10), .b(gate649inter9), .O(gate649inter11));
  nor2  gate1621(.a(gate649inter11), .b(gate649inter6), .O(gate649inter12));
  nand2 gate1622(.a(gate649inter12), .b(gate649inter1), .O(N2078));

  xor2  gate2981(.a(N290), .b(N2061), .O(gate650inter0));
  nand2 gate2982(.a(gate650inter0), .b(s_300), .O(gate650inter1));
  and2  gate2983(.a(N290), .b(N2061), .O(gate650inter2));
  inv1  gate2984(.a(s_300), .O(gate650inter3));
  inv1  gate2985(.a(s_301), .O(gate650inter4));
  nand2 gate2986(.a(gate650inter4), .b(gate650inter3), .O(gate650inter5));
  nor2  gate2987(.a(gate650inter5), .b(gate650inter2), .O(gate650inter6));
  inv1  gate2988(.a(N2061), .O(gate650inter7));
  inv1  gate2989(.a(N290), .O(gate650inter8));
  nand2 gate2990(.a(gate650inter8), .b(gate650inter7), .O(gate650inter9));
  nand2 gate2991(.a(s_301), .b(gate650inter3), .O(gate650inter10));
  nor2  gate2992(.a(gate650inter10), .b(gate650inter9), .O(gate650inter11));
  nor2  gate2993(.a(gate650inter11), .b(gate650inter6), .O(gate650inter12));
  nand2 gate2994(.a(gate650inter12), .b(gate650inter1), .O(N2081));
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );

  xor2  gate2225(.a(N915), .b(N2151), .O(gate663inter0));
  nand2 gate2226(.a(gate663inter0), .b(s_192), .O(gate663inter1));
  and2  gate2227(.a(N915), .b(N2151), .O(gate663inter2));
  inv1  gate2228(.a(s_192), .O(gate663inter3));
  inv1  gate2229(.a(s_193), .O(gate663inter4));
  nand2 gate2230(.a(gate663inter4), .b(gate663inter3), .O(gate663inter5));
  nor2  gate2231(.a(gate663inter5), .b(gate663inter2), .O(gate663inter6));
  inv1  gate2232(.a(N2151), .O(gate663inter7));
  inv1  gate2233(.a(N915), .O(gate663inter8));
  nand2 gate2234(.a(gate663inter8), .b(gate663inter7), .O(gate663inter9));
  nand2 gate2235(.a(s_193), .b(gate663inter3), .O(gate663inter10));
  nor2  gate2236(.a(gate663inter10), .b(gate663inter9), .O(gate663inter11));
  nor2  gate2237(.a(gate663inter11), .b(gate663inter6), .O(gate663inter12));
  nand2 gate2238(.a(gate663inter12), .b(gate663inter1), .O(N2214));
inv1 gate664( .a(N2151), .O(N2215) );

  xor2  gate2057(.a(N916), .b(N2148), .O(gate665inter0));
  nand2 gate2058(.a(gate665inter0), .b(s_168), .O(gate665inter1));
  and2  gate2059(.a(N916), .b(N2148), .O(gate665inter2));
  inv1  gate2060(.a(s_168), .O(gate665inter3));
  inv1  gate2061(.a(s_169), .O(gate665inter4));
  nand2 gate2062(.a(gate665inter4), .b(gate665inter3), .O(gate665inter5));
  nor2  gate2063(.a(gate665inter5), .b(gate665inter2), .O(gate665inter6));
  inv1  gate2064(.a(N2148), .O(gate665inter7));
  inv1  gate2065(.a(N916), .O(gate665inter8));
  nand2 gate2066(.a(gate665inter8), .b(gate665inter7), .O(gate665inter9));
  nand2 gate2067(.a(s_169), .b(gate665inter3), .O(gate665inter10));
  nor2  gate2068(.a(gate665inter10), .b(gate665inter9), .O(gate665inter11));
  nor2  gate2069(.a(gate665inter11), .b(gate665inter6), .O(gate665inter12));
  nand2 gate2070(.a(gate665inter12), .b(gate665inter1), .O(N2216));
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate2673(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate2674(.a(gate667inter0), .b(s_256), .O(gate667inter1));
  and2  gate2675(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate2676(.a(s_256), .O(gate667inter3));
  inv1  gate2677(.a(s_257), .O(gate667inter4));
  nand2 gate2678(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate2679(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate2680(.a(N2199), .O(gate667inter7));
  inv1  gate2681(.a(N1348), .O(gate667inter8));
  nand2 gate2682(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate2683(.a(s_257), .b(gate667inter3), .O(gate667inter10));
  nor2  gate2684(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate2685(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate2686(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );

  xor2  gate2603(.a(N1349), .b(N2196), .O(gate669inter0));
  nand2 gate2604(.a(gate669inter0), .b(s_246), .O(gate669inter1));
  and2  gate2605(.a(N1349), .b(N2196), .O(gate669inter2));
  inv1  gate2606(.a(s_246), .O(gate669inter3));
  inv1  gate2607(.a(s_247), .O(gate669inter4));
  nand2 gate2608(.a(gate669inter4), .b(gate669inter3), .O(gate669inter5));
  nor2  gate2609(.a(gate669inter5), .b(gate669inter2), .O(gate669inter6));
  inv1  gate2610(.a(N2196), .O(gate669inter7));
  inv1  gate2611(.a(N1349), .O(gate669inter8));
  nand2 gate2612(.a(gate669inter8), .b(gate669inter7), .O(gate669inter9));
  nand2 gate2613(.a(s_247), .b(gate669inter3), .O(gate669inter10));
  nor2  gate2614(.a(gate669inter10), .b(gate669inter9), .O(gate669inter11));
  nor2  gate2615(.a(gate669inter11), .b(gate669inter6), .O(gate669inter12));
  nand2 gate2616(.a(gate669inter12), .b(gate669inter1), .O(N2224));
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate3289(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate3290(.a(gate671inter0), .b(s_344), .O(gate671inter1));
  and2  gate3291(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate3292(.a(s_344), .O(gate671inter3));
  inv1  gate3293(.a(s_345), .O(gate671inter4));
  nand2 gate3294(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate3295(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate3296(.a(N2205), .O(gate671inter7));
  inv1  gate3297(.a(N913), .O(gate671inter8));
  nand2 gate3298(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate3299(.a(s_345), .b(gate671inter3), .O(gate671inter10));
  nor2  gate3300(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate3301(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate3302(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );

  xor2  gate3359(.a(N914), .b(N2202), .O(gate673inter0));
  nand2 gate3360(.a(gate673inter0), .b(s_354), .O(gate673inter1));
  and2  gate3361(.a(N914), .b(N2202), .O(gate673inter2));
  inv1  gate3362(.a(s_354), .O(gate673inter3));
  inv1  gate3363(.a(s_355), .O(gate673inter4));
  nand2 gate3364(.a(gate673inter4), .b(gate673inter3), .O(gate673inter5));
  nor2  gate3365(.a(gate673inter5), .b(gate673inter2), .O(gate673inter6));
  inv1  gate3366(.a(N2202), .O(gate673inter7));
  inv1  gate3367(.a(N914), .O(gate673inter8));
  nand2 gate3368(.a(gate673inter8), .b(gate673inter7), .O(gate673inter9));
  nand2 gate3369(.a(s_355), .b(gate673inter3), .O(gate673inter10));
  nor2  gate3370(.a(gate673inter10), .b(gate673inter9), .O(gate673inter11));
  nor2  gate3371(.a(gate673inter11), .b(gate673inter6), .O(gate673inter12));
  nand2 gate3372(.a(gate673inter12), .b(gate673inter1), .O(N2228));
inv1 gate674( .a(N2202), .O(N2229) );

  xor2  gate1259(.a(N2215), .b(N667), .O(gate675inter0));
  nand2 gate1260(.a(gate675inter0), .b(s_54), .O(gate675inter1));
  and2  gate1261(.a(N2215), .b(N667), .O(gate675inter2));
  inv1  gate1262(.a(s_54), .O(gate675inter3));
  inv1  gate1263(.a(s_55), .O(gate675inter4));
  nand2 gate1264(.a(gate675inter4), .b(gate675inter3), .O(gate675inter5));
  nor2  gate1265(.a(gate675inter5), .b(gate675inter2), .O(gate675inter6));
  inv1  gate1266(.a(N667), .O(gate675inter7));
  inv1  gate1267(.a(N2215), .O(gate675inter8));
  nand2 gate1268(.a(gate675inter8), .b(gate675inter7), .O(gate675inter9));
  nand2 gate1269(.a(s_55), .b(gate675inter3), .O(gate675inter10));
  nor2  gate1270(.a(gate675inter10), .b(gate675inter9), .O(gate675inter11));
  nor2  gate1271(.a(gate675inter11), .b(gate675inter6), .O(gate675inter12));
  nand2 gate1272(.a(gate675inter12), .b(gate675inter1), .O(N2230));

  xor2  gate2631(.a(N2217), .b(N664), .O(gate676inter0));
  nand2 gate2632(.a(gate676inter0), .b(s_250), .O(gate676inter1));
  and2  gate2633(.a(N2217), .b(N664), .O(gate676inter2));
  inv1  gate2634(.a(s_250), .O(gate676inter3));
  inv1  gate2635(.a(s_251), .O(gate676inter4));
  nand2 gate2636(.a(gate676inter4), .b(gate676inter3), .O(gate676inter5));
  nor2  gate2637(.a(gate676inter5), .b(gate676inter2), .O(gate676inter6));
  inv1  gate2638(.a(N664), .O(gate676inter7));
  inv1  gate2639(.a(N2217), .O(gate676inter8));
  nand2 gate2640(.a(gate676inter8), .b(gate676inter7), .O(gate676inter9));
  nand2 gate2641(.a(s_251), .b(gate676inter3), .O(gate676inter10));
  nor2  gate2642(.a(gate676inter10), .b(gate676inter9), .O(gate676inter11));
  nor2  gate2643(.a(gate676inter11), .b(gate676inter6), .O(gate676inter12));
  nand2 gate2644(.a(gate676inter12), .b(gate676inter1), .O(N2231));
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );

  xor2  gate3261(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate3262(.a(gate678inter0), .b(s_340), .O(gate678inter1));
  and2  gate3263(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate3264(.a(s_340), .O(gate678inter3));
  inv1  gate3265(.a(s_341), .O(gate678inter4));
  nand2 gate3266(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate3267(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate3268(.a(N1252), .O(gate678inter7));
  inv1  gate3269(.a(N2225), .O(gate678inter8));
  nand2 gate3270(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate3271(.a(s_341), .b(gate678inter3), .O(gate678inter10));
  nor2  gate3272(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate3273(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate3274(.a(gate678inter12), .b(gate678inter1), .O(N2233));

  xor2  gate937(.a(N2227), .b(N661), .O(gate679inter0));
  nand2 gate938(.a(gate679inter0), .b(s_8), .O(gate679inter1));
  and2  gate939(.a(N2227), .b(N661), .O(gate679inter2));
  inv1  gate940(.a(s_8), .O(gate679inter3));
  inv1  gate941(.a(s_9), .O(gate679inter4));
  nand2 gate942(.a(gate679inter4), .b(gate679inter3), .O(gate679inter5));
  nor2  gate943(.a(gate679inter5), .b(gate679inter2), .O(gate679inter6));
  inv1  gate944(.a(N661), .O(gate679inter7));
  inv1  gate945(.a(N2227), .O(gate679inter8));
  nand2 gate946(.a(gate679inter8), .b(gate679inter7), .O(gate679inter9));
  nand2 gate947(.a(s_9), .b(gate679inter3), .O(gate679inter10));
  nor2  gate948(.a(gate679inter10), .b(gate679inter9), .O(gate679inter11));
  nor2  gate949(.a(gate679inter11), .b(gate679inter6), .O(gate679inter12));
  nand2 gate950(.a(gate679inter12), .b(gate679inter1), .O(N2234));
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );

  xor2  gate2463(.a(N2230), .b(N2214), .O(gate681inter0));
  nand2 gate2464(.a(gate681inter0), .b(s_226), .O(gate681inter1));
  and2  gate2465(.a(N2230), .b(N2214), .O(gate681inter2));
  inv1  gate2466(.a(s_226), .O(gate681inter3));
  inv1  gate2467(.a(s_227), .O(gate681inter4));
  nand2 gate2468(.a(gate681inter4), .b(gate681inter3), .O(gate681inter5));
  nor2  gate2469(.a(gate681inter5), .b(gate681inter2), .O(gate681inter6));
  inv1  gate2470(.a(N2214), .O(gate681inter7));
  inv1  gate2471(.a(N2230), .O(gate681inter8));
  nand2 gate2472(.a(gate681inter8), .b(gate681inter7), .O(gate681inter9));
  nand2 gate2473(.a(s_227), .b(gate681inter3), .O(gate681inter10));
  nor2  gate2474(.a(gate681inter10), .b(gate681inter9), .O(gate681inter11));
  nor2  gate2475(.a(gate681inter11), .b(gate681inter6), .O(gate681inter12));
  nand2 gate2476(.a(gate681inter12), .b(gate681inter1), .O(N2236));
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );

  xor2  gate2771(.a(N2232), .b(N2222), .O(gate683inter0));
  nand2 gate2772(.a(gate683inter0), .b(s_270), .O(gate683inter1));
  and2  gate2773(.a(N2232), .b(N2222), .O(gate683inter2));
  inv1  gate2774(.a(s_270), .O(gate683inter3));
  inv1  gate2775(.a(s_271), .O(gate683inter4));
  nand2 gate2776(.a(gate683inter4), .b(gate683inter3), .O(gate683inter5));
  nor2  gate2777(.a(gate683inter5), .b(gate683inter2), .O(gate683inter6));
  inv1  gate2778(.a(N2222), .O(gate683inter7));
  inv1  gate2779(.a(N2232), .O(gate683inter8));
  nand2 gate2780(.a(gate683inter8), .b(gate683inter7), .O(gate683inter9));
  nand2 gate2781(.a(s_271), .b(gate683inter3), .O(gate683inter10));
  nor2  gate2782(.a(gate683inter10), .b(gate683inter9), .O(gate683inter11));
  nor2  gate2783(.a(gate683inter11), .b(gate683inter6), .O(gate683inter12));
  nand2 gate2784(.a(gate683inter12), .b(gate683inter1), .O(N2240));
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );

  xor2  gate2365(.a(N2235), .b(N2228), .O(gate686inter0));
  nand2 gate2366(.a(gate686inter0), .b(s_212), .O(gate686inter1));
  and2  gate2367(.a(N2235), .b(N2228), .O(gate686inter2));
  inv1  gate2368(.a(s_212), .O(gate686inter3));
  inv1  gate2369(.a(s_213), .O(gate686inter4));
  nand2 gate2370(.a(gate686inter4), .b(gate686inter3), .O(gate686inter5));
  nor2  gate2371(.a(gate686inter5), .b(gate686inter2), .O(gate686inter6));
  inv1  gate2372(.a(N2228), .O(gate686inter7));
  inv1  gate2373(.a(N2235), .O(gate686inter8));
  nand2 gate2374(.a(gate686inter8), .b(gate686inter7), .O(gate686inter9));
  nand2 gate2375(.a(s_213), .b(gate686inter3), .O(gate686inter10));
  nor2  gate2376(.a(gate686inter10), .b(gate686inter9), .O(gate686inter11));
  nor2  gate2377(.a(gate686inter11), .b(gate686inter6), .O(gate686inter12));
  nand2 gate2378(.a(gate686inter12), .b(gate686inter1), .O(N2245));
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );

  xor2  gate2813(.a(N534), .b(N2558), .O(gate750inter0));
  nand2 gate2814(.a(gate750inter0), .b(s_276), .O(gate750inter1));
  and2  gate2815(.a(N534), .b(N2558), .O(gate750inter2));
  inv1  gate2816(.a(s_276), .O(gate750inter3));
  inv1  gate2817(.a(s_277), .O(gate750inter4));
  nand2 gate2818(.a(gate750inter4), .b(gate750inter3), .O(gate750inter5));
  nor2  gate2819(.a(gate750inter5), .b(gate750inter2), .O(gate750inter6));
  inv1  gate2820(.a(N2558), .O(gate750inter7));
  inv1  gate2821(.a(N534), .O(gate750inter8));
  nand2 gate2822(.a(gate750inter8), .b(gate750inter7), .O(gate750inter9));
  nand2 gate2823(.a(s_277), .b(gate750inter3), .O(gate750inter10));
  nor2  gate2824(.a(gate750inter10), .b(gate750inter9), .O(gate750inter11));
  nor2  gate2825(.a(gate750inter11), .b(gate750inter6), .O(gate750inter12));
  nand2 gate2826(.a(gate750inter12), .b(gate750inter1), .O(N2669));
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate979(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate980(.a(gate754inter0), .b(s_14), .O(gate754inter1));
  and2  gate981(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate982(.a(s_14), .O(gate754inter3));
  inv1  gate983(.a(s_15), .O(gate754inter4));
  nand2 gate984(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate985(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate986(.a(N2564), .O(gate754inter7));
  inv1  gate987(.a(N536), .O(gate754inter8));
  nand2 gate988(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate989(.a(s_15), .b(gate754inter3), .O(gate754inter10));
  nor2  gate990(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate991(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate992(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate1091(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate1092(.a(gate756inter0), .b(s_30), .O(gate756inter1));
  and2  gate1093(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate1094(.a(s_30), .O(gate756inter3));
  inv1  gate1095(.a(s_31), .O(gate756inter4));
  nand2 gate1096(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate1097(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate1098(.a(N2567), .O(gate756inter7));
  inv1  gate1099(.a(N537), .O(gate756inter8));
  nand2 gate1100(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate1101(.a(s_31), .b(gate756inter3), .O(gate756inter10));
  nor2  gate1102(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate1103(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate1104(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );

  xor2  gate1175(.a(N548), .b(N2573), .O(gate760inter0));
  nand2 gate1176(.a(gate760inter0), .b(s_42), .O(gate760inter1));
  and2  gate1177(.a(N548), .b(N2573), .O(gate760inter2));
  inv1  gate1178(.a(s_42), .O(gate760inter3));
  inv1  gate1179(.a(s_43), .O(gate760inter4));
  nand2 gate1180(.a(gate760inter4), .b(gate760inter3), .O(gate760inter5));
  nor2  gate1181(.a(gate760inter5), .b(gate760inter2), .O(gate760inter6));
  inv1  gate1182(.a(N2573), .O(gate760inter7));
  inv1  gate1183(.a(N548), .O(gate760inter8));
  nand2 gate1184(.a(gate760inter8), .b(gate760inter7), .O(gate760inter9));
  nand2 gate1185(.a(s_43), .b(gate760inter3), .O(gate760inter10));
  nor2  gate1186(.a(gate760inter10), .b(gate760inter9), .O(gate760inter11));
  nor2  gate1187(.a(gate760inter11), .b(gate760inter6), .O(gate760inter12));
  nand2 gate1188(.a(gate760inter12), .b(gate760inter1), .O(N2688));
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );

  xor2  gate3471(.a(N2670), .b(N343), .O(gate765inter0));
  nand2 gate3472(.a(gate765inter0), .b(s_370), .O(gate765inter1));
  and2  gate3473(.a(N2670), .b(N343), .O(gate765inter2));
  inv1  gate3474(.a(s_370), .O(gate765inter3));
  inv1  gate3475(.a(s_371), .O(gate765inter4));
  nand2 gate3476(.a(gate765inter4), .b(gate765inter3), .O(gate765inter5));
  nor2  gate3477(.a(gate765inter5), .b(gate765inter2), .O(gate765inter6));
  inv1  gate3478(.a(N343), .O(gate765inter7));
  inv1  gate3479(.a(N2670), .O(gate765inter8));
  nand2 gate3480(.a(gate765inter8), .b(gate765inter7), .O(gate765inter9));
  nand2 gate3481(.a(s_371), .b(gate765inter3), .O(gate765inter10));
  nor2  gate3482(.a(gate765inter10), .b(gate765inter9), .O(gate765inter11));
  nor2  gate3483(.a(gate765inter11), .b(gate765inter6), .O(gate765inter12));
  nand2 gate3484(.a(gate765inter12), .b(gate765inter1), .O(N2720));

  xor2  gate2561(.a(N2672), .b(N346), .O(gate766inter0));
  nand2 gate2562(.a(gate766inter0), .b(s_240), .O(gate766inter1));
  and2  gate2563(.a(N2672), .b(N346), .O(gate766inter2));
  inv1  gate2564(.a(s_240), .O(gate766inter3));
  inv1  gate2565(.a(s_241), .O(gate766inter4));
  nand2 gate2566(.a(gate766inter4), .b(gate766inter3), .O(gate766inter5));
  nor2  gate2567(.a(gate766inter5), .b(gate766inter2), .O(gate766inter6));
  inv1  gate2568(.a(N346), .O(gate766inter7));
  inv1  gate2569(.a(N2672), .O(gate766inter8));
  nand2 gate2570(.a(gate766inter8), .b(gate766inter7), .O(gate766inter9));
  nand2 gate2571(.a(s_241), .b(gate766inter3), .O(gate766inter10));
  nor2  gate2572(.a(gate766inter10), .b(gate766inter9), .O(gate766inter11));
  nor2  gate2573(.a(gate766inter11), .b(gate766inter6), .O(gate766inter12));
  nand2 gate2574(.a(gate766inter12), .b(gate766inter1), .O(N2721));

  xor2  gate2267(.a(N2674), .b(N349), .O(gate767inter0));
  nand2 gate2268(.a(gate767inter0), .b(s_198), .O(gate767inter1));
  and2  gate2269(.a(N2674), .b(N349), .O(gate767inter2));
  inv1  gate2270(.a(s_198), .O(gate767inter3));
  inv1  gate2271(.a(s_199), .O(gate767inter4));
  nand2 gate2272(.a(gate767inter4), .b(gate767inter3), .O(gate767inter5));
  nor2  gate2273(.a(gate767inter5), .b(gate767inter2), .O(gate767inter6));
  inv1  gate2274(.a(N349), .O(gate767inter7));
  inv1  gate2275(.a(N2674), .O(gate767inter8));
  nand2 gate2276(.a(gate767inter8), .b(gate767inter7), .O(gate767inter9));
  nand2 gate2277(.a(s_199), .b(gate767inter3), .O(gate767inter10));
  nor2  gate2278(.a(gate767inter10), .b(gate767inter9), .O(gate767inter11));
  nor2  gate2279(.a(gate767inter11), .b(gate767inter6), .O(gate767inter12));
  nand2 gate2280(.a(gate767inter12), .b(gate767inter1), .O(N2722));

  xor2  gate2127(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate2128(.a(gate768inter0), .b(s_178), .O(gate768inter1));
  and2  gate2129(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate2130(.a(s_178), .O(gate768inter3));
  inv1  gate2131(.a(s_179), .O(gate768inter4));
  nand2 gate2132(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate2133(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate2134(.a(N352), .O(gate768inter7));
  inv1  gate2135(.a(N2676), .O(gate768inter8));
  nand2 gate2136(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate2137(.a(s_179), .b(gate768inter3), .O(gate768inter10));
  nor2  gate2138(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate2139(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate2140(.a(gate768inter12), .b(gate768inter1), .O(N2723));
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate1049(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate1050(.a(gate773inter0), .b(s_24), .O(gate773inter1));
  and2  gate1051(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate1052(.a(s_24), .O(gate773inter3));
  inv1  gate1053(.a(s_25), .O(gate773inter4));
  nand2 gate1054(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate1055(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate1056(.a(N2645), .O(gate773inter7));
  inv1  gate1057(.a(N540), .O(gate773inter8));
  nand2 gate1058(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate1059(.a(s_25), .b(gate773inter3), .O(gate773inter10));
  nor2  gate1060(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate1061(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate1062(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );

  xor2  gate1665(.a(N541), .b(N2648), .O(gate775inter0));
  nand2 gate1666(.a(gate775inter0), .b(s_112), .O(gate775inter1));
  and2  gate1667(.a(N541), .b(N2648), .O(gate775inter2));
  inv1  gate1668(.a(s_112), .O(gate775inter3));
  inv1  gate1669(.a(s_113), .O(gate775inter4));
  nand2 gate1670(.a(gate775inter4), .b(gate775inter3), .O(gate775inter5));
  nor2  gate1671(.a(gate775inter5), .b(gate775inter2), .O(gate775inter6));
  inv1  gate1672(.a(N2648), .O(gate775inter7));
  inv1  gate1673(.a(N541), .O(gate775inter8));
  nand2 gate1674(.a(gate775inter8), .b(gate775inter7), .O(gate775inter9));
  nand2 gate1675(.a(s_113), .b(gate775inter3), .O(gate775inter10));
  nor2  gate1676(.a(gate775inter10), .b(gate775inter9), .O(gate775inter11));
  nor2  gate1677(.a(gate775inter11), .b(gate775inter6), .O(gate775inter12));
  nand2 gate1678(.a(gate775inter12), .b(gate775inter1), .O(N2730));
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );

  xor2  gate1819(.a(N544), .b(N2655), .O(gate780inter0));
  nand2 gate1820(.a(gate780inter0), .b(s_134), .O(gate780inter1));
  and2  gate1821(.a(N544), .b(N2655), .O(gate780inter2));
  inv1  gate1822(.a(s_134), .O(gate780inter3));
  inv1  gate1823(.a(s_135), .O(gate780inter4));
  nand2 gate1824(.a(gate780inter4), .b(gate780inter3), .O(gate780inter5));
  nor2  gate1825(.a(gate780inter5), .b(gate780inter2), .O(gate780inter6));
  inv1  gate1826(.a(N2655), .O(gate780inter7));
  inv1  gate1827(.a(N544), .O(gate780inter8));
  nand2 gate1828(.a(gate780inter8), .b(gate780inter7), .O(gate780inter9));
  nand2 gate1829(.a(s_135), .b(gate780inter3), .O(gate780inter10));
  nor2  gate1830(.a(gate780inter10), .b(gate780inter9), .O(gate780inter11));
  nor2  gate1831(.a(gate780inter11), .b(gate780inter6), .O(gate780inter12));
  nand2 gate1832(.a(gate780inter12), .b(gate780inter1), .O(N2735));
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );

  xor2  gate2827(.a(N547), .b(N2664), .O(gate786inter0));
  nand2 gate2828(.a(gate786inter0), .b(s_278), .O(gate786inter1));
  and2  gate2829(.a(N547), .b(N2664), .O(gate786inter2));
  inv1  gate2830(.a(s_278), .O(gate786inter3));
  inv1  gate2831(.a(s_279), .O(gate786inter4));
  nand2 gate2832(.a(gate786inter4), .b(gate786inter3), .O(gate786inter5));
  nor2  gate2833(.a(gate786inter5), .b(gate786inter2), .O(gate786inter6));
  inv1  gate2834(.a(N2664), .O(gate786inter7));
  inv1  gate2835(.a(N547), .O(gate786inter8));
  nand2 gate2836(.a(gate786inter8), .b(gate786inter7), .O(gate786inter9));
  nand2 gate2837(.a(s_279), .b(gate786inter3), .O(gate786inter10));
  nor2  gate2838(.a(gate786inter10), .b(gate786inter9), .O(gate786inter11));
  nor2  gate2839(.a(gate786inter11), .b(gate786inter6), .O(gate786inter12));
  nand2 gate2840(.a(gate786inter12), .b(gate786inter1), .O(N2741));
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );

  xor2  gate1833(.a(N2691), .b(N388), .O(gate789inter0));
  nand2 gate1834(.a(gate789inter0), .b(s_136), .O(gate789inter1));
  and2  gate1835(.a(N2691), .b(N388), .O(gate789inter2));
  inv1  gate1836(.a(s_136), .O(gate789inter3));
  inv1  gate1837(.a(s_137), .O(gate789inter4));
  nand2 gate1838(.a(gate789inter4), .b(gate789inter3), .O(gate789inter5));
  nor2  gate1839(.a(gate789inter5), .b(gate789inter2), .O(gate789inter6));
  inv1  gate1840(.a(N388), .O(gate789inter7));
  inv1  gate1841(.a(N2691), .O(gate789inter8));
  nand2 gate1842(.a(gate789inter8), .b(gate789inter7), .O(gate789inter9));
  nand2 gate1843(.a(s_137), .b(gate789inter3), .O(gate789inter10));
  nor2  gate1844(.a(gate789inter10), .b(gate789inter9), .O(gate789inter11));
  nor2  gate1845(.a(gate789inter11), .b(gate789inter6), .O(gate789inter12));
  nand2 gate1846(.a(gate789inter12), .b(gate789inter1), .O(N2744));
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );

  xor2  gate1763(.a(N2720), .b(N2669), .O(gate794inter0));
  nand2 gate1764(.a(gate794inter0), .b(s_126), .O(gate794inter1));
  and2  gate1765(.a(N2720), .b(N2669), .O(gate794inter2));
  inv1  gate1766(.a(s_126), .O(gate794inter3));
  inv1  gate1767(.a(s_127), .O(gate794inter4));
  nand2 gate1768(.a(gate794inter4), .b(gate794inter3), .O(gate794inter5));
  nor2  gate1769(.a(gate794inter5), .b(gate794inter2), .O(gate794inter6));
  inv1  gate1770(.a(N2669), .O(gate794inter7));
  inv1  gate1771(.a(N2720), .O(gate794inter8));
  nand2 gate1772(.a(gate794inter8), .b(gate794inter7), .O(gate794inter9));
  nand2 gate1773(.a(s_127), .b(gate794inter3), .O(gate794inter10));
  nor2  gate1774(.a(gate794inter10), .b(gate794inter9), .O(gate794inter11));
  nor2  gate1775(.a(gate794inter11), .b(gate794inter6), .O(gate794inter12));
  nand2 gate1776(.a(gate794inter12), .b(gate794inter1), .O(N2753));
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );

  xor2  gate3163(.a(N2722), .b(N2673), .O(gate796inter0));
  nand2 gate3164(.a(gate796inter0), .b(s_326), .O(gate796inter1));
  and2  gate3165(.a(N2722), .b(N2673), .O(gate796inter2));
  inv1  gate3166(.a(s_326), .O(gate796inter3));
  inv1  gate3167(.a(s_327), .O(gate796inter4));
  nand2 gate3168(.a(gate796inter4), .b(gate796inter3), .O(gate796inter5));
  nor2  gate3169(.a(gate796inter5), .b(gate796inter2), .O(gate796inter6));
  inv1  gate3170(.a(N2673), .O(gate796inter7));
  inv1  gate3171(.a(N2722), .O(gate796inter8));
  nand2 gate3172(.a(gate796inter8), .b(gate796inter7), .O(gate796inter9));
  nand2 gate3173(.a(s_327), .b(gate796inter3), .O(gate796inter10));
  nor2  gate3174(.a(gate796inter10), .b(gate796inter9), .O(gate796inter11));
  nor2  gate3175(.a(gate796inter11), .b(gate796inter6), .O(gate796inter12));
  nand2 gate3176(.a(gate796inter12), .b(gate796inter1), .O(N2755));
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );

  xor2  gate1903(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate1904(.a(gate799inter0), .b(s_146), .O(gate799inter1));
  and2  gate1905(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate1906(.a(s_146), .O(gate799inter3));
  inv1  gate1907(.a(s_147), .O(gate799inter4));
  nand2 gate1908(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate1909(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate1910(.a(N358), .O(gate799inter7));
  inv1  gate1911(.a(N2727), .O(gate799inter8));
  nand2 gate1912(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate1913(.a(s_147), .b(gate799inter3), .O(gate799inter10));
  nor2  gate1914(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate1915(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate1916(.a(gate799inter12), .b(gate799inter1), .O(N2758));

  xor2  gate2799(.a(N2729), .b(N361), .O(gate800inter0));
  nand2 gate2800(.a(gate800inter0), .b(s_274), .O(gate800inter1));
  and2  gate2801(.a(N2729), .b(N361), .O(gate800inter2));
  inv1  gate2802(.a(s_274), .O(gate800inter3));
  inv1  gate2803(.a(s_275), .O(gate800inter4));
  nand2 gate2804(.a(gate800inter4), .b(gate800inter3), .O(gate800inter5));
  nor2  gate2805(.a(gate800inter5), .b(gate800inter2), .O(gate800inter6));
  inv1  gate2806(.a(N361), .O(gate800inter7));
  inv1  gate2807(.a(N2729), .O(gate800inter8));
  nand2 gate2808(.a(gate800inter8), .b(gate800inter7), .O(gate800inter9));
  nand2 gate2809(.a(s_275), .b(gate800inter3), .O(gate800inter10));
  nor2  gate2810(.a(gate800inter10), .b(gate800inter9), .O(gate800inter11));
  nor2  gate2811(.a(gate800inter11), .b(gate800inter6), .O(gate800inter12));
  nand2 gate2812(.a(gate800inter12), .b(gate800inter1), .O(N2759));

  xor2  gate3275(.a(N2731), .b(N364), .O(gate801inter0));
  nand2 gate3276(.a(gate801inter0), .b(s_342), .O(gate801inter1));
  and2  gate3277(.a(N2731), .b(N364), .O(gate801inter2));
  inv1  gate3278(.a(s_342), .O(gate801inter3));
  inv1  gate3279(.a(s_343), .O(gate801inter4));
  nand2 gate3280(.a(gate801inter4), .b(gate801inter3), .O(gate801inter5));
  nor2  gate3281(.a(gate801inter5), .b(gate801inter2), .O(gate801inter6));
  inv1  gate3282(.a(N364), .O(gate801inter7));
  inv1  gate3283(.a(N2731), .O(gate801inter8));
  nand2 gate3284(.a(gate801inter8), .b(gate801inter7), .O(gate801inter9));
  nand2 gate3285(.a(s_343), .b(gate801inter3), .O(gate801inter10));
  nor2  gate3286(.a(gate801inter10), .b(gate801inter9), .O(gate801inter11));
  nor2  gate3287(.a(gate801inter11), .b(gate801inter6), .O(gate801inter12));
  nand2 gate3288(.a(gate801inter12), .b(gate801inter1), .O(N2760));
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );

  xor2  gate2435(.a(N2736), .b(N373), .O(gate804inter0));
  nand2 gate2436(.a(gate804inter0), .b(s_222), .O(gate804inter1));
  and2  gate2437(.a(N2736), .b(N373), .O(gate804inter2));
  inv1  gate2438(.a(s_222), .O(gate804inter3));
  inv1  gate2439(.a(s_223), .O(gate804inter4));
  nand2 gate2440(.a(gate804inter4), .b(gate804inter3), .O(gate804inter5));
  nor2  gate2441(.a(gate804inter5), .b(gate804inter2), .O(gate804inter6));
  inv1  gate2442(.a(N373), .O(gate804inter7));
  inv1  gate2443(.a(N2736), .O(gate804inter8));
  nand2 gate2444(.a(gate804inter8), .b(gate804inter7), .O(gate804inter9));
  nand2 gate2445(.a(s_223), .b(gate804inter3), .O(gate804inter10));
  nor2  gate2446(.a(gate804inter10), .b(gate804inter9), .O(gate804inter11));
  nor2  gate2447(.a(gate804inter11), .b(gate804inter6), .O(gate804inter12));
  nand2 gate2448(.a(gate804inter12), .b(gate804inter1), .O(N2763));
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );

  xor2  gate2351(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate2352(.a(gate806inter0), .b(s_210), .O(gate806inter1));
  and2  gate2353(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate2354(.a(s_210), .O(gate806inter3));
  inv1  gate2355(.a(s_211), .O(gate806inter4));
  nand2 gate2356(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate2357(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate2358(.a(N379), .O(gate806inter7));
  inv1  gate2359(.a(N2740), .O(gate806inter8));
  nand2 gate2360(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate2361(.a(s_211), .b(gate806inter3), .O(gate806inter10));
  nor2  gate2362(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate2363(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate2364(.a(gate806inter12), .b(gate806inter1), .O(N2765));

  xor2  gate1637(.a(N2742), .b(N382), .O(gate807inter0));
  nand2 gate1638(.a(gate807inter0), .b(s_108), .O(gate807inter1));
  and2  gate1639(.a(N2742), .b(N382), .O(gate807inter2));
  inv1  gate1640(.a(s_108), .O(gate807inter3));
  inv1  gate1641(.a(s_109), .O(gate807inter4));
  nand2 gate1642(.a(gate807inter4), .b(gate807inter3), .O(gate807inter5));
  nor2  gate1643(.a(gate807inter5), .b(gate807inter2), .O(gate807inter6));
  inv1  gate1644(.a(N382), .O(gate807inter7));
  inv1  gate1645(.a(N2742), .O(gate807inter8));
  nand2 gate1646(.a(gate807inter8), .b(gate807inter7), .O(gate807inter9));
  nand2 gate1647(.a(s_109), .b(gate807inter3), .O(gate807inter10));
  nor2  gate1648(.a(gate807inter10), .b(gate807inter9), .O(gate807inter11));
  nor2  gate1649(.a(gate807inter11), .b(gate807inter6), .O(gate807inter12));
  nand2 gate1650(.a(gate807inter12), .b(gate807inter1), .O(N2766));
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );

  xor2  gate3205(.a(N2757), .b(N2724), .O(gate812inter0));
  nand2 gate3206(.a(gate812inter0), .b(s_332), .O(gate812inter1));
  and2  gate3207(.a(N2757), .b(N2724), .O(gate812inter2));
  inv1  gate3208(.a(s_332), .O(gate812inter3));
  inv1  gate3209(.a(s_333), .O(gate812inter4));
  nand2 gate3210(.a(gate812inter4), .b(gate812inter3), .O(gate812inter5));
  nor2  gate3211(.a(gate812inter5), .b(gate812inter2), .O(gate812inter6));
  inv1  gate3212(.a(N2724), .O(gate812inter7));
  inv1  gate3213(.a(N2757), .O(gate812inter8));
  nand2 gate3214(.a(gate812inter8), .b(gate812inter7), .O(gate812inter9));
  nand2 gate3215(.a(s_333), .b(gate812inter3), .O(gate812inter10));
  nor2  gate3216(.a(gate812inter10), .b(gate812inter9), .O(gate812inter11));
  nor2  gate3217(.a(gate812inter11), .b(gate812inter6), .O(gate812inter12));
  nand2 gate3218(.a(gate812inter12), .b(gate812inter1), .O(N2779));

  xor2  gate1315(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate1316(.a(gate813inter0), .b(s_62), .O(gate813inter1));
  and2  gate1317(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate1318(.a(s_62), .O(gate813inter3));
  inv1  gate1319(.a(s_63), .O(gate813inter4));
  nand2 gate1320(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate1321(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate1322(.a(N2726), .O(gate813inter7));
  inv1  gate1323(.a(N2758), .O(gate813inter8));
  nand2 gate1324(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate1325(.a(s_63), .b(gate813inter3), .O(gate813inter10));
  nor2  gate1326(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate1327(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate1328(.a(gate813inter12), .b(gate813inter1), .O(N2780));
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );

  xor2  gate1973(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate1974(.a(gate815inter0), .b(s_156), .O(gate815inter1));
  and2  gate1975(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate1976(.a(s_156), .O(gate815inter3));
  inv1  gate1977(.a(s_157), .O(gate815inter4));
  nand2 gate1978(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate1979(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate1980(.a(N2730), .O(gate815inter7));
  inv1  gate1981(.a(N2760), .O(gate815inter8));
  nand2 gate1982(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate1983(.a(s_157), .b(gate815inter3), .O(gate815inter10));
  nor2  gate1984(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate1985(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate1986(.a(gate815inter12), .b(gate815inter1), .O(N2782));

  xor2  gate1651(.a(N2761), .b(N2732), .O(gate816inter0));
  nand2 gate1652(.a(gate816inter0), .b(s_110), .O(gate816inter1));
  and2  gate1653(.a(N2761), .b(N2732), .O(gate816inter2));
  inv1  gate1654(.a(s_110), .O(gate816inter3));
  inv1  gate1655(.a(s_111), .O(gate816inter4));
  nand2 gate1656(.a(gate816inter4), .b(gate816inter3), .O(gate816inter5));
  nor2  gate1657(.a(gate816inter5), .b(gate816inter2), .O(gate816inter6));
  inv1  gate1658(.a(N2732), .O(gate816inter7));
  inv1  gate1659(.a(N2761), .O(gate816inter8));
  nand2 gate1660(.a(gate816inter8), .b(gate816inter7), .O(gate816inter9));
  nand2 gate1661(.a(s_111), .b(gate816inter3), .O(gate816inter10));
  nor2  gate1662(.a(gate816inter10), .b(gate816inter9), .O(gate816inter11));
  nor2  gate1663(.a(gate816inter11), .b(gate816inter6), .O(gate816inter12));
  nand2 gate1664(.a(gate816inter12), .b(gate816inter1), .O(N2783));

  xor2  gate1721(.a(N2763), .b(N2735), .O(gate817inter0));
  nand2 gate1722(.a(gate817inter0), .b(s_120), .O(gate817inter1));
  and2  gate1723(.a(N2763), .b(N2735), .O(gate817inter2));
  inv1  gate1724(.a(s_120), .O(gate817inter3));
  inv1  gate1725(.a(s_121), .O(gate817inter4));
  nand2 gate1726(.a(gate817inter4), .b(gate817inter3), .O(gate817inter5));
  nor2  gate1727(.a(gate817inter5), .b(gate817inter2), .O(gate817inter6));
  inv1  gate1728(.a(N2735), .O(gate817inter7));
  inv1  gate1729(.a(N2763), .O(gate817inter8));
  nand2 gate1730(.a(gate817inter8), .b(gate817inter7), .O(gate817inter9));
  nand2 gate1731(.a(s_121), .b(gate817inter3), .O(gate817inter10));
  nor2  gate1732(.a(gate817inter10), .b(gate817inter9), .O(gate817inter11));
  nor2  gate1733(.a(gate817inter11), .b(gate817inter6), .O(gate817inter12));
  nand2 gate1734(.a(gate817inter12), .b(gate817inter1), .O(N2784));
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );

  xor2  gate2939(.a(N2766), .b(N2741), .O(gate820inter0));
  nand2 gate2940(.a(gate820inter0), .b(s_294), .O(gate820inter1));
  and2  gate2941(.a(N2766), .b(N2741), .O(gate820inter2));
  inv1  gate2942(.a(s_294), .O(gate820inter3));
  inv1  gate2943(.a(s_295), .O(gate820inter4));
  nand2 gate2944(.a(gate820inter4), .b(gate820inter3), .O(gate820inter5));
  nor2  gate2945(.a(gate820inter5), .b(gate820inter2), .O(gate820inter6));
  inv1  gate2946(.a(N2741), .O(gate820inter7));
  inv1  gate2947(.a(N2766), .O(gate820inter8));
  nand2 gate2948(.a(gate820inter8), .b(gate820inter7), .O(gate820inter9));
  nand2 gate2949(.a(s_295), .b(gate820inter3), .O(gate820inter10));
  nor2  gate2950(.a(gate820inter10), .b(gate820inter9), .O(gate820inter11));
  nor2  gate2951(.a(gate820inter11), .b(gate820inter6), .O(gate820inter12));
  nand2 gate2952(.a(gate820inter12), .b(gate820inter1), .O(N2787));
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );

  xor2  gate3065(.a(N2750), .b(N2747), .O(gate822inter0));
  nand2 gate3066(.a(gate822inter0), .b(s_312), .O(gate822inter1));
  and2  gate3067(.a(N2750), .b(N2747), .O(gate822inter2));
  inv1  gate3068(.a(s_312), .O(gate822inter3));
  inv1  gate3069(.a(s_313), .O(gate822inter4));
  nand2 gate3070(.a(gate822inter4), .b(gate822inter3), .O(gate822inter5));
  nor2  gate3071(.a(gate822inter5), .b(gate822inter2), .O(gate822inter6));
  inv1  gate3072(.a(N2747), .O(gate822inter7));
  inv1  gate3073(.a(N2750), .O(gate822inter8));
  nand2 gate3074(.a(gate822inter8), .b(gate822inter7), .O(gate822inter9));
  nand2 gate3075(.a(s_313), .b(gate822inter3), .O(gate822inter10));
  nor2  gate3076(.a(gate822inter10), .b(gate822inter9), .O(gate822inter11));
  nor2  gate3077(.a(gate822inter11), .b(gate822inter6), .O(gate822inter12));
  nand2 gate3078(.a(gate822inter12), .b(gate822inter1), .O(N2789));
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );

  xor2  gate3429(.a(N2800), .b(N2384), .O(gate828inter0));
  nand2 gate3430(.a(gate828inter0), .b(s_364), .O(gate828inter1));
  and2  gate3431(.a(N2800), .b(N2384), .O(gate828inter2));
  inv1  gate3432(.a(s_364), .O(gate828inter3));
  inv1  gate3433(.a(s_365), .O(gate828inter4));
  nand2 gate3434(.a(gate828inter4), .b(gate828inter3), .O(gate828inter5));
  nor2  gate3435(.a(gate828inter5), .b(gate828inter2), .O(gate828inter6));
  inv1  gate3436(.a(N2384), .O(gate828inter7));
  inv1  gate3437(.a(N2800), .O(gate828inter8));
  nand2 gate3438(.a(gate828inter8), .b(gate828inter7), .O(gate828inter9));
  nand2 gate3439(.a(s_365), .b(gate828inter3), .O(gate828inter10));
  nor2  gate3440(.a(gate828inter10), .b(gate828inter9), .O(gate828inter11));
  nor2  gate3441(.a(gate828inter11), .b(gate828inter6), .O(gate828inter12));
  nand2 gate3442(.a(gate828inter12), .b(gate828inter1), .O(N2811));
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );

  xor2  gate2449(.a(N2810), .b(N1968), .O(gate835inter0));
  nand2 gate2450(.a(gate835inter0), .b(s_224), .O(gate835inter1));
  and2  gate2451(.a(N2810), .b(N1968), .O(gate835inter2));
  inv1  gate2452(.a(s_224), .O(gate835inter3));
  inv1  gate2453(.a(s_225), .O(gate835inter4));
  nand2 gate2454(.a(gate835inter4), .b(gate835inter3), .O(gate835inter5));
  nor2  gate2455(.a(gate835inter5), .b(gate835inter2), .O(gate835inter6));
  inv1  gate2456(.a(N1968), .O(gate835inter7));
  inv1  gate2457(.a(N2810), .O(gate835inter8));
  nand2 gate2458(.a(gate835inter8), .b(gate835inter7), .O(gate835inter9));
  nand2 gate2459(.a(s_225), .b(gate835inter3), .O(gate835inter10));
  nor2  gate2460(.a(gate835inter10), .b(gate835inter9), .O(gate835inter11));
  nor2  gate2461(.a(gate835inter11), .b(gate835inter6), .O(gate835inter12));
  nand2 gate2462(.a(gate835inter12), .b(gate835inter1), .O(N2828));
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );

  xor2  gate3051(.a(N2827), .b(N2807), .O(gate837inter0));
  nand2 gate3052(.a(gate837inter0), .b(s_310), .O(gate837inter1));
  and2  gate3053(.a(N2827), .b(N2807), .O(gate837inter2));
  inv1  gate3054(.a(s_310), .O(gate837inter3));
  inv1  gate3055(.a(s_311), .O(gate837inter4));
  nand2 gate3056(.a(gate837inter4), .b(gate837inter3), .O(gate837inter5));
  nor2  gate3057(.a(gate837inter5), .b(gate837inter2), .O(gate837inter6));
  inv1  gate3058(.a(N2807), .O(gate837inter7));
  inv1  gate3059(.a(N2827), .O(gate837inter8));
  nand2 gate3060(.a(gate837inter8), .b(gate837inter7), .O(gate837inter9));
  nand2 gate3061(.a(s_311), .b(gate837inter3), .O(gate837inter10));
  nor2  gate3062(.a(gate837inter10), .b(gate837inter9), .O(gate837inter11));
  nor2  gate3063(.a(gate837inter11), .b(gate837inter6), .O(gate837inter12));
  nand2 gate3064(.a(gate837inter12), .b(gate837inter1), .O(N2843));
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );

  xor2  gate923(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate924(.a(gate840inter0), .b(s_6), .O(gate840inter1));
  and2  gate925(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate926(.a(s_6), .O(gate840inter3));
  inv1  gate927(.a(s_7), .O(gate840inter4));
  nand2 gate928(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate929(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate930(.a(N2815), .O(gate840inter7));
  inv1  gate931(.a(N2077), .O(gate840inter8));
  nand2 gate932(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate933(.a(s_7), .b(gate840inter3), .O(gate840inter10));
  nor2  gate934(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate935(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate936(.a(gate840inter12), .b(gate840inter1), .O(N2851));

  xor2  gate2659(.a(N1915), .b(N2818), .O(gate841inter0));
  nand2 gate2660(.a(gate841inter0), .b(s_254), .O(gate841inter1));
  and2  gate2661(.a(N1915), .b(N2818), .O(gate841inter2));
  inv1  gate2662(.a(s_254), .O(gate841inter3));
  inv1  gate2663(.a(s_255), .O(gate841inter4));
  nand2 gate2664(.a(gate841inter4), .b(gate841inter3), .O(gate841inter5));
  nor2  gate2665(.a(gate841inter5), .b(gate841inter2), .O(gate841inter6));
  inv1  gate2666(.a(N2818), .O(gate841inter7));
  inv1  gate2667(.a(N1915), .O(gate841inter8));
  nand2 gate2668(.a(gate841inter8), .b(gate841inter7), .O(gate841inter9));
  nand2 gate2669(.a(s_255), .b(gate841inter3), .O(gate841inter10));
  nor2  gate2670(.a(gate841inter10), .b(gate841inter9), .O(gate841inter11));
  nor2  gate2671(.a(gate841inter11), .b(gate841inter6), .O(gate841inter12));
  nand2 gate2672(.a(gate841inter12), .b(gate841inter1), .O(N2852));
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );

  xor2  gate1105(.a(N1938), .b(N2824), .O(gate843inter0));
  nand2 gate1106(.a(gate843inter0), .b(s_32), .O(gate843inter1));
  and2  gate1107(.a(N1938), .b(N2824), .O(gate843inter2));
  inv1  gate1108(.a(s_32), .O(gate843inter3));
  inv1  gate1109(.a(s_33), .O(gate843inter4));
  nand2 gate1110(.a(gate843inter4), .b(gate843inter3), .O(gate843inter5));
  nor2  gate1111(.a(gate843inter5), .b(gate843inter2), .O(gate843inter6));
  inv1  gate1112(.a(N2824), .O(gate843inter7));
  inv1  gate1113(.a(N1938), .O(gate843inter8));
  nand2 gate1114(.a(gate843inter8), .b(gate843inter7), .O(gate843inter9));
  nand2 gate1115(.a(s_33), .b(gate843inter3), .O(gate843inter10));
  nor2  gate1116(.a(gate843inter10), .b(gate843inter9), .O(gate843inter11));
  nor2  gate1117(.a(gate843inter11), .b(gate843inter6), .O(gate843inter12));
  nand2 gate1118(.a(gate843inter12), .b(gate843inter1), .O(N2854));
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );

  xor2  gate3457(.a(N1985), .b(N2829), .O(gate850inter0));
  nand2 gate3458(.a(gate850inter0), .b(s_368), .O(gate850inter1));
  and2  gate3459(.a(N1985), .b(N2829), .O(gate850inter2));
  inv1  gate3460(.a(s_368), .O(gate850inter3));
  inv1  gate3461(.a(s_369), .O(gate850inter4));
  nand2 gate3462(.a(gate850inter4), .b(gate850inter3), .O(gate850inter5));
  nor2  gate3463(.a(gate850inter5), .b(gate850inter2), .O(gate850inter6));
  inv1  gate3464(.a(N2829), .O(gate850inter7));
  inv1  gate3465(.a(N1985), .O(gate850inter8));
  nand2 gate3466(.a(gate850inter8), .b(gate850inter7), .O(gate850inter9));
  nand2 gate3467(.a(s_369), .b(gate850inter3), .O(gate850inter10));
  nor2  gate3468(.a(gate850inter10), .b(gate850inter9), .O(gate850inter11));
  nor2  gate3469(.a(gate850inter11), .b(gate850inter6), .O(gate850inter12));
  nand2 gate3470(.a(gate850inter12), .b(gate850inter1), .O(N2863));

  xor2  gate2729(.a(N2857), .b(N2052), .O(gate851inter0));
  nand2 gate2730(.a(gate851inter0), .b(s_264), .O(gate851inter1));
  and2  gate2731(.a(N2857), .b(N2052), .O(gate851inter2));
  inv1  gate2732(.a(s_264), .O(gate851inter3));
  inv1  gate2733(.a(s_265), .O(gate851inter4));
  nand2 gate2734(.a(gate851inter4), .b(gate851inter3), .O(gate851inter5));
  nor2  gate2735(.a(gate851inter5), .b(gate851inter2), .O(gate851inter6));
  inv1  gate2736(.a(N2052), .O(gate851inter7));
  inv1  gate2737(.a(N2857), .O(gate851inter8));
  nand2 gate2738(.a(gate851inter8), .b(gate851inter7), .O(gate851inter9));
  nand2 gate2739(.a(s_265), .b(gate851inter3), .O(gate851inter10));
  nor2  gate2740(.a(gate851inter10), .b(gate851inter9), .O(gate851inter11));
  nor2  gate2741(.a(gate851inter11), .b(gate851inter6), .O(gate851inter12));
  nand2 gate2742(.a(gate851inter12), .b(gate851inter1), .O(N2866));

  xor2  gate3247(.a(N2858), .b(N2055), .O(gate852inter0));
  nand2 gate3248(.a(gate852inter0), .b(s_338), .O(gate852inter1));
  and2  gate3249(.a(N2858), .b(N2055), .O(gate852inter2));
  inv1  gate3250(.a(s_338), .O(gate852inter3));
  inv1  gate3251(.a(s_339), .O(gate852inter4));
  nand2 gate3252(.a(gate852inter4), .b(gate852inter3), .O(gate852inter5));
  nor2  gate3253(.a(gate852inter5), .b(gate852inter2), .O(gate852inter6));
  inv1  gate3254(.a(N2055), .O(gate852inter7));
  inv1  gate3255(.a(N2858), .O(gate852inter8));
  nand2 gate3256(.a(gate852inter8), .b(gate852inter7), .O(gate852inter9));
  nand2 gate3257(.a(s_339), .b(gate852inter3), .O(gate852inter10));
  nor2  gate3258(.a(gate852inter10), .b(gate852inter9), .O(gate852inter11));
  nor2  gate3259(.a(gate852inter11), .b(gate852inter6), .O(gate852inter12));
  nand2 gate3260(.a(gate852inter12), .b(gate852inter1), .O(N2867));
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );

  xor2  gate1245(.a(N887), .b(N2846), .O(gate858inter0));
  nand2 gate1246(.a(gate858inter0), .b(s_52), .O(gate858inter1));
  and2  gate1247(.a(N887), .b(N2846), .O(gate858inter2));
  inv1  gate1248(.a(s_52), .O(gate858inter3));
  inv1  gate1249(.a(s_53), .O(gate858inter4));
  nand2 gate1250(.a(gate858inter4), .b(gate858inter3), .O(gate858inter5));
  nor2  gate1251(.a(gate858inter5), .b(gate858inter2), .O(gate858inter6));
  inv1  gate1252(.a(N2846), .O(gate858inter7));
  inv1  gate1253(.a(N887), .O(gate858inter8));
  nand2 gate1254(.a(gate858inter8), .b(gate858inter7), .O(gate858inter9));
  nand2 gate1255(.a(s_53), .b(gate858inter3), .O(gate858inter10));
  nor2  gate1256(.a(gate858inter10), .b(gate858inter9), .O(gate858inter11));
  nor2  gate1257(.a(gate858inter11), .b(gate858inter6), .O(gate858inter12));
  nand2 gate1258(.a(gate858inter12), .b(gate858inter1), .O(N2873));
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate909(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate910(.a(gate860inter0), .b(s_4), .O(gate860inter1));
  and2  gate911(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate912(.a(s_4), .O(gate860inter3));
  inv1  gate913(.a(s_5), .O(gate860inter4));
  nand2 gate914(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate915(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate916(.a(N1933), .O(gate860inter7));
  inv1  gate917(.a(N2862), .O(gate860inter8));
  nand2 gate918(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate919(.a(s_5), .b(gate860inter3), .O(gate860inter10));
  nor2  gate920(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate921(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate922(.a(gate860inter12), .b(gate860inter1), .O(N2875));

  xor2  gate1581(.a(N2850), .b(N2866), .O(gate861inter0));
  nand2 gate1582(.a(gate861inter0), .b(s_100), .O(gate861inter1));
  and2  gate1583(.a(N2850), .b(N2866), .O(gate861inter2));
  inv1  gate1584(.a(s_100), .O(gate861inter3));
  inv1  gate1585(.a(s_101), .O(gate861inter4));
  nand2 gate1586(.a(gate861inter4), .b(gate861inter3), .O(gate861inter5));
  nor2  gate1587(.a(gate861inter5), .b(gate861inter2), .O(gate861inter6));
  inv1  gate1588(.a(N2866), .O(gate861inter7));
  inv1  gate1589(.a(N2850), .O(gate861inter8));
  nand2 gate1590(.a(gate861inter8), .b(gate861inter7), .O(gate861inter9));
  nand2 gate1591(.a(s_101), .b(gate861inter3), .O(gate861inter10));
  nor2  gate1592(.a(gate861inter10), .b(gate861inter9), .O(gate861inter11));
  nor2  gate1593(.a(gate861inter11), .b(gate861inter6), .O(gate861inter12));
  nand2 gate1594(.a(gate861inter12), .b(gate861inter1), .O(N2876));
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );

  xor2  gate2589(.a(N2852), .b(N2868), .O(gate863inter0));
  nand2 gate2590(.a(gate863inter0), .b(s_244), .O(gate863inter1));
  and2  gate2591(.a(N2852), .b(N2868), .O(gate863inter2));
  inv1  gate2592(.a(s_244), .O(gate863inter3));
  inv1  gate2593(.a(s_245), .O(gate863inter4));
  nand2 gate2594(.a(gate863inter4), .b(gate863inter3), .O(gate863inter5));
  nor2  gate2595(.a(gate863inter5), .b(gate863inter2), .O(gate863inter6));
  inv1  gate2596(.a(N2868), .O(gate863inter7));
  inv1  gate2597(.a(N2852), .O(gate863inter8));
  nand2 gate2598(.a(gate863inter8), .b(gate863inter7), .O(gate863inter9));
  nand2 gate2599(.a(s_245), .b(gate863inter3), .O(gate863inter10));
  nor2  gate2600(.a(gate863inter10), .b(gate863inter9), .O(gate863inter11));
  nor2  gate2601(.a(gate863inter11), .b(gate863inter6), .O(gate863inter12));
  nand2 gate2602(.a(gate863inter12), .b(gate863inter1), .O(N2878));

  xor2  gate2519(.a(N2853), .b(N2869), .O(gate864inter0));
  nand2 gate2520(.a(gate864inter0), .b(s_234), .O(gate864inter1));
  and2  gate2521(.a(N2853), .b(N2869), .O(gate864inter2));
  inv1  gate2522(.a(s_234), .O(gate864inter3));
  inv1  gate2523(.a(s_235), .O(gate864inter4));
  nand2 gate2524(.a(gate864inter4), .b(gate864inter3), .O(gate864inter5));
  nor2  gate2525(.a(gate864inter5), .b(gate864inter2), .O(gate864inter6));
  inv1  gate2526(.a(N2869), .O(gate864inter7));
  inv1  gate2527(.a(N2853), .O(gate864inter8));
  nand2 gate2528(.a(gate864inter8), .b(gate864inter7), .O(gate864inter9));
  nand2 gate2529(.a(s_235), .b(gate864inter3), .O(gate864inter10));
  nor2  gate2530(.a(gate864inter10), .b(gate864inter9), .O(gate864inter11));
  nor2  gate2531(.a(gate864inter11), .b(gate864inter6), .O(gate864inter12));
  nand2 gate2532(.a(gate864inter12), .b(gate864inter1), .O(N2879));

  xor2  gate2953(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate2954(.a(gate865inter0), .b(s_296), .O(gate865inter1));
  and2  gate2955(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate2956(.a(s_296), .O(gate865inter3));
  inv1  gate2957(.a(s_297), .O(gate865inter4));
  nand2 gate2958(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate2959(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate2960(.a(N2870), .O(gate865inter7));
  inv1  gate2961(.a(N2854), .O(gate865inter8));
  nand2 gate2962(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate2963(.a(s_297), .b(gate865inter3), .O(gate865inter10));
  nor2  gate2964(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate2965(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate2966(.a(gate865inter12), .b(gate865inter1), .O(N2880));
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate1679(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate1680(.a(gate874inter0), .b(s_114), .O(gate874inter1));
  and2  gate1681(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate1682(.a(s_114), .O(gate874inter3));
  inv1  gate1683(.a(s_115), .O(gate874inter4));
  nand2 gate1684(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate1685(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate1686(.a(N2871), .O(gate874inter7));
  inv1  gate1687(.a(N2881), .O(gate874inter8));
  nand2 gate1688(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate1689(.a(s_115), .b(gate874inter3), .O(gate874inter10));
  nor2  gate1690(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate1691(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate1692(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule