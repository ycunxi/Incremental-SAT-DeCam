module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate605inter0, gate605inter1, gate605inter2, gate605inter3, gate605inter4, gate605inter5, gate605inter6, gate605inter7, gate605inter8, gate605inter9, gate605inter10, gate605inter11, gate605inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate530inter0, gate530inter1, gate530inter2, gate530inter3, gate530inter4, gate530inter5, gate530inter6, gate530inter7, gate530inter8, gate530inter9, gate530inter10, gate530inter11, gate530inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate665inter0, gate665inter1, gate665inter2, gate665inter3, gate665inter4, gate665inter5, gate665inter6, gate665inter7, gate665inter8, gate665inter9, gate665inter10, gate665inter11, gate665inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate576inter0, gate576inter1, gate576inter2, gate576inter3, gate576inter4, gate576inter5, gate576inter6, gate576inter7, gate576inter8, gate576inter9, gate576inter10, gate576inter11, gate576inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate556inter0, gate556inter1, gate556inter2, gate556inter3, gate556inter4, gate556inter5, gate556inter6, gate556inter7, gate556inter8, gate556inter9, gate556inter10, gate556inter11, gate556inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate771inter0, gate771inter1, gate771inter2, gate771inter3, gate771inter4, gate771inter5, gate771inter6, gate771inter7, gate771inter8, gate771inter9, gate771inter10, gate771inter11, gate771inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate769inter0, gate769inter1, gate769inter2, gate769inter3, gate769inter4, gate769inter5, gate769inter6, gate769inter7, gate769inter8, gate769inter9, gate769inter10, gate769inter11, gate769inter12, gate572inter0, gate572inter1, gate572inter2, gate572inter3, gate572inter4, gate572inter5, gate572inter6, gate572inter7, gate572inter8, gate572inter9, gate572inter10, gate572inter11, gate572inter12, gate807inter0, gate807inter1, gate807inter2, gate807inter3, gate807inter4, gate807inter5, gate807inter6, gate807inter7, gate807inter8, gate807inter9, gate807inter10, gate807inter11, gate807inter12, gate543inter0, gate543inter1, gate543inter2, gate543inter3, gate543inter4, gate543inter5, gate543inter6, gate543inter7, gate543inter8, gate543inter9, gate543inter10, gate543inter11, gate543inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate673inter0, gate673inter1, gate673inter2, gate673inter3, gate673inter4, gate673inter5, gate673inter6, gate673inter7, gate673inter8, gate673inter9, gate673inter10, gate673inter11, gate673inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate671inter0, gate671inter1, gate671inter2, gate671inter3, gate671inter4, gate671inter5, gate671inter6, gate671inter7, gate671inter8, gate671inter9, gate671inter10, gate671inter11, gate671inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate824inter0, gate824inter1, gate824inter2, gate824inter3, gate824inter4, gate824inter5, gate824inter6, gate824inter7, gate824inter8, gate824inter9, gate824inter10, gate824inter11, gate824inter12, gate372inter0, gate372inter1, gate372inter2, gate372inter3, gate372inter4, gate372inter5, gate372inter6, gate372inter7, gate372inter8, gate372inter9, gate372inter10, gate372inter11, gate372inter12, gate305inter0, gate305inter1, gate305inter2, gate305inter3, gate305inter4, gate305inter5, gate305inter6, gate305inter7, gate305inter8, gate305inter9, gate305inter10, gate305inter11, gate305inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate315inter0, gate315inter1, gate315inter2, gate315inter3, gate315inter4, gate315inter5, gate315inter6, gate315inter7, gate315inter8, gate315inter9, gate315inter10, gate315inter11, gate315inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate676inter0, gate676inter1, gate676inter2, gate676inter3, gate676inter4, gate676inter5, gate676inter6, gate676inter7, gate676inter8, gate676inter9, gate676inter10, gate676inter11, gate676inter12, gate803inter0, gate803inter1, gate803inter2, gate803inter3, gate803inter4, gate803inter5, gate803inter6, gate803inter7, gate803inter8, gate803inter9, gate803inter10, gate803inter11, gate803inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate642inter0, gate642inter1, gate642inter2, gate642inter3, gate642inter4, gate642inter5, gate642inter6, gate642inter7, gate642inter8, gate642inter9, gate642inter10, gate642inter11, gate642inter12, gate835inter0, gate835inter1, gate835inter2, gate835inter3, gate835inter4, gate835inter5, gate835inter6, gate835inter7, gate835inter8, gate835inter9, gate835inter10, gate835inter11, gate835inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate809inter0, gate809inter1, gate809inter2, gate809inter3, gate809inter4, gate809inter5, gate809inter6, gate809inter7, gate809inter8, gate809inter9, gate809inter10, gate809inter11, gate809inter12, gate817inter0, gate817inter1, gate817inter2, gate817inter3, gate817inter4, gate817inter5, gate817inter6, gate817inter7, gate817inter8, gate817inter9, gate817inter10, gate817inter11, gate817inter12, gate822inter0, gate822inter1, gate822inter2, gate822inter3, gate822inter4, gate822inter5, gate822inter6, gate822inter7, gate822inter8, gate822inter9, gate822inter10, gate822inter11, gate822inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate819inter0, gate819inter1, gate819inter2, gate819inter3, gate819inter4, gate819inter5, gate819inter6, gate819inter7, gate819inter8, gate819inter9, gate819inter10, gate819inter11, gate819inter12, gate854inter0, gate854inter1, gate854inter2, gate854inter3, gate854inter4, gate854inter5, gate854inter6, gate854inter7, gate854inter8, gate854inter9, gate854inter10, gate854inter11, gate854inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate680inter0, gate680inter1, gate680inter2, gate680inter3, gate680inter4, gate680inter5, gate680inter6, gate680inter7, gate680inter8, gate680inter9, gate680inter10, gate680inter11, gate680inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate380inter0, gate380inter1, gate380inter2, gate380inter3, gate380inter4, gate380inter5, gate380inter6, gate380inter7, gate380inter8, gate380inter9, gate380inter10, gate380inter11, gate380inter12, gate563inter0, gate563inter1, gate563inter2, gate563inter3, gate563inter4, gate563inter5, gate563inter6, gate563inter7, gate563inter8, gate563inter9, gate563inter10, gate563inter11, gate563inter12, gate385inter0, gate385inter1, gate385inter2, gate385inter3, gate385inter4, gate385inter5, gate385inter6, gate385inter7, gate385inter8, gate385inter9, gate385inter10, gate385inter11, gate385inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate801inter0, gate801inter1, gate801inter2, gate801inter3, gate801inter4, gate801inter5, gate801inter6, gate801inter7, gate801inter8, gate801inter9, gate801inter10, gate801inter11, gate801inter12, gate518inter0, gate518inter1, gate518inter2, gate518inter3, gate518inter4, gate518inter5, gate518inter6, gate518inter7, gate518inter8, gate518inter9, gate518inter10, gate518inter11, gate518inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate343inter0, gate343inter1, gate343inter2, gate343inter3, gate343inter4, gate343inter5, gate343inter6, gate343inter7, gate343inter8, gate343inter9, gate343inter10, gate343inter11, gate343inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate351inter0, gate351inter1, gate351inter2, gate351inter3, gate351inter4, gate351inter5, gate351inter6, gate351inter7, gate351inter8, gate351inter9, gate351inter10, gate351inter11, gate351inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate750inter0, gate750inter1, gate750inter2, gate750inter3, gate750inter4, gate750inter5, gate750inter6, gate750inter7, gate750inter8, gate750inter9, gate750inter10, gate750inter11, gate750inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate621inter0, gate621inter1, gate621inter2, gate621inter3, gate621inter4, gate621inter5, gate621inter6, gate621inter7, gate621inter8, gate621inter9, gate621inter10, gate621inter11, gate621inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate349inter0, gate349inter1, gate349inter2, gate349inter3, gate349inter4, gate349inter5, gate349inter6, gate349inter7, gate349inter8, gate349inter9, gate349inter10, gate349inter11, gate349inter12, gate758inter0, gate758inter1, gate758inter2, gate758inter3, gate758inter4, gate758inter5, gate758inter6, gate758inter7, gate758inter8, gate758inter9, gate758inter10, gate758inter11, gate758inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12;



inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate1903(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate1904(.a(gate17inter0), .b(s_146), .O(gate17inter1));
  and2  gate1905(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate1906(.a(s_146), .O(gate17inter3));
  inv1  gate1907(.a(s_147), .O(gate17inter4));
  nand2 gate1908(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1909(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1910(.a(N63), .O(gate17inter7));
  inv1  gate1911(.a(N88), .O(gate17inter8));
  nand2 gate1912(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1913(.a(s_147), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1914(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1915(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1916(.a(gate17inter12), .b(gate17inter1), .O(N251));
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );

  xor2  gate937(.a(N331), .b(N306), .O(gate76inter0));
  nand2 gate938(.a(gate76inter0), .b(s_8), .O(gate76inter1));
  and2  gate939(.a(N331), .b(N306), .O(gate76inter2));
  inv1  gate940(.a(s_8), .O(gate76inter3));
  inv1  gate941(.a(s_9), .O(gate76inter4));
  nand2 gate942(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate943(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate944(.a(N306), .O(gate76inter7));
  inv1  gate945(.a(N331), .O(gate76inter8));
  nand2 gate946(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate947(.a(s_9), .b(gate76inter3), .O(gate76inter10));
  nor2  gate948(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate949(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate950(.a(gate76inter12), .b(gate76inter1), .O(N551));

  xor2  gate1273(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate1274(.a(gate77inter0), .b(s_56), .O(gate77inter1));
  and2  gate1275(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate1276(.a(s_56), .O(gate77inter3));
  inv1  gate1277(.a(s_57), .O(gate77inter4));
  nand2 gate1278(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1279(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1280(.a(N306), .O(gate77inter7));
  inv1  gate1281(.a(N331), .O(gate77inter8));
  nand2 gate1282(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1283(.a(s_57), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1284(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1285(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1286(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );

  xor2  gate1133(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate1134(.a(gate79inter0), .b(s_36), .O(gate79inter1));
  and2  gate1135(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate1136(.a(s_36), .O(gate79inter3));
  inv1  gate1137(.a(s_37), .O(gate79inter4));
  nand2 gate1138(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1139(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1140(.a(N306), .O(gate79inter7));
  inv1  gate1141(.a(N331), .O(gate79inter8));
  nand2 gate1142(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1143(.a(s_37), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1144(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1145(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1146(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate1203(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate1204(.a(gate96inter0), .b(s_46), .O(gate96inter1));
  and2  gate1205(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate1206(.a(s_46), .O(gate96inter3));
  inv1  gate1207(.a(s_47), .O(gate96inter4));
  nand2 gate1208(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1209(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1210(.a(N326), .O(gate96inter7));
  inv1  gate1211(.a(N277), .O(gate96inter8));
  nand2 gate1212(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1213(.a(s_47), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1214(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1215(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1216(.a(gate96inter12), .b(gate96inter1), .O(N601));

  xor2  gate1679(.a(N280), .b(N326), .O(gate97inter0));
  nand2 gate1680(.a(gate97inter0), .b(s_114), .O(gate97inter1));
  and2  gate1681(.a(N280), .b(N326), .O(gate97inter2));
  inv1  gate1682(.a(s_114), .O(gate97inter3));
  inv1  gate1683(.a(s_115), .O(gate97inter4));
  nand2 gate1684(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1685(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1686(.a(N326), .O(gate97inter7));
  inv1  gate1687(.a(N280), .O(gate97inter8));
  nand2 gate1688(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1689(.a(s_115), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1690(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1691(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1692(.a(gate97inter12), .b(gate97inter1), .O(N602));
nand2 gate98( .a(N260), .b(N72), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );

  xor2  gate993(.a(N300), .b(N256), .O(gate100inter0));
  nand2 gate994(.a(gate100inter0), .b(s_16), .O(gate100inter1));
  and2  gate995(.a(N300), .b(N256), .O(gate100inter2));
  inv1  gate996(.a(s_16), .O(gate100inter3));
  inv1  gate997(.a(s_17), .O(gate100inter4));
  nand2 gate998(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate999(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1000(.a(N256), .O(gate100inter7));
  inv1  gate1001(.a(N300), .O(gate100inter8));
  nand2 gate1002(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1003(.a(s_17), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1004(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1005(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1006(.a(gate100inter12), .b(gate100inter1), .O(N612));
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );

  xor2  gate1973(.a(N608), .b(N56), .O(gate163inter0));
  nand2 gate1974(.a(gate163inter0), .b(s_156), .O(gate163inter1));
  and2  gate1975(.a(N608), .b(N56), .O(gate163inter2));
  inv1  gate1976(.a(s_156), .O(gate163inter3));
  inv1  gate1977(.a(s_157), .O(gate163inter4));
  nand2 gate1978(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1979(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1980(.a(N56), .O(gate163inter7));
  inv1  gate1981(.a(N608), .O(gate163inter8));
  nand2 gate1982(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1983(.a(s_157), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1984(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1985(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1986(.a(gate163inter12), .b(gate163inter1), .O(N910));
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );

  xor2  gate1623(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate1624(.a(gate236inter0), .b(s_106), .O(gate236inter1));
  and2  gate1625(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate1626(.a(s_106), .O(gate236inter3));
  inv1  gate1627(.a(s_107), .O(gate236inter4));
  nand2 gate1628(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1629(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1630(.a(N622), .O(gate236inter7));
  inv1  gate1631(.a(N891), .O(gate236inter8));
  nand2 gate1632(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1633(.a(s_107), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1634(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1635(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1636(.a(gate236inter12), .b(gate236inter1), .O(N1064));
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );

  xor2  gate951(.a(N989), .b(N718), .O(gate240inter0));
  nand2 gate952(.a(gate240inter0), .b(s_10), .O(gate240inter1));
  and2  gate953(.a(N989), .b(N718), .O(gate240inter2));
  inv1  gate954(.a(s_10), .O(gate240inter3));
  inv1  gate955(.a(s_11), .O(gate240inter4));
  nand2 gate956(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate957(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate958(.a(N718), .O(gate240inter7));
  inv1  gate959(.a(N989), .O(gate240inter8));
  nand2 gate960(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate961(.a(s_11), .b(gate240inter3), .O(gate240inter10));
  nor2  gate962(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate963(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate964(.a(gate240inter12), .b(gate240inter1), .O(N1120));

  xor2  gate1105(.a(N991), .b(N727), .O(gate241inter0));
  nand2 gate1106(.a(gate241inter0), .b(s_32), .O(gate241inter1));
  and2  gate1107(.a(N991), .b(N727), .O(gate241inter2));
  inv1  gate1108(.a(s_32), .O(gate241inter3));
  inv1  gate1109(.a(s_33), .O(gate241inter4));
  nand2 gate1110(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1111(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1112(.a(N727), .O(gate241inter7));
  inv1  gate1113(.a(N991), .O(gate241inter8));
  nand2 gate1114(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1115(.a(s_33), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1116(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1117(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1118(.a(gate241inter12), .b(gate241inter1), .O(N1121));
nand2 gate242( .a(N724), .b(N992), .O(N1122) );

  xor2  gate1063(.a(N1002), .b(N739), .O(gate243inter0));
  nand2 gate1064(.a(gate243inter0), .b(s_26), .O(gate243inter1));
  and2  gate1065(.a(N1002), .b(N739), .O(gate243inter2));
  inv1  gate1066(.a(s_26), .O(gate243inter3));
  inv1  gate1067(.a(s_27), .O(gate243inter4));
  nand2 gate1068(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1069(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1070(.a(N739), .O(gate243inter7));
  inv1  gate1071(.a(N1002), .O(gate243inter8));
  nand2 gate1072(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1073(.a(s_27), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1074(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1075(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1076(.a(gate243inter12), .b(gate243inter1), .O(N1128));

  xor2  gate1525(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate1526(.a(gate244inter0), .b(s_92), .O(gate244inter1));
  and2  gate1527(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate1528(.a(s_92), .O(gate244inter3));
  inv1  gate1529(.a(s_93), .O(gate244inter4));
  nand2 gate1530(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1531(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1532(.a(N736), .O(gate244inter7));
  inv1  gate1533(.a(N1003), .O(gate244inter8));
  nand2 gate1534(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1535(.a(s_93), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1536(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1537(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1538(.a(gate244inter12), .b(gate244inter1), .O(N1129));

  xor2  gate1189(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate1190(.a(gate245inter0), .b(s_44), .O(gate245inter1));
  and2  gate1191(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate1192(.a(s_44), .O(gate245inter3));
  inv1  gate1193(.a(s_45), .O(gate245inter4));
  nand2 gate1194(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1195(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1196(.a(N745), .O(gate245inter7));
  inv1  gate1197(.a(N1005), .O(gate245inter8));
  nand2 gate1198(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1199(.a(s_45), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1200(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1201(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1202(.a(gate245inter12), .b(gate245inter1), .O(N1130));
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );

  xor2  gate1721(.a(N1009), .b(N748), .O(gate248inter0));
  nand2 gate1722(.a(gate248inter0), .b(s_120), .O(gate248inter1));
  and2  gate1723(.a(N1009), .b(N748), .O(gate248inter2));
  inv1  gate1724(.a(s_120), .O(gate248inter3));
  inv1  gate1725(.a(s_121), .O(gate248inter4));
  nand2 gate1726(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1727(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1728(.a(N748), .O(gate248inter7));
  inv1  gate1729(.a(N1009), .O(gate248inter8));
  nand2 gate1730(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1731(.a(s_121), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1732(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1733(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1734(.a(gate248inter12), .b(gate248inter1), .O(N1133));
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );

  xor2  gate1217(.a(N1068), .b(N1067), .O(gate263inter0));
  nand2 gate1218(.a(gate263inter0), .b(s_48), .O(gate263inter1));
  and2  gate1219(.a(N1068), .b(N1067), .O(gate263inter2));
  inv1  gate1220(.a(s_48), .O(gate263inter3));
  inv1  gate1221(.a(s_49), .O(gate263inter4));
  nand2 gate1222(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1223(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1224(.a(N1067), .O(gate263inter7));
  inv1  gate1225(.a(N1068), .O(gate263inter8));
  nand2 gate1226(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1227(.a(s_49), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1228(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1229(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1230(.a(gate263inter12), .b(gate263inter1), .O(N1162));
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate1763(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate1764(.a(gate277inter0), .b(s_126), .O(gate277inter1));
  and2  gate1765(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate1766(.a(s_126), .O(gate277inter3));
  inv1  gate1767(.a(s_127), .O(gate277inter4));
  nand2 gate1768(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1769(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1770(.a(N1019), .O(gate277inter7));
  inv1  gate1771(.a(N950), .O(gate277inter8));
  nand2 gate1772(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1773(.a(s_127), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1774(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1775(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1776(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );

  xor2  gate1385(.a(N958), .b(N1025), .O(gate281inter0));
  nand2 gate1386(.a(gate281inter0), .b(s_72), .O(gate281inter1));
  and2  gate1387(.a(N958), .b(N1025), .O(gate281inter2));
  inv1  gate1388(.a(s_72), .O(gate281inter3));
  inv1  gate1389(.a(s_73), .O(gate281inter4));
  nand2 gate1390(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1391(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1392(.a(N1025), .O(gate281inter7));
  inv1  gate1393(.a(N958), .O(gate281inter8));
  nand2 gate1394(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1395(.a(s_73), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1396(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1397(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1398(.a(gate281inter12), .b(gate281inter1), .O(N1216));
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );

  xor2  gate1875(.a(N972), .b(N1037), .O(gate289inter0));
  nand2 gate1876(.a(gate289inter0), .b(s_142), .O(gate289inter1));
  and2  gate1877(.a(N972), .b(N1037), .O(gate289inter2));
  inv1  gate1878(.a(s_142), .O(gate289inter3));
  inv1  gate1879(.a(s_143), .O(gate289inter4));
  nand2 gate1880(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1881(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1882(.a(N1037), .O(gate289inter7));
  inv1  gate1883(.a(N972), .O(gate289inter8));
  nand2 gate1884(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1885(.a(s_143), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1886(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1887(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1888(.a(gate289inter12), .b(gate289inter1), .O(N1224));
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );

  xor2  gate1357(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate1358(.a(gate297inter0), .b(s_68), .O(gate297inter1));
  and2  gate1359(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate1360(.a(s_68), .O(gate297inter3));
  inv1  gate1361(.a(s_69), .O(gate297inter4));
  nand2 gate1362(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate1363(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate1364(.a(N1119), .O(gate297inter7));
  inv1  gate1365(.a(N1120), .O(gate297inter8));
  nand2 gate1366(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate1367(.a(s_69), .b(gate297inter3), .O(gate297inter10));
  nor2  gate1368(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate1369(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate1370(.a(gate297inter12), .b(gate297inter1), .O(N1232));

  xor2  gate1147(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate1148(.a(gate298inter0), .b(s_38), .O(gate298inter1));
  and2  gate1149(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate1150(.a(s_38), .O(gate298inter3));
  inv1  gate1151(.a(s_39), .O(gate298inter4));
  nand2 gate1152(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate1153(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate1154(.a(N1121), .O(gate298inter7));
  inv1  gate1155(.a(N1122), .O(gate298inter8));
  nand2 gate1156(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate1157(.a(s_39), .b(gate298inter3), .O(gate298inter10));
  nor2  gate1158(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate1159(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate1160(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );

  xor2  gate1455(.a(N1131), .b(N1130), .O(gate305inter0));
  nand2 gate1456(.a(gate305inter0), .b(s_82), .O(gate305inter1));
  and2  gate1457(.a(N1131), .b(N1130), .O(gate305inter2));
  inv1  gate1458(.a(s_82), .O(gate305inter3));
  inv1  gate1459(.a(s_83), .O(gate305inter4));
  nand2 gate1460(.a(gate305inter4), .b(gate305inter3), .O(gate305inter5));
  nor2  gate1461(.a(gate305inter5), .b(gate305inter2), .O(gate305inter6));
  inv1  gate1462(.a(N1130), .O(gate305inter7));
  inv1  gate1463(.a(N1131), .O(gate305inter8));
  nand2 gate1464(.a(gate305inter8), .b(gate305inter7), .O(gate305inter9));
  nand2 gate1465(.a(s_83), .b(gate305inter3), .O(gate305inter10));
  nor2  gate1466(.a(gate305inter10), .b(gate305inter9), .O(gate305inter11));
  nor2  gate1467(.a(gate305inter11), .b(gate305inter6), .O(gate305inter12));
  nand2 gate1468(.a(gate305inter12), .b(gate305inter1), .O(N1246));
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate923(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate924(.a(gate312inter0), .b(s_6), .O(gate312inter1));
  and2  gate925(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate926(.a(s_6), .O(gate312inter3));
  inv1  gate927(.a(s_7), .O(gate312inter4));
  nand2 gate928(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate929(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate930(.a(N631), .O(gate312inter7));
  inv1  gate931(.a(N1159), .O(gate312inter8));
  nand2 gate932(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate933(.a(s_7), .b(gate312inter3), .O(gate312inter10));
  nor2  gate934(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate935(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate936(.a(gate312inter12), .b(gate312inter1), .O(N1267));
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );

  xor2  gate1511(.a(N1207), .b(N691), .O(gate314inter0));
  nand2 gate1512(.a(gate314inter0), .b(s_90), .O(gate314inter1));
  and2  gate1513(.a(N1207), .b(N691), .O(gate314inter2));
  inv1  gate1514(.a(s_90), .O(gate314inter3));
  inv1  gate1515(.a(s_91), .O(gate314inter4));
  nand2 gate1516(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate1517(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate1518(.a(N691), .O(gate314inter7));
  inv1  gate1519(.a(N1207), .O(gate314inter8));
  nand2 gate1520(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate1521(.a(s_91), .b(gate314inter3), .O(gate314inter10));
  nor2  gate1522(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate1523(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate1524(.a(gate314inter12), .b(gate314inter1), .O(N1310));

  xor2  gate1483(.a(N1209), .b(N694), .O(gate315inter0));
  nand2 gate1484(.a(gate315inter0), .b(s_86), .O(gate315inter1));
  and2  gate1485(.a(N1209), .b(N694), .O(gate315inter2));
  inv1  gate1486(.a(s_86), .O(gate315inter3));
  inv1  gate1487(.a(s_87), .O(gate315inter4));
  nand2 gate1488(.a(gate315inter4), .b(gate315inter3), .O(gate315inter5));
  nor2  gate1489(.a(gate315inter5), .b(gate315inter2), .O(gate315inter6));
  inv1  gate1490(.a(N694), .O(gate315inter7));
  inv1  gate1491(.a(N1209), .O(gate315inter8));
  nand2 gate1492(.a(gate315inter8), .b(gate315inter7), .O(gate315inter9));
  nand2 gate1493(.a(s_87), .b(gate315inter3), .O(gate315inter10));
  nor2  gate1494(.a(gate315inter10), .b(gate315inter9), .O(gate315inter11));
  nor2  gate1495(.a(gate315inter11), .b(gate315inter6), .O(gate315inter12));
  nand2 gate1496(.a(gate315inter12), .b(gate315inter1), .O(N1311));

  xor2  gate1231(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate1232(.a(gate316inter0), .b(s_50), .O(gate316inter1));
  and2  gate1233(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate1234(.a(s_50), .O(gate316inter3));
  inv1  gate1235(.a(s_51), .O(gate316inter4));
  nand2 gate1236(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate1237(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate1238(.a(N697), .O(gate316inter7));
  inv1  gate1239(.a(N1211), .O(gate316inter8));
  nand2 gate1240(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate1241(.a(s_51), .b(gate316inter3), .O(gate316inter10));
  nor2  gate1242(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate1243(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate1244(.a(gate316inter12), .b(gate316inter1), .O(N1312));

  xor2  gate2253(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate2254(.a(gate317inter0), .b(s_196), .O(gate317inter1));
  and2  gate2255(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate2256(.a(s_196), .O(gate317inter3));
  inv1  gate2257(.a(s_197), .O(gate317inter4));
  nand2 gate2258(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate2259(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate2260(.a(N700), .O(gate317inter7));
  inv1  gate2261(.a(N1213), .O(gate317inter8));
  nand2 gate2262(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate2263(.a(s_197), .b(gate317inter3), .O(gate317inter10));
  nor2  gate2264(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate2265(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate2266(.a(gate317inter12), .b(gate317inter1), .O(N1313));
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );

  xor2  gate2141(.a(N1228), .b(N715), .O(gate322inter0));
  nand2 gate2142(.a(gate322inter0), .b(s_180), .O(gate322inter1));
  and2  gate2143(.a(N1228), .b(N715), .O(gate322inter2));
  inv1  gate2144(.a(s_180), .O(gate322inter3));
  inv1  gate2145(.a(s_181), .O(gate322inter4));
  nand2 gate2146(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate2147(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate2148(.a(N715), .O(gate322inter7));
  inv1  gate2149(.a(N1228), .O(gate322inter8));
  nand2 gate2150(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate2151(.a(s_181), .b(gate322inter3), .O(gate322inter10));
  nor2  gate2152(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate2153(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate2154(.a(gate322inter12), .b(gate322inter1), .O(N1318));
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );

  xor2  gate1469(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate1470(.a(gate326inter0), .b(s_84), .O(gate326inter1));
  and2  gate1471(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate1472(.a(s_84), .O(gate326inter3));
  inv1  gate1473(.a(s_85), .O(gate326inter4));
  nand2 gate1474(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate1475(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate1476(.a(N733), .O(gate326inter7));
  inv1  gate1477(.a(N1241), .O(gate326inter8));
  nand2 gate1478(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate1479(.a(s_85), .b(gate326inter3), .O(gate326inter10));
  nor2  gate1480(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate1481(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate1482(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );

  xor2  gate2015(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate2016(.a(gate342inter0), .b(s_162), .O(gate342inter1));
  and2  gate2017(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate2018(.a(s_162), .O(gate342inter3));
  inv1  gate2019(.a(s_163), .O(gate342inter4));
  nand2 gate2020(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate2021(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate2022(.a(N1316), .O(gate342inter7));
  inv1  gate2023(.a(N1224), .O(gate342inter8));
  nand2 gate2024(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate2025(.a(s_163), .b(gate342inter3), .O(gate342inter10));
  nor2  gate2026(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate2027(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate2028(.a(gate342inter12), .b(gate342inter1), .O(N1373));

  xor2  gate2071(.a(N1226), .b(N1317), .O(gate343inter0));
  nand2 gate2072(.a(gate343inter0), .b(s_170), .O(gate343inter1));
  and2  gate2073(.a(N1226), .b(N1317), .O(gate343inter2));
  inv1  gate2074(.a(s_170), .O(gate343inter3));
  inv1  gate2075(.a(s_171), .O(gate343inter4));
  nand2 gate2076(.a(gate343inter4), .b(gate343inter3), .O(gate343inter5));
  nor2  gate2077(.a(gate343inter5), .b(gate343inter2), .O(gate343inter6));
  inv1  gate2078(.a(N1317), .O(gate343inter7));
  inv1  gate2079(.a(N1226), .O(gate343inter8));
  nand2 gate2080(.a(gate343inter8), .b(gate343inter7), .O(gate343inter9));
  nand2 gate2081(.a(s_171), .b(gate343inter3), .O(gate343inter10));
  nor2  gate2082(.a(gate343inter10), .b(gate343inter9), .O(gate343inter11));
  nor2  gate2083(.a(gate343inter11), .b(gate343inter6), .O(gate343inter12));
  nand2 gate2084(.a(gate343inter12), .b(gate343inter1), .O(N1376));
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );

  xor2  gate2183(.a(N993), .b(N1235), .O(gate349inter0));
  nand2 gate2184(.a(gate349inter0), .b(s_186), .O(gate349inter1));
  and2  gate2185(.a(N993), .b(N1235), .O(gate349inter2));
  inv1  gate2186(.a(s_186), .O(gate349inter3));
  inv1  gate2187(.a(s_187), .O(gate349inter4));
  nand2 gate2188(.a(gate349inter4), .b(gate349inter3), .O(gate349inter5));
  nor2  gate2189(.a(gate349inter5), .b(gate349inter2), .O(gate349inter6));
  inv1  gate2190(.a(N1235), .O(gate349inter7));
  inv1  gate2191(.a(N993), .O(gate349inter8));
  nand2 gate2192(.a(gate349inter8), .b(gate349inter7), .O(gate349inter9));
  nand2 gate2193(.a(s_187), .b(gate349inter3), .O(gate349inter10));
  nor2  gate2194(.a(gate349inter10), .b(gate349inter9), .O(gate349inter11));
  nor2  gate2195(.a(gate349inter11), .b(gate349inter6), .O(gate349inter12));
  nand2 gate2196(.a(gate349inter12), .b(gate349inter1), .O(N1389));
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );

  xor2  gate2099(.a(N1242), .b(N1328), .O(gate351inter0));
  nand2 gate2100(.a(gate351inter0), .b(s_174), .O(gate351inter1));
  and2  gate2101(.a(N1242), .b(N1328), .O(gate351inter2));
  inv1  gate2102(.a(s_174), .O(gate351inter3));
  inv1  gate2103(.a(s_175), .O(gate351inter4));
  nand2 gate2104(.a(gate351inter4), .b(gate351inter3), .O(gate351inter5));
  nor2  gate2105(.a(gate351inter5), .b(gate351inter2), .O(gate351inter6));
  inv1  gate2106(.a(N1328), .O(gate351inter7));
  inv1  gate2107(.a(N1242), .O(gate351inter8));
  nand2 gate2108(.a(gate351inter8), .b(gate351inter7), .O(gate351inter9));
  nand2 gate2109(.a(s_175), .b(gate351inter3), .O(gate351inter10));
  nor2  gate2110(.a(gate351inter10), .b(gate351inter9), .O(gate351inter11));
  nor2  gate2111(.a(gate351inter11), .b(gate351inter6), .O(gate351inter12));
  nand2 gate2112(.a(gate351inter12), .b(gate351inter1), .O(N1393));
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );

  xor2  gate1441(.a(N1152), .b(N1361), .O(gate372inter0));
  nand2 gate1442(.a(gate372inter0), .b(s_80), .O(gate372inter1));
  and2  gate1443(.a(N1152), .b(N1361), .O(gate372inter2));
  inv1  gate1444(.a(s_80), .O(gate372inter3));
  inv1  gate1445(.a(s_81), .O(gate372inter4));
  nand2 gate1446(.a(gate372inter4), .b(gate372inter3), .O(gate372inter5));
  nor2  gate1447(.a(gate372inter5), .b(gate372inter2), .O(gate372inter6));
  inv1  gate1448(.a(N1361), .O(gate372inter7));
  inv1  gate1449(.a(N1152), .O(gate372inter8));
  nand2 gate1450(.a(gate372inter8), .b(gate372inter7), .O(gate372inter9));
  nand2 gate1451(.a(s_81), .b(gate372inter3), .O(gate372inter10));
  nor2  gate1452(.a(gate372inter10), .b(gate372inter9), .O(gate372inter11));
  nor2  gate1453(.a(gate372inter11), .b(gate372inter6), .O(gate372inter12));
  nand2 gate1454(.a(gate372inter12), .b(gate372inter1), .O(N1451));
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate1889(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate1890(.a(gate376inter0), .b(s_144), .O(gate376inter1));
  and2  gate1891(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate1892(.a(s_144), .O(gate376inter3));
  inv1  gate1893(.a(s_145), .O(gate376inter4));
  nand2 gate1894(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate1895(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate1896(.a(N1364), .O(gate376inter7));
  inv1  gate1897(.a(N1154), .O(gate376inter8));
  nand2 gate1898(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate1899(.a(s_145), .b(gate376inter3), .O(gate376inter10));
  nor2  gate1900(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate1901(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate1902(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );

  xor2  gate1917(.a(N1157), .b(N1379), .O(gate380inter0));
  nand2 gate1918(.a(gate380inter0), .b(s_148), .O(gate380inter1));
  and2  gate1919(.a(N1157), .b(N1379), .O(gate380inter2));
  inv1  gate1920(.a(s_148), .O(gate380inter3));
  inv1  gate1921(.a(s_149), .O(gate380inter4));
  nand2 gate1922(.a(gate380inter4), .b(gate380inter3), .O(gate380inter5));
  nor2  gate1923(.a(gate380inter5), .b(gate380inter2), .O(gate380inter6));
  inv1  gate1924(.a(N1379), .O(gate380inter7));
  inv1  gate1925(.a(N1157), .O(gate380inter8));
  nand2 gate1926(.a(gate380inter8), .b(gate380inter7), .O(gate380inter9));
  nand2 gate1927(.a(s_149), .b(gate380inter3), .O(gate380inter10));
  nor2  gate1928(.a(gate380inter10), .b(gate380inter9), .O(gate380inter11));
  nor2  gate1929(.a(gate380inter11), .b(gate380inter6), .O(gate380inter12));
  nand2 gate1930(.a(gate380inter12), .b(gate380inter1), .O(N1459));
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate1581(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate1582(.a(gate383inter0), .b(s_100), .O(gate383inter1));
  and2  gate1583(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate1584(.a(s_100), .O(gate383inter3));
  inv1  gate1585(.a(s_101), .O(gate383inter4));
  nand2 gate1586(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate1587(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate1588(.a(N1393), .O(gate383inter7));
  inv1  gate1589(.a(N1161), .O(gate383inter8));
  nand2 gate1590(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate1591(.a(s_101), .b(gate383inter3), .O(gate383inter10));
  nor2  gate1592(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate1593(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate1594(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );

  xor2  gate1945(.a(N1412), .b(N1345), .O(gate385inter0));
  nand2 gate1946(.a(gate385inter0), .b(s_152), .O(gate385inter1));
  and2  gate1947(.a(N1412), .b(N1345), .O(gate385inter2));
  inv1  gate1948(.a(s_152), .O(gate385inter3));
  inv1  gate1949(.a(s_153), .O(gate385inter4));
  nand2 gate1950(.a(gate385inter4), .b(gate385inter3), .O(gate385inter5));
  nor2  gate1951(.a(gate385inter5), .b(gate385inter2), .O(gate385inter6));
  inv1  gate1952(.a(N1345), .O(gate385inter7));
  inv1  gate1953(.a(N1412), .O(gate385inter8));
  nand2 gate1954(.a(gate385inter8), .b(gate385inter7), .O(gate385inter9));
  nand2 gate1955(.a(s_153), .b(gate385inter3), .O(gate385inter10));
  nor2  gate1956(.a(gate385inter10), .b(gate385inter9), .O(gate385inter11));
  nor2  gate1957(.a(gate385inter11), .b(gate385inter6), .O(gate385inter12));
  nand2 gate1958(.a(gate385inter12), .b(gate385inter1), .O(N1464));
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );

  xor2  gate1693(.a(N1444), .b(N939), .O(gate396inter0));
  nand2 gate1694(.a(gate396inter0), .b(s_116), .O(gate396inter1));
  and2  gate1695(.a(N1444), .b(N939), .O(gate396inter2));
  inv1  gate1696(.a(s_116), .O(gate396inter3));
  inv1  gate1697(.a(s_117), .O(gate396inter4));
  nand2 gate1698(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1699(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1700(.a(N939), .O(gate396inter7));
  inv1  gate1701(.a(N1444), .O(gate396inter8));
  nand2 gate1702(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1703(.a(s_117), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1704(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1705(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1706(.a(gate396inter12), .b(gate396inter1), .O(N1487));

  xor2  gate1007(.a(N1446), .b(N935), .O(gate397inter0));
  nand2 gate1008(.a(gate397inter0), .b(s_18), .O(gate397inter1));
  and2  gate1009(.a(N1446), .b(N935), .O(gate397inter2));
  inv1  gate1010(.a(s_18), .O(gate397inter3));
  inv1  gate1011(.a(s_19), .O(gate397inter4));
  nand2 gate1012(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1013(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1014(.a(N935), .O(gate397inter7));
  inv1  gate1015(.a(N1446), .O(gate397inter8));
  nand2 gate1016(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1017(.a(s_19), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1018(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1019(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1020(.a(gate397inter12), .b(gate397inter1), .O(N1488));

  xor2  gate2169(.a(N1448), .b(N943), .O(gate398inter0));
  nand2 gate2170(.a(gate398inter0), .b(s_184), .O(gate398inter1));
  and2  gate2171(.a(N1448), .b(N943), .O(gate398inter2));
  inv1  gate2172(.a(s_184), .O(gate398inter3));
  inv1  gate2173(.a(s_185), .O(gate398inter4));
  nand2 gate2174(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2175(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2176(.a(N943), .O(gate398inter7));
  inv1  gate2177(.a(N1448), .O(gate398inter8));
  nand2 gate2178(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2179(.a(s_185), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2180(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2181(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2182(.a(gate398inter12), .b(gate398inter1), .O(N1489));
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );

  xor2  gate1497(.a(N1456), .b(N951), .O(gate403inter0));
  nand2 gate1498(.a(gate403inter0), .b(s_88), .O(gate403inter1));
  and2  gate1499(.a(N1456), .b(N951), .O(gate403inter2));
  inv1  gate1500(.a(s_88), .O(gate403inter3));
  inv1  gate1501(.a(s_89), .O(gate403inter4));
  nand2 gate1502(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1503(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1504(.a(N951), .O(gate403inter7));
  inv1  gate1505(.a(N1456), .O(gate403inter8));
  nand2 gate1506(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1507(.a(s_89), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1508(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1509(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1510(.a(gate403inter12), .b(gate403inter1), .O(N1494));

  xor2  gate1959(.a(N1458), .b(N969), .O(gate404inter0));
  nand2 gate1960(.a(gate404inter0), .b(s_154), .O(gate404inter1));
  and2  gate1961(.a(N1458), .b(N969), .O(gate404inter2));
  inv1  gate1962(.a(s_154), .O(gate404inter3));
  inv1  gate1963(.a(s_155), .O(gate404inter4));
  nand2 gate1964(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1965(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1966(.a(N969), .O(gate404inter7));
  inv1  gate1967(.a(N1458), .O(gate404inter8));
  nand2 gate1968(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1969(.a(s_155), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1970(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1971(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1972(.a(gate404inter12), .b(gate404inter1), .O(N1495));
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );

  xor2  gate1035(.a(N1487), .b(N1443), .O(gate412inter0));
  nand2 gate1036(.a(gate412inter0), .b(s_22), .O(gate412inter1));
  and2  gate1037(.a(N1487), .b(N1443), .O(gate412inter2));
  inv1  gate1038(.a(s_22), .O(gate412inter3));
  inv1  gate1039(.a(s_23), .O(gate412inter4));
  nand2 gate1040(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1041(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1042(.a(N1443), .O(gate412inter7));
  inv1  gate1043(.a(N1487), .O(gate412inter8));
  nand2 gate1044(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1045(.a(s_23), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1046(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1047(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1048(.a(gate412inter12), .b(gate412inter1), .O(N1513));

  xor2  gate2239(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate2240(.a(gate413inter0), .b(s_194), .O(gate413inter1));
  and2  gate2241(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate2242(.a(s_194), .O(gate413inter3));
  inv1  gate2243(.a(s_195), .O(gate413inter4));
  nand2 gate2244(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2245(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2246(.a(N1445), .O(gate413inter7));
  inv1  gate2247(.a(N1488), .O(gate413inter8));
  nand2 gate2248(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2249(.a(s_195), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2250(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2251(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2252(.a(gate413inter12), .b(gate413inter1), .O(N1514));
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );

  xor2  gate1861(.a(N1500), .b(N1469), .O(gate426inter0));
  nand2 gate1862(.a(gate426inter0), .b(s_140), .O(gate426inter1));
  and2  gate1863(.a(N1500), .b(N1469), .O(gate426inter2));
  inv1  gate1864(.a(s_140), .O(gate426inter3));
  inv1  gate1865(.a(s_141), .O(gate426inter4));
  nand2 gate1866(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1867(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1868(.a(N1469), .O(gate426inter7));
  inv1  gate1869(.a(N1500), .O(gate426inter8));
  nand2 gate1870(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1871(.a(s_141), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1872(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1873(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1874(.a(gate426inter12), .b(gate426inter1), .O(N1537));

  xor2  gate1567(.a(N1504), .b(N1476), .O(gate427inter0));
  nand2 gate1568(.a(gate427inter0), .b(s_98), .O(gate427inter1));
  and2  gate1569(.a(N1504), .b(N1476), .O(gate427inter2));
  inv1  gate1570(.a(s_98), .O(gate427inter3));
  inv1  gate1571(.a(s_99), .O(gate427inter4));
  nand2 gate1572(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1573(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1574(.a(N1476), .O(gate427inter7));
  inv1  gate1575(.a(N1504), .O(gate427inter8));
  nand2 gate1576(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1577(.a(s_99), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1578(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1579(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1580(.a(gate427inter12), .b(gate427inter1), .O(N1540));
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );

  xor2  gate2113(.a(N893), .b(N1596), .O(gate462inter0));
  nand2 gate2114(.a(gate462inter0), .b(s_176), .O(gate462inter1));
  and2  gate2115(.a(N893), .b(N1596), .O(gate462inter2));
  inv1  gate2116(.a(s_176), .O(gate462inter3));
  inv1  gate2117(.a(s_177), .O(gate462inter4));
  nand2 gate2118(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2119(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2120(.a(N1596), .O(gate462inter7));
  inv1  gate2121(.a(N893), .O(gate462inter8));
  nand2 gate2122(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2123(.a(s_177), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2124(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2125(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2126(.a(gate462inter12), .b(gate462inter1), .O(N1671));
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );

  xor2  gate1777(.a(N1219), .b(N1609), .O(gate468inter0));
  nand2 gate1778(.a(gate468inter0), .b(s_128), .O(gate468inter1));
  and2  gate1779(.a(N1219), .b(N1609), .O(gate468inter2));
  inv1  gate1780(.a(s_128), .O(gate468inter3));
  inv1  gate1781(.a(s_129), .O(gate468inter4));
  nand2 gate1782(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1783(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1784(.a(N1609), .O(gate468inter7));
  inv1  gate1785(.a(N1219), .O(gate468inter8));
  nand2 gate1786(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1787(.a(s_129), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1788(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1789(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1790(.a(gate468inter12), .b(gate468inter1), .O(N1680));
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );

  xor2  gate1175(.a(N1636), .b(N1594), .O(gate472inter0));
  nand2 gate1176(.a(gate472inter0), .b(s_42), .O(gate472inter1));
  and2  gate1177(.a(N1636), .b(N1594), .O(gate472inter2));
  inv1  gate1178(.a(s_42), .O(gate472inter3));
  inv1  gate1179(.a(s_43), .O(gate472inter4));
  nand2 gate1180(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1181(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1182(.a(N1594), .O(gate472inter7));
  inv1  gate1183(.a(N1636), .O(gate472inter8));
  nand2 gate1184(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1185(.a(s_43), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1186(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1187(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1188(.a(gate472inter12), .b(gate472inter1), .O(N1685));
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );

  xor2  gate909(.a(N1672), .b(N643), .O(gate476inter0));
  nand2 gate910(.a(gate476inter0), .b(s_4), .O(gate476inter1));
  and2  gate911(.a(N1672), .b(N643), .O(gate476inter2));
  inv1  gate912(.a(s_4), .O(gate476inter3));
  inv1  gate913(.a(s_5), .O(gate476inter4));
  nand2 gate914(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate915(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate916(.a(N643), .O(gate476inter7));
  inv1  gate917(.a(N1672), .O(gate476inter8));
  nand2 gate918(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate919(.a(s_5), .b(gate476inter3), .O(gate476inter10));
  nor2  gate920(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate921(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate922(.a(gate476inter12), .b(gate476inter1), .O(N1706));
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );

  xor2  gate1077(.a(N1677), .b(N1651), .O(gate480inter0));
  nand2 gate1078(.a(gate480inter0), .b(s_28), .O(gate480inter1));
  and2  gate1079(.a(N1677), .b(N1651), .O(gate480inter2));
  inv1  gate1080(.a(s_28), .O(gate480inter3));
  inv1  gate1081(.a(s_29), .O(gate480inter4));
  nand2 gate1082(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1083(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1084(.a(N1651), .O(gate480inter7));
  inv1  gate1085(.a(N1677), .O(gate480inter8));
  nand2 gate1086(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1087(.a(s_29), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1088(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1089(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1090(.a(gate480inter12), .b(gate480inter1), .O(N1710));
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );

  xor2  gate2267(.a(N1681), .b(N1031), .O(gate483inter0));
  nand2 gate2268(.a(gate483inter0), .b(s_198), .O(gate483inter1));
  and2  gate2269(.a(N1681), .b(N1031), .O(gate483inter2));
  inv1  gate2270(.a(s_198), .O(gate483inter3));
  inv1  gate2271(.a(s_199), .O(gate483inter4));
  nand2 gate2272(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2273(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2274(.a(N1031), .O(gate483inter7));
  inv1  gate2275(.a(N1681), .O(gate483inter8));
  nand2 gate2276(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2277(.a(s_199), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2278(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2279(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2280(.a(gate483inter12), .b(gate483inter1), .O(N1713));
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );

  xor2  gate965(.a(N1711), .b(N1603), .O(gate498inter0));
  nand2 gate966(.a(gate498inter0), .b(s_12), .O(gate498inter1));
  and2  gate967(.a(N1711), .b(N1603), .O(gate498inter2));
  inv1  gate968(.a(s_12), .O(gate498inter3));
  inv1  gate969(.a(s_13), .O(gate498inter4));
  nand2 gate970(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate971(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate972(.a(N1603), .O(gate498inter7));
  inv1  gate973(.a(N1711), .O(gate498inter8));
  nand2 gate974(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate975(.a(s_13), .b(gate498inter3), .O(gate498inter10));
  nor2  gate976(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate977(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate978(.a(gate498inter12), .b(gate498inter1), .O(N1747));
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );

  xor2  gate1833(.a(N1713), .b(N1680), .O(gate500inter0));
  nand2 gate1834(.a(gate500inter0), .b(s_136), .O(gate500inter1));
  and2  gate1835(.a(N1713), .b(N1680), .O(gate500inter2));
  inv1  gate1836(.a(s_136), .O(gate500inter3));
  inv1  gate1837(.a(s_137), .O(gate500inter4));
  nand2 gate1838(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1839(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1840(.a(N1680), .O(gate500inter7));
  inv1  gate1841(.a(N1713), .O(gate500inter8));
  nand2 gate1842(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1843(.a(s_137), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1844(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1845(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1846(.a(gate500inter12), .b(gate500inter1), .O(N1751));
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate1707(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate1708(.a(gate503inter0), .b(s_118), .O(gate503inter1));
  and2  gate1709(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate1710(.a(s_118), .O(gate503inter3));
  inv1  gate1711(.a(s_119), .O(gate503inter4));
  nand2 gate1712(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1713(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1714(.a(N1697), .O(gate503inter7));
  inv1  gate1715(.a(N1727), .O(gate503inter8));
  nand2 gate1716(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1717(.a(s_119), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1718(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1719(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1720(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );

  xor2  gate2001(.a(N1761), .b(N1661), .O(gate518inter0));
  nand2 gate2002(.a(gate518inter0), .b(s_160), .O(gate518inter1));
  and2  gate2003(.a(N1761), .b(N1661), .O(gate518inter2));
  inv1  gate2004(.a(s_160), .O(gate518inter3));
  inv1  gate2005(.a(s_161), .O(gate518inter4));
  nand2 gate2006(.a(gate518inter4), .b(gate518inter3), .O(gate518inter5));
  nor2  gate2007(.a(gate518inter5), .b(gate518inter2), .O(gate518inter6));
  inv1  gate2008(.a(N1661), .O(gate518inter7));
  inv1  gate2009(.a(N1761), .O(gate518inter8));
  nand2 gate2010(.a(gate518inter8), .b(gate518inter7), .O(gate518inter9));
  nand2 gate2011(.a(s_161), .b(gate518inter3), .O(gate518inter10));
  nor2  gate2012(.a(gate518inter10), .b(gate518inter9), .O(gate518inter11));
  nor2  gate2013(.a(gate518inter11), .b(gate518inter6), .O(gate518inter12));
  nand2 gate2014(.a(gate518inter12), .b(gate518inter1), .O(N1791));
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );

  xor2  gate2057(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate2058(.a(gate520inter0), .b(s_168), .O(gate520inter1));
  and2  gate2059(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate2060(.a(s_168), .O(gate520inter3));
  inv1  gate2061(.a(s_169), .O(gate520inter4));
  nand2 gate2062(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate2063(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate2064(.a(N1751), .O(gate520inter7));
  inv1  gate2065(.a(N1155), .O(gate520inter8));
  nand2 gate2066(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate2067(.a(s_169), .b(gate520inter3), .O(gate520inter10));
  nor2  gate2068(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate2069(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate2070(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate1413(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate1414(.a(gate522inter0), .b(s_76), .O(gate522inter1));
  and2  gate1415(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate1416(.a(s_76), .O(gate522inter3));
  inv1  gate1417(.a(s_77), .O(gate522inter4));
  nand2 gate1418(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate1419(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate1420(.a(N1740), .O(gate522inter7));
  inv1  gate1421(.a(N1769), .O(gate522inter8));
  nand2 gate1422(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate1423(.a(s_77), .b(gate522inter3), .O(gate522inter10));
  nor2  gate1424(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate1425(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate1426(.a(gate522inter12), .b(gate522inter1), .O(N1798));
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );

  xor2  gate1021(.a(N1764), .b(N1792), .O(gate530inter0));
  nand2 gate1022(.a(gate530inter0), .b(s_20), .O(gate530inter1));
  and2  gate1023(.a(N1764), .b(N1792), .O(gate530inter2));
  inv1  gate1024(.a(s_20), .O(gate530inter3));
  inv1  gate1025(.a(s_21), .O(gate530inter4));
  nand2 gate1026(.a(gate530inter4), .b(gate530inter3), .O(gate530inter5));
  nor2  gate1027(.a(gate530inter5), .b(gate530inter2), .O(gate530inter6));
  inv1  gate1028(.a(N1792), .O(gate530inter7));
  inv1  gate1029(.a(N1764), .O(gate530inter8));
  nand2 gate1030(.a(gate530inter8), .b(gate530inter7), .O(gate530inter9));
  nand2 gate1031(.a(s_21), .b(gate530inter3), .O(gate530inter10));
  nor2  gate1032(.a(gate530inter10), .b(gate530inter9), .O(gate530inter11));
  nor2  gate1033(.a(gate530inter11), .b(gate530inter6), .O(gate530inter12));
  nand2 gate1034(.a(gate530inter12), .b(gate530inter1), .O(N1815));
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );

  xor2  gate1343(.a(N1822), .b(N1419), .O(gate543inter0));
  nand2 gate1344(.a(gate543inter0), .b(s_66), .O(gate543inter1));
  and2  gate1345(.a(N1822), .b(N1419), .O(gate543inter2));
  inv1  gate1346(.a(s_66), .O(gate543inter3));
  inv1  gate1347(.a(s_67), .O(gate543inter4));
  nand2 gate1348(.a(gate543inter4), .b(gate543inter3), .O(gate543inter5));
  nor2  gate1349(.a(gate543inter5), .b(gate543inter2), .O(gate543inter6));
  inv1  gate1350(.a(N1419), .O(gate543inter7));
  inv1  gate1351(.a(N1822), .O(gate543inter8));
  nand2 gate1352(.a(gate543inter8), .b(gate543inter7), .O(gate543inter9));
  nand2 gate1353(.a(s_67), .b(gate543inter3), .O(gate543inter10));
  nor2  gate1354(.a(gate543inter10), .b(gate543inter9), .O(gate543inter11));
  nor2  gate1355(.a(gate543inter11), .b(gate543inter6), .O(gate543inter12));
  nand2 gate1356(.a(gate543inter12), .b(gate543inter1), .O(N1848));

  xor2  gate979(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate980(.a(gate544inter0), .b(s_14), .O(gate544inter1));
  and2  gate981(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate982(.a(s_14), .O(gate544inter3));
  inv1  gate983(.a(s_15), .O(gate544inter4));
  nand2 gate984(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate985(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate986(.a(N1416), .O(gate544inter7));
  inv1  gate987(.a(N1824), .O(gate544inter8));
  nand2 gate988(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate989(.a(s_15), .b(gate544inter3), .O(gate544inter10));
  nor2  gate990(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate991(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate992(.a(gate544inter12), .b(gate544inter1), .O(N1849));
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );

  xor2  gate1119(.a(N1837), .b(N1808), .O(gate556inter0));
  nand2 gate1120(.a(gate556inter0), .b(s_34), .O(gate556inter1));
  and2  gate1121(.a(N1837), .b(N1808), .O(gate556inter2));
  inv1  gate1122(.a(s_34), .O(gate556inter3));
  inv1  gate1123(.a(s_35), .O(gate556inter4));
  nand2 gate1124(.a(gate556inter4), .b(gate556inter3), .O(gate556inter5));
  nor2  gate1125(.a(gate556inter5), .b(gate556inter2), .O(gate556inter6));
  inv1  gate1126(.a(N1808), .O(gate556inter7));
  inv1  gate1127(.a(N1837), .O(gate556inter8));
  nand2 gate1128(.a(gate556inter8), .b(gate556inter7), .O(gate556inter9));
  nand2 gate1129(.a(s_35), .b(gate556inter3), .O(gate556inter10));
  nor2  gate1130(.a(gate556inter10), .b(gate556inter9), .O(gate556inter11));
  nor2  gate1131(.a(gate556inter11), .b(gate556inter6), .O(gate556inter12));
  nand2 gate1132(.a(gate556inter12), .b(gate556inter1), .O(N1875));
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );

  xor2  gate2281(.a(N1768), .b(N1841), .O(gate559inter0));
  nand2 gate2282(.a(gate559inter0), .b(s_200), .O(gate559inter1));
  and2  gate2283(.a(N1768), .b(N1841), .O(gate559inter2));
  inv1  gate2284(.a(s_200), .O(gate559inter3));
  inv1  gate2285(.a(s_201), .O(gate559inter4));
  nand2 gate2286(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate2287(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate2288(.a(N1841), .O(gate559inter7));
  inv1  gate2289(.a(N1768), .O(gate559inter8));
  nand2 gate2290(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate2291(.a(s_201), .b(gate559inter3), .O(gate559inter10));
  nor2  gate2292(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate2293(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate2294(.a(gate559inter12), .b(gate559inter1), .O(N1882));
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );

  xor2  gate1791(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate1792(.a(gate562inter0), .b(s_130), .O(gate562inter1));
  and2  gate1793(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate1794(.a(s_130), .O(gate562inter3));
  inv1  gate1795(.a(s_131), .O(gate562inter4));
  nand2 gate1796(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate1797(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate1798(.a(N1643), .O(gate562inter7));
  inv1  gate1799(.a(N1856), .O(gate562inter8));
  nand2 gate1800(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate1801(.a(s_131), .b(gate562inter3), .O(gate562inter10));
  nor2  gate1802(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate1803(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate1804(.a(gate562inter12), .b(gate562inter1), .O(N1885));

  xor2  gate1931(.a(N290), .b(N1830), .O(gate563inter0));
  nand2 gate1932(.a(gate563inter0), .b(s_150), .O(gate563inter1));
  and2  gate1933(.a(N290), .b(N1830), .O(gate563inter2));
  inv1  gate1934(.a(s_150), .O(gate563inter3));
  inv1  gate1935(.a(s_151), .O(gate563inter4));
  nand2 gate1936(.a(gate563inter4), .b(gate563inter3), .O(gate563inter5));
  nor2  gate1937(.a(gate563inter5), .b(gate563inter2), .O(gate563inter6));
  inv1  gate1938(.a(N1830), .O(gate563inter7));
  inv1  gate1939(.a(N290), .O(gate563inter8));
  nand2 gate1940(.a(gate563inter8), .b(gate563inter7), .O(gate563inter9));
  nand2 gate1941(.a(s_151), .b(gate563inter3), .O(gate563inter10));
  nor2  gate1942(.a(gate563inter10), .b(gate563inter9), .O(gate563inter11));
  nor2  gate1943(.a(gate563inter11), .b(gate563inter6), .O(gate563inter12));
  nand2 gate1944(.a(gate563inter12), .b(gate563inter1), .O(N1889));
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate1259(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate1260(.a(gate565inter0), .b(s_54), .O(gate565inter1));
  and2  gate1261(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate1262(.a(s_54), .O(gate565inter3));
  inv1  gate1263(.a(s_55), .O(gate565inter4));
  nand2 gate1264(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate1265(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate1266(.a(N1838), .O(gate565inter7));
  inv1  gate1267(.a(N1785), .O(gate565inter8));
  nand2 gate1268(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate1269(.a(s_55), .b(gate565inter3), .O(gate565inter10));
  nor2  gate1270(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate1271(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate1272(.a(gate565inter12), .b(gate565inter1), .O(N1896));
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );

  xor2  gate1315(.a(N1885), .b(N1855), .O(gate572inter0));
  nand2 gate1316(.a(gate572inter0), .b(s_62), .O(gate572inter1));
  and2  gate1317(.a(N1885), .b(N1855), .O(gate572inter2));
  inv1  gate1318(.a(s_62), .O(gate572inter3));
  inv1  gate1319(.a(s_63), .O(gate572inter4));
  nand2 gate1320(.a(gate572inter4), .b(gate572inter3), .O(gate572inter5));
  nor2  gate1321(.a(gate572inter5), .b(gate572inter2), .O(gate572inter6));
  inv1  gate1322(.a(N1855), .O(gate572inter7));
  inv1  gate1323(.a(N1885), .O(gate572inter8));
  nand2 gate1324(.a(gate572inter8), .b(gate572inter7), .O(gate572inter9));
  nand2 gate1325(.a(s_63), .b(gate572inter3), .O(gate572inter10));
  nor2  gate1326(.a(gate572inter10), .b(gate572inter9), .O(gate572inter11));
  nor2  gate1327(.a(gate572inter11), .b(gate572inter6), .O(gate572inter12));
  nand2 gate1328(.a(gate572inter12), .b(gate572inter1), .O(N1913));
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );

  xor2  gate1091(.a(N920), .b(N1869), .O(gate576inter0));
  nand2 gate1092(.a(gate576inter0), .b(s_30), .O(gate576inter1));
  and2  gate1093(.a(N920), .b(N1869), .O(gate576inter2));
  inv1  gate1094(.a(s_30), .O(gate576inter3));
  inv1  gate1095(.a(s_31), .O(gate576inter4));
  nand2 gate1096(.a(gate576inter4), .b(gate576inter3), .O(gate576inter5));
  nor2  gate1097(.a(gate576inter5), .b(gate576inter2), .O(gate576inter6));
  inv1  gate1098(.a(N1869), .O(gate576inter7));
  inv1  gate1099(.a(N920), .O(gate576inter8));
  nand2 gate1100(.a(gate576inter8), .b(gate576inter7), .O(gate576inter9));
  nand2 gate1101(.a(s_31), .b(gate576inter3), .O(gate576inter10));
  nor2  gate1102(.a(gate576inter10), .b(gate576inter9), .O(gate576inter11));
  nor2  gate1103(.a(gate576inter11), .b(gate576inter6), .O(gate576inter12));
  nand2 gate1104(.a(gate576inter12), .b(gate576inter1), .O(N1921));
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate2085(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate2086(.a(gate579inter0), .b(s_172), .O(gate579inter1));
  and2  gate2087(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate2088(.a(s_172), .O(gate579inter3));
  inv1  gate2089(.a(s_173), .O(gate579inter4));
  nand2 gate2090(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate2091(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate2092(.a(N1714), .O(gate579inter7));
  inv1  gate2093(.a(N1895), .O(gate579inter8));
  nand2 gate2094(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate2095(.a(s_173), .b(gate579inter3), .O(gate579inter10));
  nor2  gate2096(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate2097(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate2098(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate2211(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate2212(.a(gate596inter0), .b(s_190), .O(gate596inter1));
  and2  gate2213(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate2214(.a(s_190), .O(gate596inter3));
  inv1  gate2215(.a(s_191), .O(gate596inter4));
  nand2 gate2216(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate2217(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate2218(.a(N1930), .O(gate596inter7));
  inv1  gate2219(.a(N917), .O(gate596inter8));
  nand2 gate2220(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate2221(.a(s_191), .b(gate596inter3), .O(gate596inter10));
  nor2  gate2222(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate2223(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate2224(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );

  xor2  gate895(.a(N1937), .b(N1944), .O(gate605inter0));
  nand2 gate896(.a(gate605inter0), .b(s_2), .O(gate605inter1));
  and2  gate897(.a(N1937), .b(N1944), .O(gate605inter2));
  inv1  gate898(.a(s_2), .O(gate605inter3));
  inv1  gate899(.a(s_3), .O(gate605inter4));
  nand2 gate900(.a(gate605inter4), .b(gate605inter3), .O(gate605inter5));
  nor2  gate901(.a(gate605inter5), .b(gate605inter2), .O(gate605inter6));
  inv1  gate902(.a(N1944), .O(gate605inter7));
  inv1  gate903(.a(N1937), .O(gate605inter8));
  nand2 gate904(.a(gate605inter8), .b(gate605inter7), .O(gate605inter9));
  nand2 gate905(.a(s_3), .b(gate605inter3), .O(gate605inter10));
  nor2  gate906(.a(gate605inter10), .b(gate605inter9), .O(gate605inter11));
  nor2  gate907(.a(gate605inter11), .b(gate605inter6), .O(gate605inter12));
  nand2 gate908(.a(gate605inter12), .b(gate605inter1), .O(N2000));
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );

  xor2  gate2155(.a(N1999), .b(N1898), .O(gate621inter0));
  nand2 gate2156(.a(gate621inter0), .b(s_182), .O(gate621inter1));
  and2  gate2157(.a(N1999), .b(N1898), .O(gate621inter2));
  inv1  gate2158(.a(s_182), .O(gate621inter3));
  inv1  gate2159(.a(s_183), .O(gate621inter4));
  nand2 gate2160(.a(gate621inter4), .b(gate621inter3), .O(gate621inter5));
  nor2  gate2161(.a(gate621inter5), .b(gate621inter2), .O(gate621inter6));
  inv1  gate2162(.a(N1898), .O(gate621inter7));
  inv1  gate2163(.a(N1999), .O(gate621inter8));
  nand2 gate2164(.a(gate621inter8), .b(gate621inter7), .O(gate621inter9));
  nand2 gate2165(.a(s_183), .b(gate621inter3), .O(gate621inter10));
  nor2  gate2166(.a(gate621inter10), .b(gate621inter9), .O(gate621inter11));
  nor2  gate2167(.a(gate621inter11), .b(gate621inter6), .O(gate621inter12));
  nand2 gate2168(.a(gate621inter12), .b(gate621inter1), .O(N2020));
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );

  xor2  gate2029(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate2030(.a(gate627inter0), .b(s_164), .O(gate627inter1));
  and2  gate2031(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate2032(.a(s_164), .O(gate627inter3));
  inv1  gate2033(.a(s_165), .O(gate627inter4));
  nand2 gate2034(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate2035(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate2036(.a(N1975), .O(gate627inter7));
  inv1  gate2037(.a(N2008), .O(gate627inter8));
  nand2 gate2038(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate2039(.a(s_165), .b(gate627inter3), .O(gate627inter10));
  nor2  gate2040(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate2041(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate2042(.a(gate627inter12), .b(gate627inter1), .O(N2026));

  xor2  gate1805(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1806(.a(gate628inter0), .b(s_132), .O(gate628inter1));
  and2  gate1807(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1808(.a(s_132), .O(gate628inter3));
  inv1  gate1809(.a(s_133), .O(gate628inter4));
  nand2 gate1810(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1811(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1812(.a(N1977), .O(gate628inter7));
  inv1  gate1813(.a(N2009), .O(gate628inter8));
  nand2 gate1814(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1815(.a(s_133), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1816(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1817(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1818(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );

  xor2  gate1595(.a(N2022), .b(N2039), .O(gate642inter0));
  nand2 gate1596(.a(gate642inter0), .b(s_102), .O(gate642inter1));
  and2  gate1597(.a(N2022), .b(N2039), .O(gate642inter2));
  inv1  gate1598(.a(s_102), .O(gate642inter3));
  inv1  gate1599(.a(s_103), .O(gate642inter4));
  nand2 gate1600(.a(gate642inter4), .b(gate642inter3), .O(gate642inter5));
  nor2  gate1601(.a(gate642inter5), .b(gate642inter2), .O(gate642inter6));
  inv1  gate1602(.a(N2039), .O(gate642inter7));
  inv1  gate1603(.a(N2022), .O(gate642inter8));
  nand2 gate1604(.a(gate642inter8), .b(gate642inter7), .O(gate642inter9));
  nand2 gate1605(.a(s_103), .b(gate642inter3), .O(gate642inter10));
  nor2  gate1606(.a(gate642inter10), .b(gate642inter9), .O(gate642inter11));
  nor2  gate1607(.a(gate642inter11), .b(gate642inter6), .O(gate642inter12));
  nand2 gate1608(.a(gate642inter12), .b(gate642inter1), .O(N2061));
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );

  xor2  gate1049(.a(N916), .b(N2148), .O(gate665inter0));
  nand2 gate1050(.a(gate665inter0), .b(s_24), .O(gate665inter1));
  and2  gate1051(.a(N916), .b(N2148), .O(gate665inter2));
  inv1  gate1052(.a(s_24), .O(gate665inter3));
  inv1  gate1053(.a(s_25), .O(gate665inter4));
  nand2 gate1054(.a(gate665inter4), .b(gate665inter3), .O(gate665inter5));
  nor2  gate1055(.a(gate665inter5), .b(gate665inter2), .O(gate665inter6));
  inv1  gate1056(.a(N2148), .O(gate665inter7));
  inv1  gate1057(.a(N916), .O(gate665inter8));
  nand2 gate1058(.a(gate665inter8), .b(gate665inter7), .O(gate665inter9));
  nand2 gate1059(.a(s_25), .b(gate665inter3), .O(gate665inter10));
  nor2  gate1060(.a(gate665inter10), .b(gate665inter9), .O(gate665inter11));
  nor2  gate1061(.a(gate665inter11), .b(gate665inter6), .O(gate665inter12));
  nand2 gate1062(.a(gate665inter12), .b(gate665inter1), .O(N2216));
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );

  xor2  gate1399(.a(N913), .b(N2205), .O(gate671inter0));
  nand2 gate1400(.a(gate671inter0), .b(s_74), .O(gate671inter1));
  and2  gate1401(.a(N913), .b(N2205), .O(gate671inter2));
  inv1  gate1402(.a(s_74), .O(gate671inter3));
  inv1  gate1403(.a(s_75), .O(gate671inter4));
  nand2 gate1404(.a(gate671inter4), .b(gate671inter3), .O(gate671inter5));
  nor2  gate1405(.a(gate671inter5), .b(gate671inter2), .O(gate671inter6));
  inv1  gate1406(.a(N2205), .O(gate671inter7));
  inv1  gate1407(.a(N913), .O(gate671inter8));
  nand2 gate1408(.a(gate671inter8), .b(gate671inter7), .O(gate671inter9));
  nand2 gate1409(.a(s_75), .b(gate671inter3), .O(gate671inter10));
  nor2  gate1410(.a(gate671inter10), .b(gate671inter9), .O(gate671inter11));
  nor2  gate1411(.a(gate671inter11), .b(gate671inter6), .O(gate671inter12));
  nand2 gate1412(.a(gate671inter12), .b(gate671inter1), .O(N2226));
inv1 gate672( .a(N2205), .O(N2227) );

  xor2  gate1371(.a(N914), .b(N2202), .O(gate673inter0));
  nand2 gate1372(.a(gate673inter0), .b(s_70), .O(gate673inter1));
  and2  gate1373(.a(N914), .b(N2202), .O(gate673inter2));
  inv1  gate1374(.a(s_70), .O(gate673inter3));
  inv1  gate1375(.a(s_71), .O(gate673inter4));
  nand2 gate1376(.a(gate673inter4), .b(gate673inter3), .O(gate673inter5));
  nor2  gate1377(.a(gate673inter5), .b(gate673inter2), .O(gate673inter6));
  inv1  gate1378(.a(N2202), .O(gate673inter7));
  inv1  gate1379(.a(N914), .O(gate673inter8));
  nand2 gate1380(.a(gate673inter8), .b(gate673inter7), .O(gate673inter9));
  nand2 gate1381(.a(s_71), .b(gate673inter3), .O(gate673inter10));
  nor2  gate1382(.a(gate673inter10), .b(gate673inter9), .O(gate673inter11));
  nor2  gate1383(.a(gate673inter11), .b(gate673inter6), .O(gate673inter12));
  nand2 gate1384(.a(gate673inter12), .b(gate673inter1), .O(N2228));
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );

  xor2  gate1539(.a(N2217), .b(N664), .O(gate676inter0));
  nand2 gate1540(.a(gate676inter0), .b(s_94), .O(gate676inter1));
  and2  gate1541(.a(N2217), .b(N664), .O(gate676inter2));
  inv1  gate1542(.a(s_94), .O(gate676inter3));
  inv1  gate1543(.a(s_95), .O(gate676inter4));
  nand2 gate1544(.a(gate676inter4), .b(gate676inter3), .O(gate676inter5));
  nor2  gate1545(.a(gate676inter5), .b(gate676inter2), .O(gate676inter6));
  inv1  gate1546(.a(N664), .O(gate676inter7));
  inv1  gate1547(.a(N2217), .O(gate676inter8));
  nand2 gate1548(.a(gate676inter8), .b(gate676inter7), .O(gate676inter9));
  nand2 gate1549(.a(s_95), .b(gate676inter3), .O(gate676inter10));
  nor2  gate1550(.a(gate676inter10), .b(gate676inter9), .O(gate676inter11));
  nor2  gate1551(.a(gate676inter11), .b(gate676inter6), .O(gate676inter12));
  nand2 gate1552(.a(gate676inter12), .b(gate676inter1), .O(N2231));
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );

  xor2  gate2043(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate2044(.a(gate678inter0), .b(s_166), .O(gate678inter1));
  and2  gate2045(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate2046(.a(s_166), .O(gate678inter3));
  inv1  gate2047(.a(s_167), .O(gate678inter4));
  nand2 gate2048(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate2049(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate2050(.a(N1252), .O(gate678inter7));
  inv1  gate2051(.a(N2225), .O(gate678inter8));
  nand2 gate2052(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate2053(.a(s_167), .b(gate678inter3), .O(gate678inter10));
  nor2  gate2054(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate2055(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate2056(.a(gate678inter12), .b(gate678inter1), .O(N2233));
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );

  xor2  gate1847(.a(N2229), .b(N658), .O(gate680inter0));
  nand2 gate1848(.a(gate680inter0), .b(s_138), .O(gate680inter1));
  and2  gate1849(.a(N2229), .b(N658), .O(gate680inter2));
  inv1  gate1850(.a(s_138), .O(gate680inter3));
  inv1  gate1851(.a(s_139), .O(gate680inter4));
  nand2 gate1852(.a(gate680inter4), .b(gate680inter3), .O(gate680inter5));
  nor2  gate1853(.a(gate680inter5), .b(gate680inter2), .O(gate680inter6));
  inv1  gate1854(.a(N658), .O(gate680inter7));
  inv1  gate1855(.a(N2229), .O(gate680inter8));
  nand2 gate1856(.a(gate680inter8), .b(gate680inter7), .O(gate680inter9));
  nand2 gate1857(.a(s_139), .b(gate680inter3), .O(gate680inter10));
  nor2  gate1858(.a(gate680inter10), .b(gate680inter9), .O(gate680inter11));
  nor2  gate1859(.a(gate680inter11), .b(gate680inter6), .O(gate680inter12));
  nand2 gate1860(.a(gate680inter12), .b(gate680inter1), .O(N2235));
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );

  xor2  gate881(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate882(.a(gate684inter0), .b(s_0), .O(gate684inter1));
  and2  gate883(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate884(.a(s_0), .O(gate684inter3));
  inv1  gate885(.a(s_1), .O(gate684inter4));
  nand2 gate886(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate887(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate888(.a(N2224), .O(gate684inter7));
  inv1  gate889(.a(N2233), .O(gate684inter8));
  nand2 gate890(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate891(.a(s_1), .b(gate684inter3), .O(gate684inter10));
  nor2  gate892(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate893(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate894(.a(gate684inter12), .b(gate684inter1), .O(N2241));
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );

  xor2  gate2127(.a(N534), .b(N2558), .O(gate750inter0));
  nand2 gate2128(.a(gate750inter0), .b(s_178), .O(gate750inter1));
  and2  gate2129(.a(N534), .b(N2558), .O(gate750inter2));
  inv1  gate2130(.a(s_178), .O(gate750inter3));
  inv1  gate2131(.a(s_179), .O(gate750inter4));
  nand2 gate2132(.a(gate750inter4), .b(gate750inter3), .O(gate750inter5));
  nor2  gate2133(.a(gate750inter5), .b(gate750inter2), .O(gate750inter6));
  inv1  gate2134(.a(N2558), .O(gate750inter7));
  inv1  gate2135(.a(N534), .O(gate750inter8));
  nand2 gate2136(.a(gate750inter8), .b(gate750inter7), .O(gate750inter9));
  nand2 gate2137(.a(s_179), .b(gate750inter3), .O(gate750inter10));
  nor2  gate2138(.a(gate750inter10), .b(gate750inter9), .O(gate750inter11));
  nor2  gate2139(.a(gate750inter11), .b(gate750inter6), .O(gate750inter12));
  nand2 gate2140(.a(gate750inter12), .b(gate750inter1), .O(N2669));
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );

  xor2  gate2197(.a(N543), .b(N2570), .O(gate758inter0));
  nand2 gate2198(.a(gate758inter0), .b(s_188), .O(gate758inter1));
  and2  gate2199(.a(N543), .b(N2570), .O(gate758inter2));
  inv1  gate2200(.a(s_188), .O(gate758inter3));
  inv1  gate2201(.a(s_189), .O(gate758inter4));
  nand2 gate2202(.a(gate758inter4), .b(gate758inter3), .O(gate758inter5));
  nor2  gate2203(.a(gate758inter5), .b(gate758inter2), .O(gate758inter6));
  inv1  gate2204(.a(N2570), .O(gate758inter7));
  inv1  gate2205(.a(N543), .O(gate758inter8));
  nand2 gate2206(.a(gate758inter8), .b(gate758inter7), .O(gate758inter9));
  nand2 gate2207(.a(s_189), .b(gate758inter3), .O(gate758inter10));
  nor2  gate2208(.a(gate758inter10), .b(gate758inter9), .O(gate758inter11));
  nor2  gate2209(.a(gate758inter11), .b(gate758inter6), .O(gate758inter12));
  nand2 gate2210(.a(gate758inter12), .b(gate758inter1), .O(N2682));
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );

  xor2  gate1301(.a(N538), .b(N2639), .O(gate769inter0));
  nand2 gate1302(.a(gate769inter0), .b(s_60), .O(gate769inter1));
  and2  gate1303(.a(N538), .b(N2639), .O(gate769inter2));
  inv1  gate1304(.a(s_60), .O(gate769inter3));
  inv1  gate1305(.a(s_61), .O(gate769inter4));
  nand2 gate1306(.a(gate769inter4), .b(gate769inter3), .O(gate769inter5));
  nor2  gate1307(.a(gate769inter5), .b(gate769inter2), .O(gate769inter6));
  inv1  gate1308(.a(N2639), .O(gate769inter7));
  inv1  gate1309(.a(N538), .O(gate769inter8));
  nand2 gate1310(.a(gate769inter8), .b(gate769inter7), .O(gate769inter9));
  nand2 gate1311(.a(s_61), .b(gate769inter3), .O(gate769inter10));
  nor2  gate1312(.a(gate769inter10), .b(gate769inter9), .O(gate769inter11));
  nor2  gate1313(.a(gate769inter11), .b(gate769inter6), .O(gate769inter12));
  nand2 gate1314(.a(gate769inter12), .b(gate769inter1), .O(N2724));
inv1 gate770( .a(N2639), .O(N2725) );

  xor2  gate1245(.a(N539), .b(N2642), .O(gate771inter0));
  nand2 gate1246(.a(gate771inter0), .b(s_52), .O(gate771inter1));
  and2  gate1247(.a(N539), .b(N2642), .O(gate771inter2));
  inv1  gate1248(.a(s_52), .O(gate771inter3));
  inv1  gate1249(.a(s_53), .O(gate771inter4));
  nand2 gate1250(.a(gate771inter4), .b(gate771inter3), .O(gate771inter5));
  nor2  gate1251(.a(gate771inter5), .b(gate771inter2), .O(gate771inter6));
  inv1  gate1252(.a(N2642), .O(gate771inter7));
  inv1  gate1253(.a(N539), .O(gate771inter8));
  nand2 gate1254(.a(gate771inter8), .b(gate771inter7), .O(gate771inter9));
  nand2 gate1255(.a(s_53), .b(gate771inter3), .O(gate771inter10));
  nor2  gate1256(.a(gate771inter10), .b(gate771inter9), .O(gate771inter11));
  nor2  gate1257(.a(gate771inter11), .b(gate771inter6), .O(gate771inter12));
  nand2 gate1258(.a(gate771inter12), .b(gate771inter1), .O(N2726));
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate1819(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate1820(.a(gate788inter0), .b(s_134), .O(gate788inter1));
  and2  gate1821(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate1822(.a(s_134), .O(gate788inter3));
  inv1  gate1823(.a(s_135), .O(gate788inter4));
  nand2 gate1824(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate1825(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate1826(.a(N385), .O(gate788inter7));
  inv1  gate1827(.a(N2689), .O(gate788inter8));
  nand2 gate1828(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate1829(.a(s_135), .b(gate788inter3), .O(gate788inter10));
  nor2  gate1830(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate1831(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate1832(.a(gate788inter12), .b(gate788inter1), .O(N2743));
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );

  xor2  gate1987(.a(N2731), .b(N364), .O(gate801inter0));
  nand2 gate1988(.a(gate801inter0), .b(s_158), .O(gate801inter1));
  and2  gate1989(.a(N2731), .b(N364), .O(gate801inter2));
  inv1  gate1990(.a(s_158), .O(gate801inter3));
  inv1  gate1991(.a(s_159), .O(gate801inter4));
  nand2 gate1992(.a(gate801inter4), .b(gate801inter3), .O(gate801inter5));
  nor2  gate1993(.a(gate801inter5), .b(gate801inter2), .O(gate801inter6));
  inv1  gate1994(.a(N364), .O(gate801inter7));
  inv1  gate1995(.a(N2731), .O(gate801inter8));
  nand2 gate1996(.a(gate801inter8), .b(gate801inter7), .O(gate801inter9));
  nand2 gate1997(.a(s_159), .b(gate801inter3), .O(gate801inter10));
  nor2  gate1998(.a(gate801inter10), .b(gate801inter9), .O(gate801inter11));
  nor2  gate1999(.a(gate801inter11), .b(gate801inter6), .O(gate801inter12));
  nand2 gate2000(.a(gate801inter12), .b(gate801inter1), .O(N2760));
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );

  xor2  gate1553(.a(N2734), .b(N2682), .O(gate803inter0));
  nand2 gate1554(.a(gate803inter0), .b(s_96), .O(gate803inter1));
  and2  gate1555(.a(N2734), .b(N2682), .O(gate803inter2));
  inv1  gate1556(.a(s_96), .O(gate803inter3));
  inv1  gate1557(.a(s_97), .O(gate803inter4));
  nand2 gate1558(.a(gate803inter4), .b(gate803inter3), .O(gate803inter5));
  nor2  gate1559(.a(gate803inter5), .b(gate803inter2), .O(gate803inter6));
  inv1  gate1560(.a(N2682), .O(gate803inter7));
  inv1  gate1561(.a(N2734), .O(gate803inter8));
  nand2 gate1562(.a(gate803inter8), .b(gate803inter7), .O(gate803inter9));
  nand2 gate1563(.a(s_97), .b(gate803inter3), .O(gate803inter10));
  nor2  gate1564(.a(gate803inter10), .b(gate803inter9), .O(gate803inter11));
  nor2  gate1565(.a(gate803inter11), .b(gate803inter6), .O(gate803inter12));
  nand2 gate1566(.a(gate803inter12), .b(gate803inter1), .O(N2762));
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );

  xor2  gate1329(.a(N2742), .b(N382), .O(gate807inter0));
  nand2 gate1330(.a(gate807inter0), .b(s_64), .O(gate807inter1));
  and2  gate1331(.a(N2742), .b(N382), .O(gate807inter2));
  inv1  gate1332(.a(s_64), .O(gate807inter3));
  inv1  gate1333(.a(s_65), .O(gate807inter4));
  nand2 gate1334(.a(gate807inter4), .b(gate807inter3), .O(gate807inter5));
  nor2  gate1335(.a(gate807inter5), .b(gate807inter2), .O(gate807inter6));
  inv1  gate1336(.a(N382), .O(gate807inter7));
  inv1  gate1337(.a(N2742), .O(gate807inter8));
  nand2 gate1338(.a(gate807inter8), .b(gate807inter7), .O(gate807inter9));
  nand2 gate1339(.a(s_65), .b(gate807inter3), .O(gate807inter10));
  nor2  gate1340(.a(gate807inter10), .b(gate807inter9), .O(gate807inter11));
  nor2  gate1341(.a(gate807inter11), .b(gate807inter6), .O(gate807inter12));
  nand2 gate1342(.a(gate807inter12), .b(gate807inter1), .O(N2766));
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );

  xor2  gate1637(.a(N2744), .b(N2690), .O(gate809inter0));
  nand2 gate1638(.a(gate809inter0), .b(s_108), .O(gate809inter1));
  and2  gate1639(.a(N2744), .b(N2690), .O(gate809inter2));
  inv1  gate1640(.a(s_108), .O(gate809inter3));
  inv1  gate1641(.a(s_109), .O(gate809inter4));
  nand2 gate1642(.a(gate809inter4), .b(gate809inter3), .O(gate809inter5));
  nor2  gate1643(.a(gate809inter5), .b(gate809inter2), .O(gate809inter6));
  inv1  gate1644(.a(N2690), .O(gate809inter7));
  inv1  gate1645(.a(N2744), .O(gate809inter8));
  nand2 gate1646(.a(gate809inter8), .b(gate809inter7), .O(gate809inter9));
  nand2 gate1647(.a(s_109), .b(gate809inter3), .O(gate809inter10));
  nor2  gate1648(.a(gate809inter10), .b(gate809inter9), .O(gate809inter11));
  nor2  gate1649(.a(gate809inter11), .b(gate809inter6), .O(gate809inter12));
  nand2 gate1650(.a(gate809inter12), .b(gate809inter1), .O(N2768));
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );

  xor2  gate1161(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate1162(.a(gate813inter0), .b(s_40), .O(gate813inter1));
  and2  gate1163(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate1164(.a(s_40), .O(gate813inter3));
  inv1  gate1165(.a(s_41), .O(gate813inter4));
  nand2 gate1166(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate1167(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate1168(.a(N2726), .O(gate813inter7));
  inv1  gate1169(.a(N2758), .O(gate813inter8));
  nand2 gate1170(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate1171(.a(s_41), .b(gate813inter3), .O(gate813inter10));
  nor2  gate1172(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate1173(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate1174(.a(gate813inter12), .b(gate813inter1), .O(N2780));
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );

  xor2  gate2225(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate2226(.a(gate815inter0), .b(s_192), .O(gate815inter1));
  and2  gate2227(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate2228(.a(s_192), .O(gate815inter3));
  inv1  gate2229(.a(s_193), .O(gate815inter4));
  nand2 gate2230(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate2231(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate2232(.a(N2730), .O(gate815inter7));
  inv1  gate2233(.a(N2760), .O(gate815inter8));
  nand2 gate2234(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate2235(.a(s_193), .b(gate815inter3), .O(gate815inter10));
  nor2  gate2236(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate2237(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate2238(.a(gate815inter12), .b(gate815inter1), .O(N2782));
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );

  xor2  gate1651(.a(N2763), .b(N2735), .O(gate817inter0));
  nand2 gate1652(.a(gate817inter0), .b(s_110), .O(gate817inter1));
  and2  gate1653(.a(N2763), .b(N2735), .O(gate817inter2));
  inv1  gate1654(.a(s_110), .O(gate817inter3));
  inv1  gate1655(.a(s_111), .O(gate817inter4));
  nand2 gate1656(.a(gate817inter4), .b(gate817inter3), .O(gate817inter5));
  nor2  gate1657(.a(gate817inter5), .b(gate817inter2), .O(gate817inter6));
  inv1  gate1658(.a(N2735), .O(gate817inter7));
  inv1  gate1659(.a(N2763), .O(gate817inter8));
  nand2 gate1660(.a(gate817inter8), .b(gate817inter7), .O(gate817inter9));
  nand2 gate1661(.a(s_111), .b(gate817inter3), .O(gate817inter10));
  nor2  gate1662(.a(gate817inter10), .b(gate817inter9), .O(gate817inter11));
  nor2  gate1663(.a(gate817inter11), .b(gate817inter6), .O(gate817inter12));
  nand2 gate1664(.a(gate817inter12), .b(gate817inter1), .O(N2784));
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );

  xor2  gate1735(.a(N2765), .b(N2739), .O(gate819inter0));
  nand2 gate1736(.a(gate819inter0), .b(s_122), .O(gate819inter1));
  and2  gate1737(.a(N2765), .b(N2739), .O(gate819inter2));
  inv1  gate1738(.a(s_122), .O(gate819inter3));
  inv1  gate1739(.a(s_123), .O(gate819inter4));
  nand2 gate1740(.a(gate819inter4), .b(gate819inter3), .O(gate819inter5));
  nor2  gate1741(.a(gate819inter5), .b(gate819inter2), .O(gate819inter6));
  inv1  gate1742(.a(N2739), .O(gate819inter7));
  inv1  gate1743(.a(N2765), .O(gate819inter8));
  nand2 gate1744(.a(gate819inter8), .b(gate819inter7), .O(gate819inter9));
  nand2 gate1745(.a(s_123), .b(gate819inter3), .O(gate819inter10));
  nor2  gate1746(.a(gate819inter10), .b(gate819inter9), .O(gate819inter11));
  nor2  gate1747(.a(gate819inter11), .b(gate819inter6), .O(gate819inter12));
  nand2 gate1748(.a(gate819inter12), .b(gate819inter1), .O(N2786));
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );

  xor2  gate1665(.a(N2750), .b(N2747), .O(gate822inter0));
  nand2 gate1666(.a(gate822inter0), .b(s_112), .O(gate822inter1));
  and2  gate1667(.a(N2750), .b(N2747), .O(gate822inter2));
  inv1  gate1668(.a(s_112), .O(gate822inter3));
  inv1  gate1669(.a(s_113), .O(gate822inter4));
  nand2 gate1670(.a(gate822inter4), .b(gate822inter3), .O(gate822inter5));
  nor2  gate1671(.a(gate822inter5), .b(gate822inter2), .O(gate822inter6));
  inv1  gate1672(.a(N2747), .O(gate822inter7));
  inv1  gate1673(.a(N2750), .O(gate822inter8));
  nand2 gate1674(.a(gate822inter8), .b(gate822inter7), .O(gate822inter9));
  nand2 gate1675(.a(s_113), .b(gate822inter3), .O(gate822inter10));
  nor2  gate1676(.a(gate822inter10), .b(gate822inter9), .O(gate822inter11));
  nor2  gate1677(.a(gate822inter11), .b(gate822inter6), .O(gate822inter12));
  nand2 gate1678(.a(gate822inter12), .b(gate822inter1), .O(N2789));
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );

  xor2  gate1427(.a(N2018), .b(N2773), .O(gate824inter0));
  nand2 gate1428(.a(gate824inter0), .b(s_78), .O(gate824inter1));
  and2  gate1429(.a(N2018), .b(N2773), .O(gate824inter2));
  inv1  gate1430(.a(s_78), .O(gate824inter3));
  inv1  gate1431(.a(s_79), .O(gate824inter4));
  nand2 gate1432(.a(gate824inter4), .b(gate824inter3), .O(gate824inter5));
  nor2  gate1433(.a(gate824inter5), .b(gate824inter2), .O(gate824inter6));
  inv1  gate1434(.a(N2773), .O(gate824inter7));
  inv1  gate1435(.a(N2018), .O(gate824inter8));
  nand2 gate1436(.a(gate824inter8), .b(gate824inter7), .O(gate824inter9));
  nand2 gate1437(.a(s_79), .b(gate824inter3), .O(gate824inter10));
  nor2  gate1438(.a(gate824inter10), .b(gate824inter9), .O(gate824inter11));
  nor2  gate1439(.a(gate824inter11), .b(gate824inter6), .O(gate824inter12));
  nand2 gate1440(.a(gate824inter12), .b(gate824inter1), .O(N2807));
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );

  xor2  gate1609(.a(N2810), .b(N1968), .O(gate835inter0));
  nand2 gate1610(.a(gate835inter0), .b(s_104), .O(gate835inter1));
  and2  gate1611(.a(N2810), .b(N1968), .O(gate835inter2));
  inv1  gate1612(.a(s_104), .O(gate835inter3));
  inv1  gate1613(.a(s_105), .O(gate835inter4));
  nand2 gate1614(.a(gate835inter4), .b(gate835inter3), .O(gate835inter5));
  nor2  gate1615(.a(gate835inter5), .b(gate835inter2), .O(gate835inter6));
  inv1  gate1616(.a(N1968), .O(gate835inter7));
  inv1  gate1617(.a(N2810), .O(gate835inter8));
  nand2 gate1618(.a(gate835inter8), .b(gate835inter7), .O(gate835inter9));
  nand2 gate1619(.a(s_105), .b(gate835inter3), .O(gate835inter10));
  nor2  gate1620(.a(gate835inter10), .b(gate835inter9), .O(gate835inter11));
  nor2  gate1621(.a(gate835inter11), .b(gate835inter6), .O(gate835inter12));
  nand2 gate1622(.a(gate835inter12), .b(gate835inter1), .O(N2828));
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );

  xor2  gate1749(.a(N2860), .b(N1818), .O(gate854inter0));
  nand2 gate1750(.a(gate854inter0), .b(s_124), .O(gate854inter1));
  and2  gate1751(.a(N2860), .b(N1818), .O(gate854inter2));
  inv1  gate1752(.a(s_124), .O(gate854inter3));
  inv1  gate1753(.a(s_125), .O(gate854inter4));
  nand2 gate1754(.a(gate854inter4), .b(gate854inter3), .O(gate854inter5));
  nor2  gate1755(.a(gate854inter5), .b(gate854inter2), .O(gate854inter6));
  inv1  gate1756(.a(N1818), .O(gate854inter7));
  inv1  gate1757(.a(N2860), .O(gate854inter8));
  nand2 gate1758(.a(gate854inter8), .b(gate854inter7), .O(gate854inter9));
  nand2 gate1759(.a(s_125), .b(gate854inter3), .O(gate854inter10));
  nor2  gate1760(.a(gate854inter10), .b(gate854inter9), .O(gate854inter11));
  nor2  gate1761(.a(gate854inter11), .b(gate854inter6), .O(gate854inter12));
  nand2 gate1762(.a(gate854inter12), .b(gate854inter1), .O(N2869));
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate1287(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate1288(.a(gate860inter0), .b(s_58), .O(gate860inter1));
  and2  gate1289(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate1290(.a(s_58), .O(gate860inter3));
  inv1  gate1291(.a(s_59), .O(gate860inter4));
  nand2 gate1292(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate1293(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate1294(.a(N1933), .O(gate860inter7));
  inv1  gate1295(.a(N2862), .O(gate860inter8));
  nand2 gate1296(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate1297(.a(s_59), .b(gate860inter3), .O(gate860inter10));
  nor2  gate1298(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate1299(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate1300(.a(gate860inter12), .b(gate860inter1), .O(N2875));
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule