module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1121(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1122(.a(gate13inter0), .b(s_82), .O(gate13inter1));
  and2  gate1123(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1124(.a(s_82), .O(gate13inter3));
  inv1  gate1125(.a(s_83), .O(gate13inter4));
  nand2 gate1126(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1127(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1128(.a(G9), .O(gate13inter7));
  inv1  gate1129(.a(G10), .O(gate13inter8));
  nand2 gate1130(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1131(.a(s_83), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1132(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1133(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1134(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1317(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1318(.a(gate15inter0), .b(s_110), .O(gate15inter1));
  and2  gate1319(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1320(.a(s_110), .O(gate15inter3));
  inv1  gate1321(.a(s_111), .O(gate15inter4));
  nand2 gate1322(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1323(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1324(.a(G13), .O(gate15inter7));
  inv1  gate1325(.a(G14), .O(gate15inter8));
  nand2 gate1326(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1327(.a(s_111), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1328(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1329(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1330(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2563(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2564(.a(gate17inter0), .b(s_288), .O(gate17inter1));
  and2  gate2565(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2566(.a(s_288), .O(gate17inter3));
  inv1  gate2567(.a(s_289), .O(gate17inter4));
  nand2 gate2568(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2569(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2570(.a(G17), .O(gate17inter7));
  inv1  gate2571(.a(G18), .O(gate17inter8));
  nand2 gate2572(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2573(.a(s_289), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2574(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2575(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2576(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate3193(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate3194(.a(gate18inter0), .b(s_378), .O(gate18inter1));
  and2  gate3195(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate3196(.a(s_378), .O(gate18inter3));
  inv1  gate3197(.a(s_379), .O(gate18inter4));
  nand2 gate3198(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate3199(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate3200(.a(G19), .O(gate18inter7));
  inv1  gate3201(.a(G20), .O(gate18inter8));
  nand2 gate3202(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate3203(.a(s_379), .b(gate18inter3), .O(gate18inter10));
  nor2  gate3204(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate3205(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate3206(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1947(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1948(.a(gate20inter0), .b(s_200), .O(gate20inter1));
  and2  gate1949(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1950(.a(s_200), .O(gate20inter3));
  inv1  gate1951(.a(s_201), .O(gate20inter4));
  nand2 gate1952(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1953(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1954(.a(G23), .O(gate20inter7));
  inv1  gate1955(.a(G24), .O(gate20inter8));
  nand2 gate1956(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1957(.a(s_201), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1958(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1959(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1960(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2815(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2816(.a(gate22inter0), .b(s_324), .O(gate22inter1));
  and2  gate2817(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2818(.a(s_324), .O(gate22inter3));
  inv1  gate2819(.a(s_325), .O(gate22inter4));
  nand2 gate2820(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2821(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2822(.a(G27), .O(gate22inter7));
  inv1  gate2823(.a(G28), .O(gate22inter8));
  nand2 gate2824(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2825(.a(s_325), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2826(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2827(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2828(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate547(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate548(.a(gate27inter0), .b(s_0), .O(gate27inter1));
  and2  gate549(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate550(.a(s_0), .O(gate27inter3));
  inv1  gate551(.a(s_1), .O(gate27inter4));
  nand2 gate552(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate553(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate554(.a(G2), .O(gate27inter7));
  inv1  gate555(.a(G6), .O(gate27inter8));
  nand2 gate556(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate557(.a(s_1), .b(gate27inter3), .O(gate27inter10));
  nor2  gate558(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate559(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate560(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1233(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1234(.a(gate31inter0), .b(s_98), .O(gate31inter1));
  and2  gate1235(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1236(.a(s_98), .O(gate31inter3));
  inv1  gate1237(.a(s_99), .O(gate31inter4));
  nand2 gate1238(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1239(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1240(.a(G4), .O(gate31inter7));
  inv1  gate1241(.a(G8), .O(gate31inter8));
  nand2 gate1242(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1243(.a(s_99), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1244(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1245(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1246(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate771(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate772(.a(gate40inter0), .b(s_32), .O(gate40inter1));
  and2  gate773(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate774(.a(s_32), .O(gate40inter3));
  inv1  gate775(.a(s_33), .O(gate40inter4));
  nand2 gate776(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate777(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate778(.a(G28), .O(gate40inter7));
  inv1  gate779(.a(G32), .O(gate40inter8));
  nand2 gate780(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate781(.a(s_33), .b(gate40inter3), .O(gate40inter10));
  nor2  gate782(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate783(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate784(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2955(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2956(.a(gate41inter0), .b(s_344), .O(gate41inter1));
  and2  gate2957(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2958(.a(s_344), .O(gate41inter3));
  inv1  gate2959(.a(s_345), .O(gate41inter4));
  nand2 gate2960(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2961(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2962(.a(G1), .O(gate41inter7));
  inv1  gate2963(.a(G266), .O(gate41inter8));
  nand2 gate2964(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2965(.a(s_345), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2966(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2967(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2968(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1429(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1430(.a(gate44inter0), .b(s_126), .O(gate44inter1));
  and2  gate1431(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1432(.a(s_126), .O(gate44inter3));
  inv1  gate1433(.a(s_127), .O(gate44inter4));
  nand2 gate1434(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1435(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1436(.a(G4), .O(gate44inter7));
  inv1  gate1437(.a(G269), .O(gate44inter8));
  nand2 gate1438(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1439(.a(s_127), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1440(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1441(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1442(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1107(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1108(.a(gate46inter0), .b(s_80), .O(gate46inter1));
  and2  gate1109(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1110(.a(s_80), .O(gate46inter3));
  inv1  gate1111(.a(s_81), .O(gate46inter4));
  nand2 gate1112(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1113(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1114(.a(G6), .O(gate46inter7));
  inv1  gate1115(.a(G272), .O(gate46inter8));
  nand2 gate1116(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1117(.a(s_81), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1118(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1119(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1120(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1415(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1416(.a(gate47inter0), .b(s_124), .O(gate47inter1));
  and2  gate1417(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1418(.a(s_124), .O(gate47inter3));
  inv1  gate1419(.a(s_125), .O(gate47inter4));
  nand2 gate1420(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1421(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1422(.a(G7), .O(gate47inter7));
  inv1  gate1423(.a(G275), .O(gate47inter8));
  nand2 gate1424(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1425(.a(s_125), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1426(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1427(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1428(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2521(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2522(.a(gate48inter0), .b(s_282), .O(gate48inter1));
  and2  gate2523(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2524(.a(s_282), .O(gate48inter3));
  inv1  gate2525(.a(s_283), .O(gate48inter4));
  nand2 gate2526(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2527(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2528(.a(G8), .O(gate48inter7));
  inv1  gate2529(.a(G275), .O(gate48inter8));
  nand2 gate2530(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2531(.a(s_283), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2532(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2533(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2534(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate757(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate758(.a(gate49inter0), .b(s_30), .O(gate49inter1));
  and2  gate759(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate760(.a(s_30), .O(gate49inter3));
  inv1  gate761(.a(s_31), .O(gate49inter4));
  nand2 gate762(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate763(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate764(.a(G9), .O(gate49inter7));
  inv1  gate765(.a(G278), .O(gate49inter8));
  nand2 gate766(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate767(.a(s_31), .b(gate49inter3), .O(gate49inter10));
  nor2  gate768(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate769(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate770(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2367(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2368(.a(gate50inter0), .b(s_260), .O(gate50inter1));
  and2  gate2369(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2370(.a(s_260), .O(gate50inter3));
  inv1  gate2371(.a(s_261), .O(gate50inter4));
  nand2 gate2372(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2373(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2374(.a(G10), .O(gate50inter7));
  inv1  gate2375(.a(G278), .O(gate50inter8));
  nand2 gate2376(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2377(.a(s_261), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2378(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2379(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2380(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2675(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2676(.a(gate52inter0), .b(s_304), .O(gate52inter1));
  and2  gate2677(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2678(.a(s_304), .O(gate52inter3));
  inv1  gate2679(.a(s_305), .O(gate52inter4));
  nand2 gate2680(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2681(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2682(.a(G12), .O(gate52inter7));
  inv1  gate2683(.a(G281), .O(gate52inter8));
  nand2 gate2684(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2685(.a(s_305), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2686(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2687(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2688(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate2269(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2270(.a(gate53inter0), .b(s_246), .O(gate53inter1));
  and2  gate2271(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2272(.a(s_246), .O(gate53inter3));
  inv1  gate2273(.a(s_247), .O(gate53inter4));
  nand2 gate2274(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2275(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2276(.a(G13), .O(gate53inter7));
  inv1  gate2277(.a(G284), .O(gate53inter8));
  nand2 gate2278(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2279(.a(s_247), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2280(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2281(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2282(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1765(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1766(.a(gate54inter0), .b(s_174), .O(gate54inter1));
  and2  gate1767(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1768(.a(s_174), .O(gate54inter3));
  inv1  gate1769(.a(s_175), .O(gate54inter4));
  nand2 gate1770(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1771(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1772(.a(G14), .O(gate54inter7));
  inv1  gate1773(.a(G284), .O(gate54inter8));
  nand2 gate1774(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1775(.a(s_175), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1776(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1777(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1778(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate3151(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate3152(.a(gate55inter0), .b(s_372), .O(gate55inter1));
  and2  gate3153(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate3154(.a(s_372), .O(gate55inter3));
  inv1  gate3155(.a(s_373), .O(gate55inter4));
  nand2 gate3156(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate3157(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate3158(.a(G15), .O(gate55inter7));
  inv1  gate3159(.a(G287), .O(gate55inter8));
  nand2 gate3160(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate3161(.a(s_373), .b(gate55inter3), .O(gate55inter10));
  nor2  gate3162(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate3163(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate3164(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate939(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate940(.a(gate56inter0), .b(s_56), .O(gate56inter1));
  and2  gate941(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate942(.a(s_56), .O(gate56inter3));
  inv1  gate943(.a(s_57), .O(gate56inter4));
  nand2 gate944(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate945(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate946(.a(G16), .O(gate56inter7));
  inv1  gate947(.a(G287), .O(gate56inter8));
  nand2 gate948(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate949(.a(s_57), .b(gate56inter3), .O(gate56inter10));
  nor2  gate950(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate951(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate952(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate2199(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2200(.a(gate57inter0), .b(s_236), .O(gate57inter1));
  and2  gate2201(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2202(.a(s_236), .O(gate57inter3));
  inv1  gate2203(.a(s_237), .O(gate57inter4));
  nand2 gate2204(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2205(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2206(.a(G17), .O(gate57inter7));
  inv1  gate2207(.a(G290), .O(gate57inter8));
  nand2 gate2208(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2209(.a(s_237), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2210(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2211(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2212(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2381(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2382(.a(gate62inter0), .b(s_262), .O(gate62inter1));
  and2  gate2383(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2384(.a(s_262), .O(gate62inter3));
  inv1  gate2385(.a(s_263), .O(gate62inter4));
  nand2 gate2386(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2387(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2388(.a(G22), .O(gate62inter7));
  inv1  gate2389(.a(G296), .O(gate62inter8));
  nand2 gate2390(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2391(.a(s_263), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2392(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2393(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2394(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate3179(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate3180(.a(gate64inter0), .b(s_376), .O(gate64inter1));
  and2  gate3181(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate3182(.a(s_376), .O(gate64inter3));
  inv1  gate3183(.a(s_377), .O(gate64inter4));
  nand2 gate3184(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate3185(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate3186(.a(G24), .O(gate64inter7));
  inv1  gate3187(.a(G299), .O(gate64inter8));
  nand2 gate3188(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate3189(.a(s_377), .b(gate64inter3), .O(gate64inter10));
  nor2  gate3190(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate3191(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate3192(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2647(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2648(.a(gate67inter0), .b(s_300), .O(gate67inter1));
  and2  gate2649(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2650(.a(s_300), .O(gate67inter3));
  inv1  gate2651(.a(s_301), .O(gate67inter4));
  nand2 gate2652(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2653(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2654(.a(G27), .O(gate67inter7));
  inv1  gate2655(.a(G305), .O(gate67inter8));
  nand2 gate2656(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2657(.a(s_301), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2658(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2659(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2660(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate3137(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate3138(.a(gate68inter0), .b(s_370), .O(gate68inter1));
  and2  gate3139(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate3140(.a(s_370), .O(gate68inter3));
  inv1  gate3141(.a(s_371), .O(gate68inter4));
  nand2 gate3142(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate3143(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate3144(.a(G28), .O(gate68inter7));
  inv1  gate3145(.a(G305), .O(gate68inter8));
  nand2 gate3146(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate3147(.a(s_371), .b(gate68inter3), .O(gate68inter10));
  nor2  gate3148(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate3149(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate3150(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate2899(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2900(.a(gate69inter0), .b(s_336), .O(gate69inter1));
  and2  gate2901(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2902(.a(s_336), .O(gate69inter3));
  inv1  gate2903(.a(s_337), .O(gate69inter4));
  nand2 gate2904(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2905(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2906(.a(G29), .O(gate69inter7));
  inv1  gate2907(.a(G308), .O(gate69inter8));
  nand2 gate2908(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2909(.a(s_337), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2910(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2911(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2912(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate897(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate898(.a(gate70inter0), .b(s_50), .O(gate70inter1));
  and2  gate899(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate900(.a(s_50), .O(gate70inter3));
  inv1  gate901(.a(s_51), .O(gate70inter4));
  nand2 gate902(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate903(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate904(.a(G30), .O(gate70inter7));
  inv1  gate905(.a(G308), .O(gate70inter8));
  nand2 gate906(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate907(.a(s_51), .b(gate70inter3), .O(gate70inter10));
  nor2  gate908(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate909(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate910(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1779(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1780(.a(gate74inter0), .b(s_176), .O(gate74inter1));
  and2  gate1781(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1782(.a(s_176), .O(gate74inter3));
  inv1  gate1783(.a(s_177), .O(gate74inter4));
  nand2 gate1784(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1785(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1786(.a(G5), .O(gate74inter7));
  inv1  gate1787(.a(G314), .O(gate74inter8));
  nand2 gate1788(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1789(.a(s_177), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1790(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1791(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1792(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1919(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1920(.a(gate76inter0), .b(s_196), .O(gate76inter1));
  and2  gate1921(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1922(.a(s_196), .O(gate76inter3));
  inv1  gate1923(.a(s_197), .O(gate76inter4));
  nand2 gate1924(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1925(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1926(.a(G13), .O(gate76inter7));
  inv1  gate1927(.a(G317), .O(gate76inter8));
  nand2 gate1928(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1929(.a(s_197), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1930(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1931(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1932(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1695(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1696(.a(gate80inter0), .b(s_164), .O(gate80inter1));
  and2  gate1697(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1698(.a(s_164), .O(gate80inter3));
  inv1  gate1699(.a(s_165), .O(gate80inter4));
  nand2 gate1700(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1701(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1702(.a(G14), .O(gate80inter7));
  inv1  gate1703(.a(G323), .O(gate80inter8));
  nand2 gate1704(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1705(.a(s_165), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1706(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1707(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1708(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2185(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2186(.a(gate82inter0), .b(s_234), .O(gate82inter1));
  and2  gate2187(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2188(.a(s_234), .O(gate82inter3));
  inv1  gate2189(.a(s_235), .O(gate82inter4));
  nand2 gate2190(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2191(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2192(.a(G7), .O(gate82inter7));
  inv1  gate2193(.a(G326), .O(gate82inter8));
  nand2 gate2194(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2195(.a(s_235), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2196(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2197(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2198(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1191(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1192(.a(gate83inter0), .b(s_92), .O(gate83inter1));
  and2  gate1193(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1194(.a(s_92), .O(gate83inter3));
  inv1  gate1195(.a(s_93), .O(gate83inter4));
  nand2 gate1196(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1197(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1198(.a(G11), .O(gate83inter7));
  inv1  gate1199(.a(G329), .O(gate83inter8));
  nand2 gate1200(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1201(.a(s_93), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1202(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1203(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1204(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1989(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1990(.a(gate90inter0), .b(s_206), .O(gate90inter1));
  and2  gate1991(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1992(.a(s_206), .O(gate90inter3));
  inv1  gate1993(.a(s_207), .O(gate90inter4));
  nand2 gate1994(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1995(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1996(.a(G21), .O(gate90inter7));
  inv1  gate1997(.a(G338), .O(gate90inter8));
  nand2 gate1998(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1999(.a(s_207), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2000(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2001(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2002(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2115(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2116(.a(gate91inter0), .b(s_224), .O(gate91inter1));
  and2  gate2117(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2118(.a(s_224), .O(gate91inter3));
  inv1  gate2119(.a(s_225), .O(gate91inter4));
  nand2 gate2120(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2121(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2122(.a(G25), .O(gate91inter7));
  inv1  gate2123(.a(G341), .O(gate91inter8));
  nand2 gate2124(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2125(.a(s_225), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2126(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2127(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2128(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2829(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2830(.a(gate92inter0), .b(s_326), .O(gate92inter1));
  and2  gate2831(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2832(.a(s_326), .O(gate92inter3));
  inv1  gate2833(.a(s_327), .O(gate92inter4));
  nand2 gate2834(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2835(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2836(.a(G29), .O(gate92inter7));
  inv1  gate2837(.a(G341), .O(gate92inter8));
  nand2 gate2838(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2839(.a(s_327), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2840(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2841(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2842(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate3095(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate3096(.a(gate95inter0), .b(s_364), .O(gate95inter1));
  and2  gate3097(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate3098(.a(s_364), .O(gate95inter3));
  inv1  gate3099(.a(s_365), .O(gate95inter4));
  nand2 gate3100(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate3101(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate3102(.a(G26), .O(gate95inter7));
  inv1  gate3103(.a(G347), .O(gate95inter8));
  nand2 gate3104(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate3105(.a(s_365), .b(gate95inter3), .O(gate95inter10));
  nor2  gate3106(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate3107(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate3108(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate981(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate982(.a(gate100inter0), .b(s_62), .O(gate100inter1));
  and2  gate983(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate984(.a(s_62), .O(gate100inter3));
  inv1  gate985(.a(s_63), .O(gate100inter4));
  nand2 gate986(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate987(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate988(.a(G31), .O(gate100inter7));
  inv1  gate989(.a(G353), .O(gate100inter8));
  nand2 gate990(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate991(.a(s_63), .b(gate100inter3), .O(gate100inter10));
  nor2  gate992(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate993(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate994(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1457(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1458(.a(gate102inter0), .b(s_130), .O(gate102inter1));
  and2  gate1459(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1460(.a(s_130), .O(gate102inter3));
  inv1  gate1461(.a(s_131), .O(gate102inter4));
  nand2 gate1462(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1463(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1464(.a(G24), .O(gate102inter7));
  inv1  gate1465(.a(G356), .O(gate102inter8));
  nand2 gate1466(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1467(.a(s_131), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1468(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1469(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1470(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2731(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2732(.a(gate104inter0), .b(s_312), .O(gate104inter1));
  and2  gate2733(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2734(.a(s_312), .O(gate104inter3));
  inv1  gate2735(.a(s_313), .O(gate104inter4));
  nand2 gate2736(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2737(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2738(.a(G32), .O(gate104inter7));
  inv1  gate2739(.a(G359), .O(gate104inter8));
  nand2 gate2740(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2741(.a(s_313), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2742(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2743(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2744(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2339(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2340(.a(gate106inter0), .b(s_256), .O(gate106inter1));
  and2  gate2341(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2342(.a(s_256), .O(gate106inter3));
  inv1  gate2343(.a(s_257), .O(gate106inter4));
  nand2 gate2344(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2345(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2346(.a(G364), .O(gate106inter7));
  inv1  gate2347(.a(G365), .O(gate106inter8));
  nand2 gate2348(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2349(.a(s_257), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2350(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2351(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2352(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2213(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2214(.a(gate107inter0), .b(s_238), .O(gate107inter1));
  and2  gate2215(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2216(.a(s_238), .O(gate107inter3));
  inv1  gate2217(.a(s_239), .O(gate107inter4));
  nand2 gate2218(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2219(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2220(.a(G366), .O(gate107inter7));
  inv1  gate2221(.a(G367), .O(gate107inter8));
  nand2 gate2222(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2223(.a(s_239), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2224(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2225(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2226(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate3081(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate3082(.a(gate108inter0), .b(s_362), .O(gate108inter1));
  and2  gate3083(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate3084(.a(s_362), .O(gate108inter3));
  inv1  gate3085(.a(s_363), .O(gate108inter4));
  nand2 gate3086(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate3087(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate3088(.a(G368), .O(gate108inter7));
  inv1  gate3089(.a(G369), .O(gate108inter8));
  nand2 gate3090(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate3091(.a(s_363), .b(gate108inter3), .O(gate108inter10));
  nor2  gate3092(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate3093(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate3094(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1905(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1906(.a(gate110inter0), .b(s_194), .O(gate110inter1));
  and2  gate1907(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1908(.a(s_194), .O(gate110inter3));
  inv1  gate1909(.a(s_195), .O(gate110inter4));
  nand2 gate1910(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1911(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1912(.a(G372), .O(gate110inter7));
  inv1  gate1913(.a(G373), .O(gate110inter8));
  nand2 gate1914(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1915(.a(s_195), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1916(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1917(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1918(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2773(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2774(.a(gate118inter0), .b(s_318), .O(gate118inter1));
  and2  gate2775(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2776(.a(s_318), .O(gate118inter3));
  inv1  gate2777(.a(s_319), .O(gate118inter4));
  nand2 gate2778(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2779(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2780(.a(G388), .O(gate118inter7));
  inv1  gate2781(.a(G389), .O(gate118inter8));
  nand2 gate2782(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2783(.a(s_319), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2784(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2785(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2786(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2045(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2046(.a(gate119inter0), .b(s_214), .O(gate119inter1));
  and2  gate2047(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2048(.a(s_214), .O(gate119inter3));
  inv1  gate2049(.a(s_215), .O(gate119inter4));
  nand2 gate2050(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2051(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2052(.a(G390), .O(gate119inter7));
  inv1  gate2053(.a(G391), .O(gate119inter8));
  nand2 gate2054(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2055(.a(s_215), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2056(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2057(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2058(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2241(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2242(.a(gate122inter0), .b(s_242), .O(gate122inter1));
  and2  gate2243(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2244(.a(s_242), .O(gate122inter3));
  inv1  gate2245(.a(s_243), .O(gate122inter4));
  nand2 gate2246(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2247(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2248(.a(G396), .O(gate122inter7));
  inv1  gate2249(.a(G397), .O(gate122inter8));
  nand2 gate2250(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2251(.a(s_243), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2252(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2253(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2254(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1639(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1640(.a(gate123inter0), .b(s_156), .O(gate123inter1));
  and2  gate1641(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1642(.a(s_156), .O(gate123inter3));
  inv1  gate1643(.a(s_157), .O(gate123inter4));
  nand2 gate1644(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1645(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1646(.a(G398), .O(gate123inter7));
  inv1  gate1647(.a(G399), .O(gate123inter8));
  nand2 gate1648(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1649(.a(s_157), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1650(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1651(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1652(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2437(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2438(.a(gate125inter0), .b(s_270), .O(gate125inter1));
  and2  gate2439(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2440(.a(s_270), .O(gate125inter3));
  inv1  gate2441(.a(s_271), .O(gate125inter4));
  nand2 gate2442(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2443(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2444(.a(G402), .O(gate125inter7));
  inv1  gate2445(.a(G403), .O(gate125inter8));
  nand2 gate2446(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2447(.a(s_271), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2448(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2449(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2450(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1219(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1220(.a(gate128inter0), .b(s_96), .O(gate128inter1));
  and2  gate1221(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1222(.a(s_96), .O(gate128inter3));
  inv1  gate1223(.a(s_97), .O(gate128inter4));
  nand2 gate1224(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1225(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1226(.a(G408), .O(gate128inter7));
  inv1  gate1227(.a(G409), .O(gate128inter8));
  nand2 gate1228(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1229(.a(s_97), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1230(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1231(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1232(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate575(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate576(.a(gate132inter0), .b(s_4), .O(gate132inter1));
  and2  gate577(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate578(.a(s_4), .O(gate132inter3));
  inv1  gate579(.a(s_5), .O(gate132inter4));
  nand2 gate580(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate581(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate582(.a(G416), .O(gate132inter7));
  inv1  gate583(.a(G417), .O(gate132inter8));
  nand2 gate584(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate585(.a(s_5), .b(gate132inter3), .O(gate132inter10));
  nor2  gate586(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate587(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate588(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2353(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2354(.a(gate133inter0), .b(s_258), .O(gate133inter1));
  and2  gate2355(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2356(.a(s_258), .O(gate133inter3));
  inv1  gate2357(.a(s_259), .O(gate133inter4));
  nand2 gate2358(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2359(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2360(.a(G418), .O(gate133inter7));
  inv1  gate2361(.a(G419), .O(gate133inter8));
  nand2 gate2362(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2363(.a(s_259), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2364(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2365(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2366(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1975(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1976(.a(gate135inter0), .b(s_204), .O(gate135inter1));
  and2  gate1977(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1978(.a(s_204), .O(gate135inter3));
  inv1  gate1979(.a(s_205), .O(gate135inter4));
  nand2 gate1980(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1981(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1982(.a(G422), .O(gate135inter7));
  inv1  gate1983(.a(G423), .O(gate135inter8));
  nand2 gate1984(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1985(.a(s_205), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1986(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1987(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1988(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1653(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1654(.a(gate136inter0), .b(s_158), .O(gate136inter1));
  and2  gate1655(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1656(.a(s_158), .O(gate136inter3));
  inv1  gate1657(.a(s_159), .O(gate136inter4));
  nand2 gate1658(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1659(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1660(.a(G424), .O(gate136inter7));
  inv1  gate1661(.a(G425), .O(gate136inter8));
  nand2 gate1662(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1663(.a(s_159), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1664(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1665(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1666(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1205(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1206(.a(gate137inter0), .b(s_94), .O(gate137inter1));
  and2  gate1207(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1208(.a(s_94), .O(gate137inter3));
  inv1  gate1209(.a(s_95), .O(gate137inter4));
  nand2 gate1210(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1211(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1212(.a(G426), .O(gate137inter7));
  inv1  gate1213(.a(G429), .O(gate137inter8));
  nand2 gate1214(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1215(.a(s_95), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1216(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1217(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1218(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1667(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1668(.a(gate138inter0), .b(s_160), .O(gate138inter1));
  and2  gate1669(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1670(.a(s_160), .O(gate138inter3));
  inv1  gate1671(.a(s_161), .O(gate138inter4));
  nand2 gate1672(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1673(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1674(.a(G432), .O(gate138inter7));
  inv1  gate1675(.a(G435), .O(gate138inter8));
  nand2 gate1676(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1677(.a(s_161), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1678(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1679(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1680(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2591(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2592(.a(gate141inter0), .b(s_292), .O(gate141inter1));
  and2  gate2593(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2594(.a(s_292), .O(gate141inter3));
  inv1  gate2595(.a(s_293), .O(gate141inter4));
  nand2 gate2596(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2597(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2598(.a(G450), .O(gate141inter7));
  inv1  gate2599(.a(G453), .O(gate141inter8));
  nand2 gate2600(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2601(.a(s_293), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2602(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2603(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2604(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate2913(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2914(.a(gate142inter0), .b(s_338), .O(gate142inter1));
  and2  gate2915(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2916(.a(s_338), .O(gate142inter3));
  inv1  gate2917(.a(s_339), .O(gate142inter4));
  nand2 gate2918(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2919(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2920(.a(G456), .O(gate142inter7));
  inv1  gate2921(.a(G459), .O(gate142inter8));
  nand2 gate2922(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2923(.a(s_339), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2924(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2925(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2926(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1835(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1836(.a(gate143inter0), .b(s_184), .O(gate143inter1));
  and2  gate1837(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1838(.a(s_184), .O(gate143inter3));
  inv1  gate1839(.a(s_185), .O(gate143inter4));
  nand2 gate1840(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1841(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1842(.a(G462), .O(gate143inter7));
  inv1  gate1843(.a(G465), .O(gate143inter8));
  nand2 gate1844(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1845(.a(s_185), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1846(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1847(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1848(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1681(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1682(.a(gate144inter0), .b(s_162), .O(gate144inter1));
  and2  gate1683(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1684(.a(s_162), .O(gate144inter3));
  inv1  gate1685(.a(s_163), .O(gate144inter4));
  nand2 gate1686(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1687(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1688(.a(G468), .O(gate144inter7));
  inv1  gate1689(.a(G471), .O(gate144inter8));
  nand2 gate1690(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1691(.a(s_163), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1692(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1693(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1694(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2535(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2536(.a(gate145inter0), .b(s_284), .O(gate145inter1));
  and2  gate2537(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2538(.a(s_284), .O(gate145inter3));
  inv1  gate2539(.a(s_285), .O(gate145inter4));
  nand2 gate2540(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2541(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2542(.a(G474), .O(gate145inter7));
  inv1  gate2543(.a(G477), .O(gate145inter8));
  nand2 gate2544(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2545(.a(s_285), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2546(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2547(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2548(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate3109(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate3110(.a(gate147inter0), .b(s_366), .O(gate147inter1));
  and2  gate3111(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate3112(.a(s_366), .O(gate147inter3));
  inv1  gate3113(.a(s_367), .O(gate147inter4));
  nand2 gate3114(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate3115(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate3116(.a(G486), .O(gate147inter7));
  inv1  gate3117(.a(G489), .O(gate147inter8));
  nand2 gate3118(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate3119(.a(s_367), .b(gate147inter3), .O(gate147inter10));
  nor2  gate3120(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate3121(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate3122(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate2661(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2662(.a(gate148inter0), .b(s_302), .O(gate148inter1));
  and2  gate2663(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2664(.a(s_302), .O(gate148inter3));
  inv1  gate2665(.a(s_303), .O(gate148inter4));
  nand2 gate2666(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2667(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2668(.a(G492), .O(gate148inter7));
  inv1  gate2669(.a(G495), .O(gate148inter8));
  nand2 gate2670(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2671(.a(s_303), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2672(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2673(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2674(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate701(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate702(.a(gate149inter0), .b(s_22), .O(gate149inter1));
  and2  gate703(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate704(.a(s_22), .O(gate149inter3));
  inv1  gate705(.a(s_23), .O(gate149inter4));
  nand2 gate706(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate707(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate708(.a(G498), .O(gate149inter7));
  inv1  gate709(.a(G501), .O(gate149inter8));
  nand2 gate710(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate711(.a(s_23), .b(gate149inter3), .O(gate149inter10));
  nor2  gate712(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate713(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate714(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2983(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2984(.a(gate150inter0), .b(s_348), .O(gate150inter1));
  and2  gate2985(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2986(.a(s_348), .O(gate150inter3));
  inv1  gate2987(.a(s_349), .O(gate150inter4));
  nand2 gate2988(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2989(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2990(.a(G504), .O(gate150inter7));
  inv1  gate2991(.a(G507), .O(gate150inter8));
  nand2 gate2992(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2993(.a(s_349), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2994(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2995(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2996(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1709(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1710(.a(gate151inter0), .b(s_166), .O(gate151inter1));
  and2  gate1711(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1712(.a(s_166), .O(gate151inter3));
  inv1  gate1713(.a(s_167), .O(gate151inter4));
  nand2 gate1714(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1715(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1716(.a(G510), .O(gate151inter7));
  inv1  gate1717(.a(G513), .O(gate151inter8));
  nand2 gate1718(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1719(.a(s_167), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1720(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1721(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1722(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2577(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2578(.a(gate154inter0), .b(s_290), .O(gate154inter1));
  and2  gate2579(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2580(.a(s_290), .O(gate154inter3));
  inv1  gate2581(.a(s_291), .O(gate154inter4));
  nand2 gate2582(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2583(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2584(.a(G429), .O(gate154inter7));
  inv1  gate2585(.a(G522), .O(gate154inter8));
  nand2 gate2586(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2587(.a(s_291), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2588(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2589(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2590(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate855(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate856(.a(gate157inter0), .b(s_44), .O(gate157inter1));
  and2  gate857(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate858(.a(s_44), .O(gate157inter3));
  inv1  gate859(.a(s_45), .O(gate157inter4));
  nand2 gate860(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate861(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate862(.a(G438), .O(gate157inter7));
  inv1  gate863(.a(G528), .O(gate157inter8));
  nand2 gate864(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate865(.a(s_45), .b(gate157inter3), .O(gate157inter10));
  nor2  gate866(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate867(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate868(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1163(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1164(.a(gate159inter0), .b(s_88), .O(gate159inter1));
  and2  gate1165(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1166(.a(s_88), .O(gate159inter3));
  inv1  gate1167(.a(s_89), .O(gate159inter4));
  nand2 gate1168(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1169(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1170(.a(G444), .O(gate159inter7));
  inv1  gate1171(.a(G531), .O(gate159inter8));
  nand2 gate1172(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1173(.a(s_89), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1174(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1175(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1176(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2395(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2396(.a(gate160inter0), .b(s_264), .O(gate160inter1));
  and2  gate2397(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2398(.a(s_264), .O(gate160inter3));
  inv1  gate2399(.a(s_265), .O(gate160inter4));
  nand2 gate2400(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2401(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2402(.a(G447), .O(gate160inter7));
  inv1  gate2403(.a(G531), .O(gate160inter8));
  nand2 gate2404(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2405(.a(s_265), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2406(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2407(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2408(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate799(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate800(.a(gate165inter0), .b(s_36), .O(gate165inter1));
  and2  gate801(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate802(.a(s_36), .O(gate165inter3));
  inv1  gate803(.a(s_37), .O(gate165inter4));
  nand2 gate804(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate805(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate806(.a(G462), .O(gate165inter7));
  inv1  gate807(.a(G540), .O(gate165inter8));
  nand2 gate808(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate809(.a(s_37), .b(gate165inter3), .O(gate165inter10));
  nor2  gate810(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate811(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate812(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1177(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1178(.a(gate166inter0), .b(s_90), .O(gate166inter1));
  and2  gate1179(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1180(.a(s_90), .O(gate166inter3));
  inv1  gate1181(.a(s_91), .O(gate166inter4));
  nand2 gate1182(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1183(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1184(.a(G465), .O(gate166inter7));
  inv1  gate1185(.a(G540), .O(gate166inter8));
  nand2 gate1186(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1187(.a(s_91), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1188(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1189(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1190(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2507(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2508(.a(gate167inter0), .b(s_280), .O(gate167inter1));
  and2  gate2509(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2510(.a(s_280), .O(gate167inter3));
  inv1  gate2511(.a(s_281), .O(gate167inter4));
  nand2 gate2512(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2513(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2514(.a(G468), .O(gate167inter7));
  inv1  gate2515(.a(G543), .O(gate167inter8));
  nand2 gate2516(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2517(.a(s_281), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2518(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2519(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2520(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1597(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1598(.a(gate169inter0), .b(s_150), .O(gate169inter1));
  and2  gate1599(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1600(.a(s_150), .O(gate169inter3));
  inv1  gate1601(.a(s_151), .O(gate169inter4));
  nand2 gate1602(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1603(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1604(.a(G474), .O(gate169inter7));
  inv1  gate1605(.a(G546), .O(gate169inter8));
  nand2 gate1606(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1607(.a(s_151), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1608(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1609(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1610(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate645(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate646(.a(gate171inter0), .b(s_14), .O(gate171inter1));
  and2  gate647(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate648(.a(s_14), .O(gate171inter3));
  inv1  gate649(.a(s_15), .O(gate171inter4));
  nand2 gate650(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate651(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate652(.a(G480), .O(gate171inter7));
  inv1  gate653(.a(G549), .O(gate171inter8));
  nand2 gate654(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate655(.a(s_15), .b(gate171inter3), .O(gate171inter10));
  nor2  gate656(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate657(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate658(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate729(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate730(.a(gate172inter0), .b(s_26), .O(gate172inter1));
  and2  gate731(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate732(.a(s_26), .O(gate172inter3));
  inv1  gate733(.a(s_27), .O(gate172inter4));
  nand2 gate734(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate735(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate736(.a(G483), .O(gate172inter7));
  inv1  gate737(.a(G549), .O(gate172inter8));
  nand2 gate738(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate739(.a(s_27), .b(gate172inter3), .O(gate172inter10));
  nor2  gate740(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate741(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate742(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1877(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1878(.a(gate173inter0), .b(s_190), .O(gate173inter1));
  and2  gate1879(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1880(.a(s_190), .O(gate173inter3));
  inv1  gate1881(.a(s_191), .O(gate173inter4));
  nand2 gate1882(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1883(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1884(.a(G486), .O(gate173inter7));
  inv1  gate1885(.a(G552), .O(gate173inter8));
  nand2 gate1886(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1887(.a(s_191), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1888(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1889(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1890(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2059(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2060(.a(gate174inter0), .b(s_216), .O(gate174inter1));
  and2  gate2061(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2062(.a(s_216), .O(gate174inter3));
  inv1  gate2063(.a(s_217), .O(gate174inter4));
  nand2 gate2064(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2065(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2066(.a(G489), .O(gate174inter7));
  inv1  gate2067(.a(G552), .O(gate174inter8));
  nand2 gate2068(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2069(.a(s_217), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2070(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2071(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2072(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1849(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1850(.a(gate175inter0), .b(s_186), .O(gate175inter1));
  and2  gate1851(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1852(.a(s_186), .O(gate175inter3));
  inv1  gate1853(.a(s_187), .O(gate175inter4));
  nand2 gate1854(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1855(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1856(.a(G492), .O(gate175inter7));
  inv1  gate1857(.a(G555), .O(gate175inter8));
  nand2 gate1858(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1859(.a(s_187), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1860(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1861(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1862(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1527(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1528(.a(gate177inter0), .b(s_140), .O(gate177inter1));
  and2  gate1529(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1530(.a(s_140), .O(gate177inter3));
  inv1  gate1531(.a(s_141), .O(gate177inter4));
  nand2 gate1532(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1533(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1534(.a(G498), .O(gate177inter7));
  inv1  gate1535(.a(G558), .O(gate177inter8));
  nand2 gate1536(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1537(.a(s_141), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1538(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1539(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1540(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2969(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2970(.a(gate181inter0), .b(s_346), .O(gate181inter1));
  and2  gate2971(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2972(.a(s_346), .O(gate181inter3));
  inv1  gate2973(.a(s_347), .O(gate181inter4));
  nand2 gate2974(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2975(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2976(.a(G510), .O(gate181inter7));
  inv1  gate2977(.a(G564), .O(gate181inter8));
  nand2 gate2978(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2979(.a(s_347), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2980(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2981(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2982(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2227(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2228(.a(gate184inter0), .b(s_240), .O(gate184inter1));
  and2  gate2229(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2230(.a(s_240), .O(gate184inter3));
  inv1  gate2231(.a(s_241), .O(gate184inter4));
  nand2 gate2232(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2233(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2234(.a(G519), .O(gate184inter7));
  inv1  gate2235(.a(G567), .O(gate184inter8));
  nand2 gate2236(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2237(.a(s_241), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2238(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2239(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2240(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2689(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2690(.a(gate185inter0), .b(s_306), .O(gate185inter1));
  and2  gate2691(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2692(.a(s_306), .O(gate185inter3));
  inv1  gate2693(.a(s_307), .O(gate185inter4));
  nand2 gate2694(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2695(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2696(.a(G570), .O(gate185inter7));
  inv1  gate2697(.a(G571), .O(gate185inter8));
  nand2 gate2698(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2699(.a(s_307), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2700(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2701(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2702(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1303(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1304(.a(gate189inter0), .b(s_108), .O(gate189inter1));
  and2  gate1305(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1306(.a(s_108), .O(gate189inter3));
  inv1  gate1307(.a(s_109), .O(gate189inter4));
  nand2 gate1308(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1309(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1310(.a(G578), .O(gate189inter7));
  inv1  gate1311(.a(G579), .O(gate189inter8));
  nand2 gate1312(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1313(.a(s_109), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1314(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1315(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1316(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1583(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1584(.a(gate190inter0), .b(s_148), .O(gate190inter1));
  and2  gate1585(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1586(.a(s_148), .O(gate190inter3));
  inv1  gate1587(.a(s_149), .O(gate190inter4));
  nand2 gate1588(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1589(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1590(.a(G580), .O(gate190inter7));
  inv1  gate1591(.a(G581), .O(gate190inter8));
  nand2 gate1592(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1593(.a(s_149), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1594(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1595(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1596(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1289(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1290(.a(gate192inter0), .b(s_106), .O(gate192inter1));
  and2  gate1291(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1292(.a(s_106), .O(gate192inter3));
  inv1  gate1293(.a(s_107), .O(gate192inter4));
  nand2 gate1294(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1295(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1296(.a(G584), .O(gate192inter7));
  inv1  gate1297(.a(G585), .O(gate192inter8));
  nand2 gate1298(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1299(.a(s_107), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1300(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1301(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1302(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate2787(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2788(.a(gate196inter0), .b(s_320), .O(gate196inter1));
  and2  gate2789(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2790(.a(s_320), .O(gate196inter3));
  inv1  gate2791(.a(s_321), .O(gate196inter4));
  nand2 gate2792(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2793(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2794(.a(G592), .O(gate196inter7));
  inv1  gate2795(.a(G593), .O(gate196inter8));
  nand2 gate2796(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2797(.a(s_321), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2798(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2799(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2800(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1079(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1080(.a(gate198inter0), .b(s_76), .O(gate198inter1));
  and2  gate1081(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1082(.a(s_76), .O(gate198inter3));
  inv1  gate1083(.a(s_77), .O(gate198inter4));
  nand2 gate1084(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1085(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1086(.a(G596), .O(gate198inter7));
  inv1  gate1087(.a(G597), .O(gate198inter8));
  nand2 gate1088(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1089(.a(s_77), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1090(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1091(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1092(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1359(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1360(.a(gate199inter0), .b(s_116), .O(gate199inter1));
  and2  gate1361(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1362(.a(s_116), .O(gate199inter3));
  inv1  gate1363(.a(s_117), .O(gate199inter4));
  nand2 gate1364(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1365(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1366(.a(G598), .O(gate199inter7));
  inv1  gate1367(.a(G599), .O(gate199inter8));
  nand2 gate1368(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1369(.a(s_117), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1370(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1371(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1372(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate2885(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2886(.a(gate200inter0), .b(s_334), .O(gate200inter1));
  and2  gate2887(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2888(.a(s_334), .O(gate200inter3));
  inv1  gate2889(.a(s_335), .O(gate200inter4));
  nand2 gate2890(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2891(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2892(.a(G600), .O(gate200inter7));
  inv1  gate2893(.a(G601), .O(gate200inter8));
  nand2 gate2894(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2895(.a(s_335), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2896(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2897(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2898(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2451(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2452(.a(gate202inter0), .b(s_272), .O(gate202inter1));
  and2  gate2453(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2454(.a(s_272), .O(gate202inter3));
  inv1  gate2455(.a(s_273), .O(gate202inter4));
  nand2 gate2456(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2457(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2458(.a(G612), .O(gate202inter7));
  inv1  gate2459(.a(G617), .O(gate202inter8));
  nand2 gate2460(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2461(.a(s_273), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2462(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2463(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2464(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1737(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1738(.a(gate203inter0), .b(s_170), .O(gate203inter1));
  and2  gate1739(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1740(.a(s_170), .O(gate203inter3));
  inv1  gate1741(.a(s_171), .O(gate203inter4));
  nand2 gate1742(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1743(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1744(.a(G602), .O(gate203inter7));
  inv1  gate1745(.a(G612), .O(gate203inter8));
  nand2 gate1746(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1747(.a(s_171), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1748(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1749(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1750(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2087(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2088(.a(gate208inter0), .b(s_220), .O(gate208inter1));
  and2  gate2089(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2090(.a(s_220), .O(gate208inter3));
  inv1  gate2091(.a(s_221), .O(gate208inter4));
  nand2 gate2092(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2093(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2094(.a(G627), .O(gate208inter7));
  inv1  gate2095(.a(G637), .O(gate208inter8));
  nand2 gate2096(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2097(.a(s_221), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2098(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2099(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2100(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2717(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2718(.a(gate212inter0), .b(s_310), .O(gate212inter1));
  and2  gate2719(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2720(.a(s_310), .O(gate212inter3));
  inv1  gate2721(.a(s_311), .O(gate212inter4));
  nand2 gate2722(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2723(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2724(.a(G617), .O(gate212inter7));
  inv1  gate2725(.a(G669), .O(gate212inter8));
  nand2 gate2726(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2727(.a(s_311), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2728(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2729(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2730(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1569(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1570(.a(gate217inter0), .b(s_146), .O(gate217inter1));
  and2  gate1571(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1572(.a(s_146), .O(gate217inter3));
  inv1  gate1573(.a(s_147), .O(gate217inter4));
  nand2 gate1574(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1575(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1576(.a(G622), .O(gate217inter7));
  inv1  gate1577(.a(G678), .O(gate217inter8));
  nand2 gate1578(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1579(.a(s_147), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1580(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1581(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1582(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1793(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1794(.a(gate218inter0), .b(s_178), .O(gate218inter1));
  and2  gate1795(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1796(.a(s_178), .O(gate218inter3));
  inv1  gate1797(.a(s_179), .O(gate218inter4));
  nand2 gate1798(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1799(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1800(.a(G627), .O(gate218inter7));
  inv1  gate1801(.a(G678), .O(gate218inter8));
  nand2 gate1802(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1803(.a(s_179), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1804(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1805(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1806(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2157(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2158(.a(gate225inter0), .b(s_230), .O(gate225inter1));
  and2  gate2159(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2160(.a(s_230), .O(gate225inter3));
  inv1  gate2161(.a(s_231), .O(gate225inter4));
  nand2 gate2162(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2163(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2164(.a(G690), .O(gate225inter7));
  inv1  gate2165(.a(G691), .O(gate225inter8));
  nand2 gate2166(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2167(.a(s_231), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2168(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2169(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2170(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate603(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate604(.a(gate226inter0), .b(s_8), .O(gate226inter1));
  and2  gate605(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate606(.a(s_8), .O(gate226inter3));
  inv1  gate607(.a(s_9), .O(gate226inter4));
  nand2 gate608(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate609(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate610(.a(G692), .O(gate226inter7));
  inv1  gate611(.a(G693), .O(gate226inter8));
  nand2 gate612(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate613(.a(s_9), .b(gate226inter3), .O(gate226inter10));
  nor2  gate614(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate615(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate616(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1387(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1388(.a(gate233inter0), .b(s_120), .O(gate233inter1));
  and2  gate1389(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1390(.a(s_120), .O(gate233inter3));
  inv1  gate1391(.a(s_121), .O(gate233inter4));
  nand2 gate1392(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1393(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1394(.a(G242), .O(gate233inter7));
  inv1  gate1395(.a(G718), .O(gate233inter8));
  nand2 gate1396(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1397(.a(s_121), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1398(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1399(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1400(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate785(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate786(.a(gate234inter0), .b(s_34), .O(gate234inter1));
  and2  gate787(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate788(.a(s_34), .O(gate234inter3));
  inv1  gate789(.a(s_35), .O(gate234inter4));
  nand2 gate790(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate791(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate792(.a(G245), .O(gate234inter7));
  inv1  gate793(.a(G721), .O(gate234inter8));
  nand2 gate794(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate795(.a(s_35), .b(gate234inter3), .O(gate234inter10));
  nor2  gate796(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate797(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate798(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate673(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate674(.a(gate242inter0), .b(s_18), .O(gate242inter1));
  and2  gate675(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate676(.a(s_18), .O(gate242inter3));
  inv1  gate677(.a(s_19), .O(gate242inter4));
  nand2 gate678(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate679(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate680(.a(G718), .O(gate242inter7));
  inv1  gate681(.a(G730), .O(gate242inter8));
  nand2 gate682(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate683(.a(s_19), .b(gate242inter3), .O(gate242inter10));
  nor2  gate684(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate685(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate686(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1961(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1962(.a(gate243inter0), .b(s_202), .O(gate243inter1));
  and2  gate1963(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1964(.a(s_202), .O(gate243inter3));
  inv1  gate1965(.a(s_203), .O(gate243inter4));
  nand2 gate1966(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1967(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1968(.a(G245), .O(gate243inter7));
  inv1  gate1969(.a(G733), .O(gate243inter8));
  nand2 gate1970(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1971(.a(s_203), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1972(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1973(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1974(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2143(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2144(.a(gate245inter0), .b(s_228), .O(gate245inter1));
  and2  gate2145(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2146(.a(s_228), .O(gate245inter3));
  inv1  gate2147(.a(s_229), .O(gate245inter4));
  nand2 gate2148(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2149(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2150(.a(G248), .O(gate245inter7));
  inv1  gate2151(.a(G736), .O(gate245inter8));
  nand2 gate2152(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2153(.a(s_229), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2154(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2155(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2156(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1471(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1472(.a(gate246inter0), .b(s_132), .O(gate246inter1));
  and2  gate1473(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1474(.a(s_132), .O(gate246inter3));
  inv1  gate1475(.a(s_133), .O(gate246inter4));
  nand2 gate1476(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1477(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1478(.a(G724), .O(gate246inter7));
  inv1  gate1479(.a(G736), .O(gate246inter8));
  nand2 gate1480(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1481(.a(s_133), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1482(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1483(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1484(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate2311(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2312(.a(gate247inter0), .b(s_252), .O(gate247inter1));
  and2  gate2313(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2314(.a(s_252), .O(gate247inter3));
  inv1  gate2315(.a(s_253), .O(gate247inter4));
  nand2 gate2316(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2317(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2318(.a(G251), .O(gate247inter7));
  inv1  gate2319(.a(G739), .O(gate247inter8));
  nand2 gate2320(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2321(.a(s_253), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2322(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2323(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2324(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2479(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2480(.a(gate248inter0), .b(s_276), .O(gate248inter1));
  and2  gate2481(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2482(.a(s_276), .O(gate248inter3));
  inv1  gate2483(.a(s_277), .O(gate248inter4));
  nand2 gate2484(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2485(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2486(.a(G727), .O(gate248inter7));
  inv1  gate2487(.a(G739), .O(gate248inter8));
  nand2 gate2488(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2489(.a(s_277), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2490(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2491(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2492(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2493(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2494(.a(gate250inter0), .b(s_278), .O(gate250inter1));
  and2  gate2495(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2496(.a(s_278), .O(gate250inter3));
  inv1  gate2497(.a(s_279), .O(gate250inter4));
  nand2 gate2498(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2499(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2500(.a(G706), .O(gate250inter7));
  inv1  gate2501(.a(G742), .O(gate250inter8));
  nand2 gate2502(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2503(.a(s_279), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2504(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2505(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2506(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1513(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1514(.a(gate253inter0), .b(s_138), .O(gate253inter1));
  and2  gate1515(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1516(.a(s_138), .O(gate253inter3));
  inv1  gate1517(.a(s_139), .O(gate253inter4));
  nand2 gate1518(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1519(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1520(.a(G260), .O(gate253inter7));
  inv1  gate1521(.a(G748), .O(gate253inter8));
  nand2 gate1522(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1523(.a(s_139), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1524(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1525(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1526(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate2423(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2424(.a(gate254inter0), .b(s_268), .O(gate254inter1));
  and2  gate2425(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2426(.a(s_268), .O(gate254inter3));
  inv1  gate2427(.a(s_269), .O(gate254inter4));
  nand2 gate2428(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2429(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2430(.a(G712), .O(gate254inter7));
  inv1  gate2431(.a(G748), .O(gate254inter8));
  nand2 gate2432(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2433(.a(s_269), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2434(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2435(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2436(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1863(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1864(.a(gate255inter0), .b(s_188), .O(gate255inter1));
  and2  gate1865(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1866(.a(s_188), .O(gate255inter3));
  inv1  gate1867(.a(s_189), .O(gate255inter4));
  nand2 gate1868(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1869(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1870(.a(G263), .O(gate255inter7));
  inv1  gate1871(.a(G751), .O(gate255inter8));
  nand2 gate1872(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1873(.a(s_189), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1874(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1875(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1876(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2633(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2634(.a(gate257inter0), .b(s_298), .O(gate257inter1));
  and2  gate2635(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2636(.a(s_298), .O(gate257inter3));
  inv1  gate2637(.a(s_299), .O(gate257inter4));
  nand2 gate2638(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2639(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2640(.a(G754), .O(gate257inter7));
  inv1  gate2641(.a(G755), .O(gate257inter8));
  nand2 gate2642(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2643(.a(s_299), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2644(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2645(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2646(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1611(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1612(.a(gate263inter0), .b(s_152), .O(gate263inter1));
  and2  gate1613(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1614(.a(s_152), .O(gate263inter3));
  inv1  gate1615(.a(s_153), .O(gate263inter4));
  nand2 gate1616(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1617(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1618(.a(G766), .O(gate263inter7));
  inv1  gate1619(.a(G767), .O(gate263inter8));
  nand2 gate1620(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1621(.a(s_153), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1622(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1623(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1624(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1093(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1094(.a(gate264inter0), .b(s_78), .O(gate264inter1));
  and2  gate1095(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1096(.a(s_78), .O(gate264inter3));
  inv1  gate1097(.a(s_79), .O(gate264inter4));
  nand2 gate1098(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1099(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1100(.a(G768), .O(gate264inter7));
  inv1  gate1101(.a(G769), .O(gate264inter8));
  nand2 gate1102(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1103(.a(s_79), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1104(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1105(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1106(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate2255(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2256(.a(gate265inter0), .b(s_244), .O(gate265inter1));
  and2  gate2257(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2258(.a(s_244), .O(gate265inter3));
  inv1  gate2259(.a(s_245), .O(gate265inter4));
  nand2 gate2260(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2261(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2262(.a(G642), .O(gate265inter7));
  inv1  gate2263(.a(G770), .O(gate265inter8));
  nand2 gate2264(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2265(.a(s_245), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2266(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2267(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2268(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate715(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate716(.a(gate270inter0), .b(s_24), .O(gate270inter1));
  and2  gate717(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate718(.a(s_24), .O(gate270inter3));
  inv1  gate719(.a(s_25), .O(gate270inter4));
  nand2 gate720(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate721(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate722(.a(G657), .O(gate270inter7));
  inv1  gate723(.a(G785), .O(gate270inter8));
  nand2 gate724(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate725(.a(s_25), .b(gate270inter3), .O(gate270inter10));
  nor2  gate726(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate727(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate728(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1275(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1276(.a(gate271inter0), .b(s_104), .O(gate271inter1));
  and2  gate1277(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1278(.a(s_104), .O(gate271inter3));
  inv1  gate1279(.a(s_105), .O(gate271inter4));
  nand2 gate1280(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1281(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1282(.a(G660), .O(gate271inter7));
  inv1  gate1283(.a(G788), .O(gate271inter8));
  nand2 gate1284(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1285(.a(s_105), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1286(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1287(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1288(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1499(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1500(.a(gate272inter0), .b(s_136), .O(gate272inter1));
  and2  gate1501(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1502(.a(s_136), .O(gate272inter3));
  inv1  gate1503(.a(s_137), .O(gate272inter4));
  nand2 gate1504(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1505(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1506(.a(G663), .O(gate272inter7));
  inv1  gate1507(.a(G791), .O(gate272inter8));
  nand2 gate1508(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1509(.a(s_137), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1510(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1511(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1512(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate3039(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate3040(.a(gate273inter0), .b(s_356), .O(gate273inter1));
  and2  gate3041(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate3042(.a(s_356), .O(gate273inter3));
  inv1  gate3043(.a(s_357), .O(gate273inter4));
  nand2 gate3044(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate3045(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate3046(.a(G642), .O(gate273inter7));
  inv1  gate3047(.a(G794), .O(gate273inter8));
  nand2 gate3048(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate3049(.a(s_357), .b(gate273inter3), .O(gate273inter10));
  nor2  gate3050(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate3051(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate3052(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1009(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1010(.a(gate274inter0), .b(s_66), .O(gate274inter1));
  and2  gate1011(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1012(.a(s_66), .O(gate274inter3));
  inv1  gate1013(.a(s_67), .O(gate274inter4));
  nand2 gate1014(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1015(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1016(.a(G770), .O(gate274inter7));
  inv1  gate1017(.a(G794), .O(gate274inter8));
  nand2 gate1018(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1019(.a(s_67), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1020(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1021(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1022(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1891(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1892(.a(gate275inter0), .b(s_192), .O(gate275inter1));
  and2  gate1893(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1894(.a(s_192), .O(gate275inter3));
  inv1  gate1895(.a(s_193), .O(gate275inter4));
  nand2 gate1896(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1897(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1898(.a(G645), .O(gate275inter7));
  inv1  gate1899(.a(G797), .O(gate275inter8));
  nand2 gate1900(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1901(.a(s_193), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1902(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1903(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1904(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate925(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate926(.a(gate278inter0), .b(s_54), .O(gate278inter1));
  and2  gate927(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate928(.a(s_54), .O(gate278inter3));
  inv1  gate929(.a(s_55), .O(gate278inter4));
  nand2 gate930(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate931(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate932(.a(G776), .O(gate278inter7));
  inv1  gate933(.a(G800), .O(gate278inter8));
  nand2 gate934(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate935(.a(s_55), .b(gate278inter3), .O(gate278inter10));
  nor2  gate936(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate937(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate938(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2297(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2298(.a(gate283inter0), .b(s_250), .O(gate283inter1));
  and2  gate2299(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2300(.a(s_250), .O(gate283inter3));
  inv1  gate2301(.a(s_251), .O(gate283inter4));
  nand2 gate2302(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2303(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2304(.a(G657), .O(gate283inter7));
  inv1  gate2305(.a(G809), .O(gate283inter8));
  nand2 gate2306(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2307(.a(s_251), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2308(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2309(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2310(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate631(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate632(.a(gate284inter0), .b(s_12), .O(gate284inter1));
  and2  gate633(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate634(.a(s_12), .O(gate284inter3));
  inv1  gate635(.a(s_13), .O(gate284inter4));
  nand2 gate636(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate637(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate638(.a(G785), .O(gate284inter7));
  inv1  gate639(.a(G809), .O(gate284inter8));
  nand2 gate640(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate641(.a(s_13), .b(gate284inter3), .O(gate284inter10));
  nor2  gate642(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate643(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate644(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2857(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2858(.a(gate285inter0), .b(s_330), .O(gate285inter1));
  and2  gate2859(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2860(.a(s_330), .O(gate285inter3));
  inv1  gate2861(.a(s_331), .O(gate285inter4));
  nand2 gate2862(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2863(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2864(.a(G660), .O(gate285inter7));
  inv1  gate2865(.a(G812), .O(gate285inter8));
  nand2 gate2866(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2867(.a(s_331), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2868(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2869(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2870(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate841(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate842(.a(gate287inter0), .b(s_42), .O(gate287inter1));
  and2  gate843(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate844(.a(s_42), .O(gate287inter3));
  inv1  gate845(.a(s_43), .O(gate287inter4));
  nand2 gate846(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate847(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate848(.a(G663), .O(gate287inter7));
  inv1  gate849(.a(G815), .O(gate287inter8));
  nand2 gate850(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate851(.a(s_43), .b(gate287inter3), .O(gate287inter10));
  nor2  gate852(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate853(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate854(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2759(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2760(.a(gate289inter0), .b(s_316), .O(gate289inter1));
  and2  gate2761(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2762(.a(s_316), .O(gate289inter3));
  inv1  gate2763(.a(s_317), .O(gate289inter4));
  nand2 gate2764(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2765(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2766(.a(G818), .O(gate289inter7));
  inv1  gate2767(.a(G819), .O(gate289inter8));
  nand2 gate2768(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2769(.a(s_317), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2770(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2771(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2772(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2031(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2032(.a(gate293inter0), .b(s_212), .O(gate293inter1));
  and2  gate2033(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2034(.a(s_212), .O(gate293inter3));
  inv1  gate2035(.a(s_213), .O(gate293inter4));
  nand2 gate2036(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2037(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2038(.a(G828), .O(gate293inter7));
  inv1  gate2039(.a(G829), .O(gate293inter8));
  nand2 gate2040(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2041(.a(s_213), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2042(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2043(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2044(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate3067(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate3068(.a(gate294inter0), .b(s_360), .O(gate294inter1));
  and2  gate3069(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate3070(.a(s_360), .O(gate294inter3));
  inv1  gate3071(.a(s_361), .O(gate294inter4));
  nand2 gate3072(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate3073(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate3074(.a(G832), .O(gate294inter7));
  inv1  gate3075(.a(G833), .O(gate294inter8));
  nand2 gate3076(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate3077(.a(s_361), .b(gate294inter3), .O(gate294inter10));
  nor2  gate3078(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate3079(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate3080(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate3123(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate3124(.a(gate387inter0), .b(s_368), .O(gate387inter1));
  and2  gate3125(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate3126(.a(s_368), .O(gate387inter3));
  inv1  gate3127(.a(s_369), .O(gate387inter4));
  nand2 gate3128(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate3129(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate3130(.a(G1), .O(gate387inter7));
  inv1  gate3131(.a(G1036), .O(gate387inter8));
  nand2 gate3132(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate3133(.a(s_369), .b(gate387inter3), .O(gate387inter10));
  nor2  gate3134(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate3135(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate3136(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1051(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1052(.a(gate389inter0), .b(s_72), .O(gate389inter1));
  and2  gate1053(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1054(.a(s_72), .O(gate389inter3));
  inv1  gate1055(.a(s_73), .O(gate389inter4));
  nand2 gate1056(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1057(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1058(.a(G3), .O(gate389inter7));
  inv1  gate1059(.a(G1042), .O(gate389inter8));
  nand2 gate1060(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1061(.a(s_73), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1062(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1063(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1064(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1247(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1248(.a(gate390inter0), .b(s_100), .O(gate390inter1));
  and2  gate1249(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1250(.a(s_100), .O(gate390inter3));
  inv1  gate1251(.a(s_101), .O(gate390inter4));
  nand2 gate1252(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1253(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1254(.a(G4), .O(gate390inter7));
  inv1  gate1255(.a(G1045), .O(gate390inter8));
  nand2 gate1256(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1257(.a(s_101), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1258(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1259(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1260(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2409(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2410(.a(gate394inter0), .b(s_266), .O(gate394inter1));
  and2  gate2411(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2412(.a(s_266), .O(gate394inter3));
  inv1  gate2413(.a(s_267), .O(gate394inter4));
  nand2 gate2414(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2415(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2416(.a(G8), .O(gate394inter7));
  inv1  gate2417(.a(G1057), .O(gate394inter8));
  nand2 gate2418(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2419(.a(s_267), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2420(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2421(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2422(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate2927(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2928(.a(gate395inter0), .b(s_340), .O(gate395inter1));
  and2  gate2929(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2930(.a(s_340), .O(gate395inter3));
  inv1  gate2931(.a(s_341), .O(gate395inter4));
  nand2 gate2932(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2933(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2934(.a(G9), .O(gate395inter7));
  inv1  gate2935(.a(G1060), .O(gate395inter8));
  nand2 gate2936(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2937(.a(s_341), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2938(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2939(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2940(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate589(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate590(.a(gate399inter0), .b(s_6), .O(gate399inter1));
  and2  gate591(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate592(.a(s_6), .O(gate399inter3));
  inv1  gate593(.a(s_7), .O(gate399inter4));
  nand2 gate594(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate595(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate596(.a(G13), .O(gate399inter7));
  inv1  gate597(.a(G1072), .O(gate399inter8));
  nand2 gate598(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate599(.a(s_7), .b(gate399inter3), .O(gate399inter10));
  nor2  gate600(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate601(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate602(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate743(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate744(.a(gate402inter0), .b(s_28), .O(gate402inter1));
  and2  gate745(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate746(.a(s_28), .O(gate402inter3));
  inv1  gate747(.a(s_29), .O(gate402inter4));
  nand2 gate748(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate749(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate750(.a(G16), .O(gate402inter7));
  inv1  gate751(.a(G1081), .O(gate402inter8));
  nand2 gate752(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate753(.a(s_29), .b(gate402inter3), .O(gate402inter10));
  nor2  gate754(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate755(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate756(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1821(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1822(.a(gate404inter0), .b(s_182), .O(gate404inter1));
  and2  gate1823(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1824(.a(s_182), .O(gate404inter3));
  inv1  gate1825(.a(s_183), .O(gate404inter4));
  nand2 gate1826(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1827(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1828(.a(G18), .O(gate404inter7));
  inv1  gate1829(.a(G1087), .O(gate404inter8));
  nand2 gate1830(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1831(.a(s_183), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1832(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1833(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1834(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate3053(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate3054(.a(gate405inter0), .b(s_358), .O(gate405inter1));
  and2  gate3055(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate3056(.a(s_358), .O(gate405inter3));
  inv1  gate3057(.a(s_359), .O(gate405inter4));
  nand2 gate3058(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate3059(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate3060(.a(G19), .O(gate405inter7));
  inv1  gate3061(.a(G1090), .O(gate405inter8));
  nand2 gate3062(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate3063(.a(s_359), .b(gate405inter3), .O(gate405inter10));
  nor2  gate3064(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate3065(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate3066(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2073(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2074(.a(gate406inter0), .b(s_218), .O(gate406inter1));
  and2  gate2075(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2076(.a(s_218), .O(gate406inter3));
  inv1  gate2077(.a(s_219), .O(gate406inter4));
  nand2 gate2078(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2079(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2080(.a(G20), .O(gate406inter7));
  inv1  gate2081(.a(G1093), .O(gate406inter8));
  nand2 gate2082(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2083(.a(s_219), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2084(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2085(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2086(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2465(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2466(.a(gate408inter0), .b(s_274), .O(gate408inter1));
  and2  gate2467(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2468(.a(s_274), .O(gate408inter3));
  inv1  gate2469(.a(s_275), .O(gate408inter4));
  nand2 gate2470(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2471(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2472(.a(G22), .O(gate408inter7));
  inv1  gate2473(.a(G1099), .O(gate408inter8));
  nand2 gate2474(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2475(.a(s_275), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2476(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2477(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2478(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1065(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1066(.a(gate409inter0), .b(s_74), .O(gate409inter1));
  and2  gate1067(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1068(.a(s_74), .O(gate409inter3));
  inv1  gate1069(.a(s_75), .O(gate409inter4));
  nand2 gate1070(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1071(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1072(.a(G23), .O(gate409inter7));
  inv1  gate1073(.a(G1102), .O(gate409inter8));
  nand2 gate1074(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1075(.a(s_75), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1076(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1077(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1078(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1149(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1150(.a(gate410inter0), .b(s_86), .O(gate410inter1));
  and2  gate1151(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1152(.a(s_86), .O(gate410inter3));
  inv1  gate1153(.a(s_87), .O(gate410inter4));
  nand2 gate1154(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1155(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1156(.a(G24), .O(gate410inter7));
  inv1  gate1157(.a(G1105), .O(gate410inter8));
  nand2 gate1158(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1159(.a(s_87), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1160(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1161(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1162(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2801(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2802(.a(gate412inter0), .b(s_322), .O(gate412inter1));
  and2  gate2803(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2804(.a(s_322), .O(gate412inter3));
  inv1  gate2805(.a(s_323), .O(gate412inter4));
  nand2 gate2806(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2807(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2808(.a(G26), .O(gate412inter7));
  inv1  gate2809(.a(G1111), .O(gate412inter8));
  nand2 gate2810(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2811(.a(s_323), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2812(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2813(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2814(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1443(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1444(.a(gate413inter0), .b(s_128), .O(gate413inter1));
  and2  gate1445(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1446(.a(s_128), .O(gate413inter3));
  inv1  gate1447(.a(s_129), .O(gate413inter4));
  nand2 gate1448(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1449(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1450(.a(G27), .O(gate413inter7));
  inv1  gate1451(.a(G1114), .O(gate413inter8));
  nand2 gate1452(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1453(.a(s_129), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1454(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1455(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1456(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate911(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate912(.a(gate415inter0), .b(s_52), .O(gate415inter1));
  and2  gate913(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate914(.a(s_52), .O(gate415inter3));
  inv1  gate915(.a(s_53), .O(gate415inter4));
  nand2 gate916(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate917(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate918(.a(G29), .O(gate415inter7));
  inv1  gate919(.a(G1120), .O(gate415inter8));
  nand2 gate920(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate921(.a(s_53), .b(gate415inter3), .O(gate415inter10));
  nor2  gate922(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate923(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate924(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1555(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1556(.a(gate419inter0), .b(s_144), .O(gate419inter1));
  and2  gate1557(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1558(.a(s_144), .O(gate419inter3));
  inv1  gate1559(.a(s_145), .O(gate419inter4));
  nand2 gate1560(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1561(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1562(.a(G1), .O(gate419inter7));
  inv1  gate1563(.a(G1132), .O(gate419inter8));
  nand2 gate1564(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1565(.a(s_145), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1566(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1567(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1568(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1331(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1332(.a(gate420inter0), .b(s_112), .O(gate420inter1));
  and2  gate1333(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1334(.a(s_112), .O(gate420inter3));
  inv1  gate1335(.a(s_113), .O(gate420inter4));
  nand2 gate1336(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1337(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1338(.a(G1036), .O(gate420inter7));
  inv1  gate1339(.a(G1132), .O(gate420inter8));
  nand2 gate1340(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1341(.a(s_113), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1342(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1343(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1344(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2283(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2284(.a(gate428inter0), .b(s_248), .O(gate428inter1));
  and2  gate2285(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2286(.a(s_248), .O(gate428inter3));
  inv1  gate2287(.a(s_249), .O(gate428inter4));
  nand2 gate2288(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2289(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2290(.a(G1048), .O(gate428inter7));
  inv1  gate2291(.a(G1144), .O(gate428inter8));
  nand2 gate2292(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2293(.a(s_249), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2294(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2295(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2296(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1345(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1346(.a(gate429inter0), .b(s_114), .O(gate429inter1));
  and2  gate1347(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1348(.a(s_114), .O(gate429inter3));
  inv1  gate1349(.a(s_115), .O(gate429inter4));
  nand2 gate1350(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1351(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1352(.a(G6), .O(gate429inter7));
  inv1  gate1353(.a(G1147), .O(gate429inter8));
  nand2 gate1354(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1355(.a(s_115), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1356(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1357(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1358(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate3165(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate3166(.a(gate430inter0), .b(s_374), .O(gate430inter1));
  and2  gate3167(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate3168(.a(s_374), .O(gate430inter3));
  inv1  gate3169(.a(s_375), .O(gate430inter4));
  nand2 gate3170(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate3171(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate3172(.a(G1051), .O(gate430inter7));
  inv1  gate3173(.a(G1147), .O(gate430inter8));
  nand2 gate3174(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate3175(.a(s_375), .b(gate430inter3), .O(gate430inter10));
  nor2  gate3176(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate3177(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate3178(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2703(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2704(.a(gate431inter0), .b(s_308), .O(gate431inter1));
  and2  gate2705(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2706(.a(s_308), .O(gate431inter3));
  inv1  gate2707(.a(s_309), .O(gate431inter4));
  nand2 gate2708(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2709(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2710(.a(G7), .O(gate431inter7));
  inv1  gate2711(.a(G1150), .O(gate431inter8));
  nand2 gate2712(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2713(.a(s_309), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2714(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2715(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2716(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2745(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2746(.a(gate432inter0), .b(s_314), .O(gate432inter1));
  and2  gate2747(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2748(.a(s_314), .O(gate432inter3));
  inv1  gate2749(.a(s_315), .O(gate432inter4));
  nand2 gate2750(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2751(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2752(.a(G1054), .O(gate432inter7));
  inv1  gate2753(.a(G1150), .O(gate432inter8));
  nand2 gate2754(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2755(.a(s_315), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2756(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2757(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2758(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate869(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate870(.a(gate433inter0), .b(s_46), .O(gate433inter1));
  and2  gate871(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate872(.a(s_46), .O(gate433inter3));
  inv1  gate873(.a(s_47), .O(gate433inter4));
  nand2 gate874(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate875(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate876(.a(G8), .O(gate433inter7));
  inv1  gate877(.a(G1153), .O(gate433inter8));
  nand2 gate878(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate879(.a(s_47), .b(gate433inter3), .O(gate433inter10));
  nor2  gate880(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate881(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate882(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1135(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1136(.a(gate434inter0), .b(s_84), .O(gate434inter1));
  and2  gate1137(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1138(.a(s_84), .O(gate434inter3));
  inv1  gate1139(.a(s_85), .O(gate434inter4));
  nand2 gate1140(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1141(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1142(.a(G1057), .O(gate434inter7));
  inv1  gate1143(.a(G1153), .O(gate434inter8));
  nand2 gate1144(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1145(.a(s_85), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1146(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1147(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1148(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1541(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1542(.a(gate437inter0), .b(s_142), .O(gate437inter1));
  and2  gate1543(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1544(.a(s_142), .O(gate437inter3));
  inv1  gate1545(.a(s_143), .O(gate437inter4));
  nand2 gate1546(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1547(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1548(.a(G10), .O(gate437inter7));
  inv1  gate1549(.a(G1159), .O(gate437inter8));
  nand2 gate1550(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1551(.a(s_143), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1552(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1553(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1554(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate813(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate814(.a(gate439inter0), .b(s_38), .O(gate439inter1));
  and2  gate815(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate816(.a(s_38), .O(gate439inter3));
  inv1  gate817(.a(s_39), .O(gate439inter4));
  nand2 gate818(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate819(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate820(.a(G11), .O(gate439inter7));
  inv1  gate821(.a(G1162), .O(gate439inter8));
  nand2 gate822(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate823(.a(s_39), .b(gate439inter3), .O(gate439inter10));
  nor2  gate824(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate825(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate826(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate995(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate996(.a(gate440inter0), .b(s_64), .O(gate440inter1));
  and2  gate997(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate998(.a(s_64), .O(gate440inter3));
  inv1  gate999(.a(s_65), .O(gate440inter4));
  nand2 gate1000(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1001(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1002(.a(G1066), .O(gate440inter7));
  inv1  gate1003(.a(G1162), .O(gate440inter8));
  nand2 gate1004(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1005(.a(s_65), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1006(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1007(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1008(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2017(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2018(.a(gate442inter0), .b(s_210), .O(gate442inter1));
  and2  gate2019(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2020(.a(s_210), .O(gate442inter3));
  inv1  gate2021(.a(s_211), .O(gate442inter4));
  nand2 gate2022(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2023(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2024(.a(G1069), .O(gate442inter7));
  inv1  gate2025(.a(G1165), .O(gate442inter8));
  nand2 gate2026(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2027(.a(s_211), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2028(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2029(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2030(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1807(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1808(.a(gate444inter0), .b(s_180), .O(gate444inter1));
  and2  gate1809(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1810(.a(s_180), .O(gate444inter3));
  inv1  gate1811(.a(s_181), .O(gate444inter4));
  nand2 gate1812(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1813(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1814(.a(G1072), .O(gate444inter7));
  inv1  gate1815(.a(G1168), .O(gate444inter8));
  nand2 gate1816(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1817(.a(s_181), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1818(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1819(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1820(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate687(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate688(.a(gate445inter0), .b(s_20), .O(gate445inter1));
  and2  gate689(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate690(.a(s_20), .O(gate445inter3));
  inv1  gate691(.a(s_21), .O(gate445inter4));
  nand2 gate692(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate693(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate694(.a(G14), .O(gate445inter7));
  inv1  gate695(.a(G1171), .O(gate445inter8));
  nand2 gate696(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate697(.a(s_21), .b(gate445inter3), .O(gate445inter10));
  nor2  gate698(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate699(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate700(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate2003(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2004(.a(gate447inter0), .b(s_208), .O(gate447inter1));
  and2  gate2005(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2006(.a(s_208), .O(gate447inter3));
  inv1  gate2007(.a(s_209), .O(gate447inter4));
  nand2 gate2008(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2009(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2010(.a(G15), .O(gate447inter7));
  inv1  gate2011(.a(G1174), .O(gate447inter8));
  nand2 gate2012(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2013(.a(s_209), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2014(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2015(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2016(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate617(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate618(.a(gate448inter0), .b(s_10), .O(gate448inter1));
  and2  gate619(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate620(.a(s_10), .O(gate448inter3));
  inv1  gate621(.a(s_11), .O(gate448inter4));
  nand2 gate622(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate623(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate624(.a(G1078), .O(gate448inter7));
  inv1  gate625(.a(G1174), .O(gate448inter8));
  nand2 gate626(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate627(.a(s_11), .b(gate448inter3), .O(gate448inter10));
  nor2  gate628(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate629(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate630(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1037(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1038(.a(gate449inter0), .b(s_70), .O(gate449inter1));
  and2  gate1039(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1040(.a(s_70), .O(gate449inter3));
  inv1  gate1041(.a(s_71), .O(gate449inter4));
  nand2 gate1042(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1043(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1044(.a(G16), .O(gate449inter7));
  inv1  gate1045(.a(G1177), .O(gate449inter8));
  nand2 gate1046(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1047(.a(s_71), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1048(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1049(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1050(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1261(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1262(.a(gate450inter0), .b(s_102), .O(gate450inter1));
  and2  gate1263(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1264(.a(s_102), .O(gate450inter3));
  inv1  gate1265(.a(s_103), .O(gate450inter4));
  nand2 gate1266(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1267(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1268(.a(G1081), .O(gate450inter7));
  inv1  gate1269(.a(G1177), .O(gate450inter8));
  nand2 gate1270(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1271(.a(s_103), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1272(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1273(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1274(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1373(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1374(.a(gate451inter0), .b(s_118), .O(gate451inter1));
  and2  gate1375(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1376(.a(s_118), .O(gate451inter3));
  inv1  gate1377(.a(s_119), .O(gate451inter4));
  nand2 gate1378(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1379(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1380(.a(G17), .O(gate451inter7));
  inv1  gate1381(.a(G1180), .O(gate451inter8));
  nand2 gate1382(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1383(.a(s_119), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1384(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1385(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1386(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate953(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate954(.a(gate452inter0), .b(s_58), .O(gate452inter1));
  and2  gate955(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate956(.a(s_58), .O(gate452inter3));
  inv1  gate957(.a(s_59), .O(gate452inter4));
  nand2 gate958(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate959(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate960(.a(G1084), .O(gate452inter7));
  inv1  gate961(.a(G1180), .O(gate452inter8));
  nand2 gate962(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate963(.a(s_59), .b(gate452inter3), .O(gate452inter10));
  nor2  gate964(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate965(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate966(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2619(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2620(.a(gate455inter0), .b(s_296), .O(gate455inter1));
  and2  gate2621(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2622(.a(s_296), .O(gate455inter3));
  inv1  gate2623(.a(s_297), .O(gate455inter4));
  nand2 gate2624(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2625(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2626(.a(G19), .O(gate455inter7));
  inv1  gate2627(.a(G1186), .O(gate455inter8));
  nand2 gate2628(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2629(.a(s_297), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2630(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2631(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2632(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate827(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate828(.a(gate458inter0), .b(s_40), .O(gate458inter1));
  and2  gate829(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate830(.a(s_40), .O(gate458inter3));
  inv1  gate831(.a(s_41), .O(gate458inter4));
  nand2 gate832(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate833(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate834(.a(G1093), .O(gate458inter7));
  inv1  gate835(.a(G1189), .O(gate458inter8));
  nand2 gate836(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate837(.a(s_41), .b(gate458inter3), .O(gate458inter10));
  nor2  gate838(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate839(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate840(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1625(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1626(.a(gate459inter0), .b(s_154), .O(gate459inter1));
  and2  gate1627(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1628(.a(s_154), .O(gate459inter3));
  inv1  gate1629(.a(s_155), .O(gate459inter4));
  nand2 gate1630(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1631(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1632(.a(G21), .O(gate459inter7));
  inv1  gate1633(.a(G1192), .O(gate459inter8));
  nand2 gate1634(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1635(.a(s_155), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1636(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1637(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1638(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate561(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate562(.a(gate460inter0), .b(s_2), .O(gate460inter1));
  and2  gate563(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate564(.a(s_2), .O(gate460inter3));
  inv1  gate565(.a(s_3), .O(gate460inter4));
  nand2 gate566(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate567(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate568(.a(G1096), .O(gate460inter7));
  inv1  gate569(.a(G1192), .O(gate460inter8));
  nand2 gate570(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate571(.a(s_3), .b(gate460inter3), .O(gate460inter10));
  nor2  gate572(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate573(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate574(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate967(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate968(.a(gate461inter0), .b(s_60), .O(gate461inter1));
  and2  gate969(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate970(.a(s_60), .O(gate461inter3));
  inv1  gate971(.a(s_61), .O(gate461inter4));
  nand2 gate972(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate973(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate974(.a(G22), .O(gate461inter7));
  inv1  gate975(.a(G1195), .O(gate461inter8));
  nand2 gate976(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate977(.a(s_61), .b(gate461inter3), .O(gate461inter10));
  nor2  gate978(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate979(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate980(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate3011(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate3012(.a(gate466inter0), .b(s_352), .O(gate466inter1));
  and2  gate3013(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate3014(.a(s_352), .O(gate466inter3));
  inv1  gate3015(.a(s_353), .O(gate466inter4));
  nand2 gate3016(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate3017(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate3018(.a(G1105), .O(gate466inter7));
  inv1  gate3019(.a(G1201), .O(gate466inter8));
  nand2 gate3020(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate3021(.a(s_353), .b(gate466inter3), .O(gate466inter10));
  nor2  gate3022(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate3023(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate3024(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1401(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1402(.a(gate468inter0), .b(s_122), .O(gate468inter1));
  and2  gate1403(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1404(.a(s_122), .O(gate468inter3));
  inv1  gate1405(.a(s_123), .O(gate468inter4));
  nand2 gate1406(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1407(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1408(.a(G1108), .O(gate468inter7));
  inv1  gate1409(.a(G1204), .O(gate468inter8));
  nand2 gate1410(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1411(.a(s_123), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1412(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1413(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1414(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate2549(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2550(.a(gate469inter0), .b(s_286), .O(gate469inter1));
  and2  gate2551(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2552(.a(s_286), .O(gate469inter3));
  inv1  gate2553(.a(s_287), .O(gate469inter4));
  nand2 gate2554(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2555(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2556(.a(G26), .O(gate469inter7));
  inv1  gate2557(.a(G1207), .O(gate469inter8));
  nand2 gate2558(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2559(.a(s_287), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2560(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2561(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2562(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate3207(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate3208(.a(gate473inter0), .b(s_380), .O(gate473inter1));
  and2  gate3209(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate3210(.a(s_380), .O(gate473inter3));
  inv1  gate3211(.a(s_381), .O(gate473inter4));
  nand2 gate3212(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate3213(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate3214(.a(G28), .O(gate473inter7));
  inv1  gate3215(.a(G1213), .O(gate473inter8));
  nand2 gate3216(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate3217(.a(s_381), .b(gate473inter3), .O(gate473inter10));
  nor2  gate3218(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate3219(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate3220(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2605(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2606(.a(gate478inter0), .b(s_294), .O(gate478inter1));
  and2  gate2607(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2608(.a(s_294), .O(gate478inter3));
  inv1  gate2609(.a(s_295), .O(gate478inter4));
  nand2 gate2610(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2611(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2612(.a(G1123), .O(gate478inter7));
  inv1  gate2613(.a(G1219), .O(gate478inter8));
  nand2 gate2614(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2615(.a(s_295), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2616(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2617(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2618(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2871(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2872(.a(gate479inter0), .b(s_332), .O(gate479inter1));
  and2  gate2873(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2874(.a(s_332), .O(gate479inter3));
  inv1  gate2875(.a(s_333), .O(gate479inter4));
  nand2 gate2876(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2877(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2878(.a(G31), .O(gate479inter7));
  inv1  gate2879(.a(G1222), .O(gate479inter8));
  nand2 gate2880(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2881(.a(s_333), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2882(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2883(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2884(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1723(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1724(.a(gate480inter0), .b(s_168), .O(gate480inter1));
  and2  gate1725(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1726(.a(s_168), .O(gate480inter3));
  inv1  gate1727(.a(s_169), .O(gate480inter4));
  nand2 gate1728(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1729(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1730(.a(G1126), .O(gate480inter7));
  inv1  gate1731(.a(G1222), .O(gate480inter8));
  nand2 gate1732(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1733(.a(s_169), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1734(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1735(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1736(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate3025(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate3026(.a(gate486inter0), .b(s_354), .O(gate486inter1));
  and2  gate3027(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate3028(.a(s_354), .O(gate486inter3));
  inv1  gate3029(.a(s_355), .O(gate486inter4));
  nand2 gate3030(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate3031(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate3032(.a(G1234), .O(gate486inter7));
  inv1  gate3033(.a(G1235), .O(gate486inter8));
  nand2 gate3034(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate3035(.a(s_355), .b(gate486inter3), .O(gate486inter10));
  nor2  gate3036(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate3037(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate3038(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2325(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2326(.a(gate489inter0), .b(s_254), .O(gate489inter1));
  and2  gate2327(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2328(.a(s_254), .O(gate489inter3));
  inv1  gate2329(.a(s_255), .O(gate489inter4));
  nand2 gate2330(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2331(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2332(.a(G1240), .O(gate489inter7));
  inv1  gate2333(.a(G1241), .O(gate489inter8));
  nand2 gate2334(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2335(.a(s_255), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2336(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2337(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2338(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1751(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1752(.a(gate494inter0), .b(s_172), .O(gate494inter1));
  and2  gate1753(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1754(.a(s_172), .O(gate494inter3));
  inv1  gate1755(.a(s_173), .O(gate494inter4));
  nand2 gate1756(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1757(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1758(.a(G1250), .O(gate494inter7));
  inv1  gate1759(.a(G1251), .O(gate494inter8));
  nand2 gate1760(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1761(.a(s_173), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1762(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1763(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1764(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2101(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2102(.a(gate495inter0), .b(s_222), .O(gate495inter1));
  and2  gate2103(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2104(.a(s_222), .O(gate495inter3));
  inv1  gate2105(.a(s_223), .O(gate495inter4));
  nand2 gate2106(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2107(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2108(.a(G1252), .O(gate495inter7));
  inv1  gate2109(.a(G1253), .O(gate495inter8));
  nand2 gate2110(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2111(.a(s_223), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2112(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2113(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2114(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate2997(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2998(.a(gate496inter0), .b(s_350), .O(gate496inter1));
  and2  gate2999(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate3000(.a(s_350), .O(gate496inter3));
  inv1  gate3001(.a(s_351), .O(gate496inter4));
  nand2 gate3002(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate3003(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate3004(.a(G1254), .O(gate496inter7));
  inv1  gate3005(.a(G1255), .O(gate496inter8));
  nand2 gate3006(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate3007(.a(s_351), .b(gate496inter3), .O(gate496inter10));
  nor2  gate3008(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate3009(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate3010(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate2843(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2844(.a(gate498inter0), .b(s_328), .O(gate498inter1));
  and2  gate2845(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2846(.a(s_328), .O(gate498inter3));
  inv1  gate2847(.a(s_329), .O(gate498inter4));
  nand2 gate2848(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2849(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2850(.a(G1258), .O(gate498inter7));
  inv1  gate2851(.a(G1259), .O(gate498inter8));
  nand2 gate2852(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2853(.a(s_329), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2854(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2855(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2856(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate2941(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2942(.a(gate499inter0), .b(s_342), .O(gate499inter1));
  and2  gate2943(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2944(.a(s_342), .O(gate499inter3));
  inv1  gate2945(.a(s_343), .O(gate499inter4));
  nand2 gate2946(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2947(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2948(.a(G1260), .O(gate499inter7));
  inv1  gate2949(.a(G1261), .O(gate499inter8));
  nand2 gate2950(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2951(.a(s_343), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2952(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2953(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2954(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2171(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2172(.a(gate500inter0), .b(s_232), .O(gate500inter1));
  and2  gate2173(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2174(.a(s_232), .O(gate500inter3));
  inv1  gate2175(.a(s_233), .O(gate500inter4));
  nand2 gate2176(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2177(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2178(.a(G1262), .O(gate500inter7));
  inv1  gate2179(.a(G1263), .O(gate500inter8));
  nand2 gate2180(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2181(.a(s_233), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2182(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2183(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2184(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2129(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2130(.a(gate501inter0), .b(s_226), .O(gate501inter1));
  and2  gate2131(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2132(.a(s_226), .O(gate501inter3));
  inv1  gate2133(.a(s_227), .O(gate501inter4));
  nand2 gate2134(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2135(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2136(.a(G1264), .O(gate501inter7));
  inv1  gate2137(.a(G1265), .O(gate501inter8));
  nand2 gate2138(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2139(.a(s_227), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2140(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2141(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2142(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1485(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1486(.a(gate503inter0), .b(s_134), .O(gate503inter1));
  and2  gate1487(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1488(.a(s_134), .O(gate503inter3));
  inv1  gate1489(.a(s_135), .O(gate503inter4));
  nand2 gate1490(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1491(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1492(.a(G1268), .O(gate503inter7));
  inv1  gate1493(.a(G1269), .O(gate503inter8));
  nand2 gate1494(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1495(.a(s_135), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1496(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1497(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1498(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate883(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate884(.a(gate504inter0), .b(s_48), .O(gate504inter1));
  and2  gate885(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate886(.a(s_48), .O(gate504inter3));
  inv1  gate887(.a(s_49), .O(gate504inter4));
  nand2 gate888(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate889(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate890(.a(G1270), .O(gate504inter7));
  inv1  gate891(.a(G1271), .O(gate504inter8));
  nand2 gate892(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate893(.a(s_49), .b(gate504inter3), .O(gate504inter10));
  nor2  gate894(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate895(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate896(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate659(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate660(.a(gate512inter0), .b(s_16), .O(gate512inter1));
  and2  gate661(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate662(.a(s_16), .O(gate512inter3));
  inv1  gate663(.a(s_17), .O(gate512inter4));
  nand2 gate664(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate665(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate666(.a(G1286), .O(gate512inter7));
  inv1  gate667(.a(G1287), .O(gate512inter8));
  nand2 gate668(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate669(.a(s_17), .b(gate512inter3), .O(gate512inter10));
  nor2  gate670(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate671(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate672(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1023(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1024(.a(gate513inter0), .b(s_68), .O(gate513inter1));
  and2  gate1025(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1026(.a(s_68), .O(gate513inter3));
  inv1  gate1027(.a(s_69), .O(gate513inter4));
  nand2 gate1028(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1029(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1030(.a(G1288), .O(gate513inter7));
  inv1  gate1031(.a(G1289), .O(gate513inter8));
  nand2 gate1032(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1033(.a(s_69), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1034(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1035(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1036(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1933(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1934(.a(gate514inter0), .b(s_198), .O(gate514inter1));
  and2  gate1935(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1936(.a(s_198), .O(gate514inter3));
  inv1  gate1937(.a(s_199), .O(gate514inter4));
  nand2 gate1938(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1939(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1940(.a(G1290), .O(gate514inter7));
  inv1  gate1941(.a(G1291), .O(gate514inter8));
  nand2 gate1942(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1943(.a(s_199), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1944(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1945(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1946(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule