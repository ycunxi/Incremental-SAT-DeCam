module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1611(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1612(.a(gate11inter0), .b(s_152), .O(gate11inter1));
  and2  gate1613(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1614(.a(s_152), .O(gate11inter3));
  inv1  gate1615(.a(s_153), .O(gate11inter4));
  nand2 gate1616(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1617(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1618(.a(G5), .O(gate11inter7));
  inv1  gate1619(.a(G6), .O(gate11inter8));
  nand2 gate1620(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1621(.a(s_153), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1622(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1623(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1624(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate743(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate744(.a(gate17inter0), .b(s_28), .O(gate17inter1));
  and2  gate745(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate746(.a(s_28), .O(gate17inter3));
  inv1  gate747(.a(s_29), .O(gate17inter4));
  nand2 gate748(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate749(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate750(.a(G17), .O(gate17inter7));
  inv1  gate751(.a(G18), .O(gate17inter8));
  nand2 gate752(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate753(.a(s_29), .b(gate17inter3), .O(gate17inter10));
  nor2  gate754(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate755(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate756(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate925(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate926(.a(gate18inter0), .b(s_54), .O(gate18inter1));
  and2  gate927(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate928(.a(s_54), .O(gate18inter3));
  inv1  gate929(.a(s_55), .O(gate18inter4));
  nand2 gate930(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate931(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate932(.a(G19), .O(gate18inter7));
  inv1  gate933(.a(G20), .O(gate18inter8));
  nand2 gate934(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate935(.a(s_55), .b(gate18inter3), .O(gate18inter10));
  nor2  gate936(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate937(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate938(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1709(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1710(.a(gate22inter0), .b(s_166), .O(gate22inter1));
  and2  gate1711(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1712(.a(s_166), .O(gate22inter3));
  inv1  gate1713(.a(s_167), .O(gate22inter4));
  nand2 gate1714(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1715(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1716(.a(G27), .O(gate22inter7));
  inv1  gate1717(.a(G28), .O(gate22inter8));
  nand2 gate1718(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1719(.a(s_167), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1720(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1721(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1722(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate589(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate590(.a(gate24inter0), .b(s_6), .O(gate24inter1));
  and2  gate591(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate592(.a(s_6), .O(gate24inter3));
  inv1  gate593(.a(s_7), .O(gate24inter4));
  nand2 gate594(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate595(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate596(.a(G31), .O(gate24inter7));
  inv1  gate597(.a(G32), .O(gate24inter8));
  nand2 gate598(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate599(.a(s_7), .b(gate24inter3), .O(gate24inter10));
  nor2  gate600(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate601(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate602(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1975(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1976(.a(gate25inter0), .b(s_204), .O(gate25inter1));
  and2  gate1977(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1978(.a(s_204), .O(gate25inter3));
  inv1  gate1979(.a(s_205), .O(gate25inter4));
  nand2 gate1980(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1981(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1982(.a(G1), .O(gate25inter7));
  inv1  gate1983(.a(G5), .O(gate25inter8));
  nand2 gate1984(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1985(.a(s_205), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1986(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1987(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1988(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1765(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1766(.a(gate31inter0), .b(s_174), .O(gate31inter1));
  and2  gate1767(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1768(.a(s_174), .O(gate31inter3));
  inv1  gate1769(.a(s_175), .O(gate31inter4));
  nand2 gate1770(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1771(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1772(.a(G4), .O(gate31inter7));
  inv1  gate1773(.a(G8), .O(gate31inter8));
  nand2 gate1774(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1775(.a(s_175), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1776(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1777(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1778(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1415(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1416(.a(gate32inter0), .b(s_124), .O(gate32inter1));
  and2  gate1417(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1418(.a(s_124), .O(gate32inter3));
  inv1  gate1419(.a(s_125), .O(gate32inter4));
  nand2 gate1420(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1421(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1422(.a(G12), .O(gate32inter7));
  inv1  gate1423(.a(G16), .O(gate32inter8));
  nand2 gate1424(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1425(.a(s_125), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1426(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1427(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1428(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate827(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate828(.a(gate33inter0), .b(s_40), .O(gate33inter1));
  and2  gate829(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate830(.a(s_40), .O(gate33inter3));
  inv1  gate831(.a(s_41), .O(gate33inter4));
  nand2 gate832(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate833(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate834(.a(G17), .O(gate33inter7));
  inv1  gate835(.a(G21), .O(gate33inter8));
  nand2 gate836(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate837(.a(s_41), .b(gate33inter3), .O(gate33inter10));
  nor2  gate838(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate839(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate840(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1443(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1444(.a(gate36inter0), .b(s_128), .O(gate36inter1));
  and2  gate1445(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1446(.a(s_128), .O(gate36inter3));
  inv1  gate1447(.a(s_129), .O(gate36inter4));
  nand2 gate1448(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1449(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1450(.a(G26), .O(gate36inter7));
  inv1  gate1451(.a(G30), .O(gate36inter8));
  nand2 gate1452(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1453(.a(s_129), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1454(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1455(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1456(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate757(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate758(.a(gate41inter0), .b(s_30), .O(gate41inter1));
  and2  gate759(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate760(.a(s_30), .O(gate41inter3));
  inv1  gate761(.a(s_31), .O(gate41inter4));
  nand2 gate762(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate763(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate764(.a(G1), .O(gate41inter7));
  inv1  gate765(.a(G266), .O(gate41inter8));
  nand2 gate766(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate767(.a(s_31), .b(gate41inter3), .O(gate41inter10));
  nor2  gate768(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate769(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate770(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate799(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate800(.a(gate42inter0), .b(s_36), .O(gate42inter1));
  and2  gate801(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate802(.a(s_36), .O(gate42inter3));
  inv1  gate803(.a(s_37), .O(gate42inter4));
  nand2 gate804(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate805(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate806(.a(G2), .O(gate42inter7));
  inv1  gate807(.a(G266), .O(gate42inter8));
  nand2 gate808(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate809(.a(s_37), .b(gate42inter3), .O(gate42inter10));
  nor2  gate810(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate811(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate812(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1219(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1220(.a(gate48inter0), .b(s_96), .O(gate48inter1));
  and2  gate1221(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1222(.a(s_96), .O(gate48inter3));
  inv1  gate1223(.a(s_97), .O(gate48inter4));
  nand2 gate1224(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1225(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1226(.a(G8), .O(gate48inter7));
  inv1  gate1227(.a(G275), .O(gate48inter8));
  nand2 gate1228(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1229(.a(s_97), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1230(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1231(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1232(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate995(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate996(.a(gate54inter0), .b(s_64), .O(gate54inter1));
  and2  gate997(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate998(.a(s_64), .O(gate54inter3));
  inv1  gate999(.a(s_65), .O(gate54inter4));
  nand2 gate1000(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1001(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1002(.a(G14), .O(gate54inter7));
  inv1  gate1003(.a(G284), .O(gate54inter8));
  nand2 gate1004(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1005(.a(s_65), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1006(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1007(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1008(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1289(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1290(.a(gate58inter0), .b(s_106), .O(gate58inter1));
  and2  gate1291(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1292(.a(s_106), .O(gate58inter3));
  inv1  gate1293(.a(s_107), .O(gate58inter4));
  nand2 gate1294(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1295(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1296(.a(G18), .O(gate58inter7));
  inv1  gate1297(.a(G290), .O(gate58inter8));
  nand2 gate1298(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1299(.a(s_107), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1300(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1301(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1302(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1331(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1332(.a(gate59inter0), .b(s_112), .O(gate59inter1));
  and2  gate1333(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1334(.a(s_112), .O(gate59inter3));
  inv1  gate1335(.a(s_113), .O(gate59inter4));
  nand2 gate1336(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1337(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1338(.a(G19), .O(gate59inter7));
  inv1  gate1339(.a(G293), .O(gate59inter8));
  nand2 gate1340(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1341(.a(s_113), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1342(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1343(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1344(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate701(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate702(.a(gate60inter0), .b(s_22), .O(gate60inter1));
  and2  gate703(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate704(.a(s_22), .O(gate60inter3));
  inv1  gate705(.a(s_23), .O(gate60inter4));
  nand2 gate706(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate707(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate708(.a(G20), .O(gate60inter7));
  inv1  gate709(.a(G293), .O(gate60inter8));
  nand2 gate710(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate711(.a(s_23), .b(gate60inter3), .O(gate60inter10));
  nor2  gate712(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate713(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate714(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate841(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate842(.a(gate62inter0), .b(s_42), .O(gate62inter1));
  and2  gate843(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate844(.a(s_42), .O(gate62inter3));
  inv1  gate845(.a(s_43), .O(gate62inter4));
  nand2 gate846(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate847(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate848(.a(G22), .O(gate62inter7));
  inv1  gate849(.a(G296), .O(gate62inter8));
  nand2 gate850(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate851(.a(s_43), .b(gate62inter3), .O(gate62inter10));
  nor2  gate852(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate853(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate854(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1527(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1528(.a(gate63inter0), .b(s_140), .O(gate63inter1));
  and2  gate1529(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1530(.a(s_140), .O(gate63inter3));
  inv1  gate1531(.a(s_141), .O(gate63inter4));
  nand2 gate1532(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1533(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1534(.a(G23), .O(gate63inter7));
  inv1  gate1535(.a(G299), .O(gate63inter8));
  nand2 gate1536(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1537(.a(s_141), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1538(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1539(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1540(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate939(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate940(.a(gate66inter0), .b(s_56), .O(gate66inter1));
  and2  gate941(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate942(.a(s_56), .O(gate66inter3));
  inv1  gate943(.a(s_57), .O(gate66inter4));
  nand2 gate944(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate945(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate946(.a(G26), .O(gate66inter7));
  inv1  gate947(.a(G302), .O(gate66inter8));
  nand2 gate948(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate949(.a(s_57), .b(gate66inter3), .O(gate66inter10));
  nor2  gate950(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate951(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate952(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2087(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2088(.a(gate77inter0), .b(s_220), .O(gate77inter1));
  and2  gate2089(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2090(.a(s_220), .O(gate77inter3));
  inv1  gate2091(.a(s_221), .O(gate77inter4));
  nand2 gate2092(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2093(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2094(.a(G2), .O(gate77inter7));
  inv1  gate2095(.a(G320), .O(gate77inter8));
  nand2 gate2096(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2097(.a(s_221), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2098(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2099(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2100(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate715(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate716(.a(gate81inter0), .b(s_24), .O(gate81inter1));
  and2  gate717(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate718(.a(s_24), .O(gate81inter3));
  inv1  gate719(.a(s_25), .O(gate81inter4));
  nand2 gate720(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate721(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate722(.a(G3), .O(gate81inter7));
  inv1  gate723(.a(G326), .O(gate81inter8));
  nand2 gate724(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate725(.a(s_25), .b(gate81inter3), .O(gate81inter10));
  nor2  gate726(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate727(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate728(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate813(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate814(.a(gate82inter0), .b(s_38), .O(gate82inter1));
  and2  gate815(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate816(.a(s_38), .O(gate82inter3));
  inv1  gate817(.a(s_39), .O(gate82inter4));
  nand2 gate818(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate819(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate820(.a(G7), .O(gate82inter7));
  inv1  gate821(.a(G326), .O(gate82inter8));
  nand2 gate822(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate823(.a(s_39), .b(gate82inter3), .O(gate82inter10));
  nor2  gate824(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate825(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate826(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate967(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate968(.a(gate87inter0), .b(s_60), .O(gate87inter1));
  and2  gate969(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate970(.a(s_60), .O(gate87inter3));
  inv1  gate971(.a(s_61), .O(gate87inter4));
  nand2 gate972(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate973(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate974(.a(G12), .O(gate87inter7));
  inv1  gate975(.a(G335), .O(gate87inter8));
  nand2 gate976(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate977(.a(s_61), .b(gate87inter3), .O(gate87inter10));
  nor2  gate978(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate979(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate980(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1793(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1794(.a(gate88inter0), .b(s_178), .O(gate88inter1));
  and2  gate1795(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1796(.a(s_178), .O(gate88inter3));
  inv1  gate1797(.a(s_179), .O(gate88inter4));
  nand2 gate1798(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1799(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1800(.a(G16), .O(gate88inter7));
  inv1  gate1801(.a(G335), .O(gate88inter8));
  nand2 gate1802(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1803(.a(s_179), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1804(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1805(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1806(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1093(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1094(.a(gate93inter0), .b(s_78), .O(gate93inter1));
  and2  gate1095(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1096(.a(s_78), .O(gate93inter3));
  inv1  gate1097(.a(s_79), .O(gate93inter4));
  nand2 gate1098(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1099(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1100(.a(G18), .O(gate93inter7));
  inv1  gate1101(.a(G344), .O(gate93inter8));
  nand2 gate1102(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1103(.a(s_79), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1104(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1105(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1106(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1457(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1458(.a(gate107inter0), .b(s_130), .O(gate107inter1));
  and2  gate1459(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1460(.a(s_130), .O(gate107inter3));
  inv1  gate1461(.a(s_131), .O(gate107inter4));
  nand2 gate1462(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1463(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1464(.a(G366), .O(gate107inter7));
  inv1  gate1465(.a(G367), .O(gate107inter8));
  nand2 gate1466(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1467(.a(s_131), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1468(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1469(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1470(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1863(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1864(.a(gate108inter0), .b(s_188), .O(gate108inter1));
  and2  gate1865(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1866(.a(s_188), .O(gate108inter3));
  inv1  gate1867(.a(s_189), .O(gate108inter4));
  nand2 gate1868(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1869(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1870(.a(G368), .O(gate108inter7));
  inv1  gate1871(.a(G369), .O(gate108inter8));
  nand2 gate1872(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1873(.a(s_189), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1874(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1875(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1876(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1625(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1626(.a(gate110inter0), .b(s_154), .O(gate110inter1));
  and2  gate1627(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1628(.a(s_154), .O(gate110inter3));
  inv1  gate1629(.a(s_155), .O(gate110inter4));
  nand2 gate1630(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1631(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1632(.a(G372), .O(gate110inter7));
  inv1  gate1633(.a(G373), .O(gate110inter8));
  nand2 gate1634(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1635(.a(s_155), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1636(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1637(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1638(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2073(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2074(.a(gate112inter0), .b(s_218), .O(gate112inter1));
  and2  gate2075(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2076(.a(s_218), .O(gate112inter3));
  inv1  gate2077(.a(s_219), .O(gate112inter4));
  nand2 gate2078(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2079(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2080(.a(G376), .O(gate112inter7));
  inv1  gate2081(.a(G377), .O(gate112inter8));
  nand2 gate2082(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2083(.a(s_219), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2084(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2085(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2086(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate883(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate884(.a(gate113inter0), .b(s_48), .O(gate113inter1));
  and2  gate885(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate886(.a(s_48), .O(gate113inter3));
  inv1  gate887(.a(s_49), .O(gate113inter4));
  nand2 gate888(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate889(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate890(.a(G378), .O(gate113inter7));
  inv1  gate891(.a(G379), .O(gate113inter8));
  nand2 gate892(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate893(.a(s_49), .b(gate113inter3), .O(gate113inter10));
  nor2  gate894(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate895(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate896(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1065(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1066(.a(gate115inter0), .b(s_74), .O(gate115inter1));
  and2  gate1067(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1068(.a(s_74), .O(gate115inter3));
  inv1  gate1069(.a(s_75), .O(gate115inter4));
  nand2 gate1070(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1071(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1072(.a(G382), .O(gate115inter7));
  inv1  gate1073(.a(G383), .O(gate115inter8));
  nand2 gate1074(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1075(.a(s_75), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1076(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1077(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1078(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1359(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1360(.a(gate131inter0), .b(s_116), .O(gate131inter1));
  and2  gate1361(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1362(.a(s_116), .O(gate131inter3));
  inv1  gate1363(.a(s_117), .O(gate131inter4));
  nand2 gate1364(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1365(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1366(.a(G414), .O(gate131inter7));
  inv1  gate1367(.a(G415), .O(gate131inter8));
  nand2 gate1368(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1369(.a(s_117), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1370(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1371(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1372(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1947(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1948(.a(gate134inter0), .b(s_200), .O(gate134inter1));
  and2  gate1949(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1950(.a(s_200), .O(gate134inter3));
  inv1  gate1951(.a(s_201), .O(gate134inter4));
  nand2 gate1952(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1953(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1954(.a(G420), .O(gate134inter7));
  inv1  gate1955(.a(G421), .O(gate134inter8));
  nand2 gate1956(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1957(.a(s_201), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1958(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1959(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1960(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1919(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1920(.a(gate136inter0), .b(s_196), .O(gate136inter1));
  and2  gate1921(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1922(.a(s_196), .O(gate136inter3));
  inv1  gate1923(.a(s_197), .O(gate136inter4));
  nand2 gate1924(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1925(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1926(.a(G424), .O(gate136inter7));
  inv1  gate1927(.a(G425), .O(gate136inter8));
  nand2 gate1928(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1929(.a(s_197), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1930(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1931(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1932(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1429(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1430(.a(gate142inter0), .b(s_126), .O(gate142inter1));
  and2  gate1431(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1432(.a(s_126), .O(gate142inter3));
  inv1  gate1433(.a(s_127), .O(gate142inter4));
  nand2 gate1434(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1435(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1436(.a(G456), .O(gate142inter7));
  inv1  gate1437(.a(G459), .O(gate142inter8));
  nand2 gate1438(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1439(.a(s_127), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1440(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1441(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1442(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate897(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate898(.a(gate143inter0), .b(s_50), .O(gate143inter1));
  and2  gate899(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate900(.a(s_50), .O(gate143inter3));
  inv1  gate901(.a(s_51), .O(gate143inter4));
  nand2 gate902(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate903(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate904(.a(G462), .O(gate143inter7));
  inv1  gate905(.a(G465), .O(gate143inter8));
  nand2 gate906(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate907(.a(s_51), .b(gate143inter3), .O(gate143inter10));
  nor2  gate908(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate909(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate910(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate673(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate674(.a(gate150inter0), .b(s_18), .O(gate150inter1));
  and2  gate675(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate676(.a(s_18), .O(gate150inter3));
  inv1  gate677(.a(s_19), .O(gate150inter4));
  nand2 gate678(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate679(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate680(.a(G504), .O(gate150inter7));
  inv1  gate681(.a(G507), .O(gate150inter8));
  nand2 gate682(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate683(.a(s_19), .b(gate150inter3), .O(gate150inter10));
  nor2  gate684(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate685(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate686(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1471(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1472(.a(gate151inter0), .b(s_132), .O(gate151inter1));
  and2  gate1473(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1474(.a(s_132), .O(gate151inter3));
  inv1  gate1475(.a(s_133), .O(gate151inter4));
  nand2 gate1476(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1477(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1478(.a(G510), .O(gate151inter7));
  inv1  gate1479(.a(G513), .O(gate151inter8));
  nand2 gate1480(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1481(.a(s_133), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1482(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1483(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1484(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1639(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1640(.a(gate154inter0), .b(s_156), .O(gate154inter1));
  and2  gate1641(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1642(.a(s_156), .O(gate154inter3));
  inv1  gate1643(.a(s_157), .O(gate154inter4));
  nand2 gate1644(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1645(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1646(.a(G429), .O(gate154inter7));
  inv1  gate1647(.a(G522), .O(gate154inter8));
  nand2 gate1648(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1649(.a(s_157), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1650(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1651(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1652(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1555(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1556(.a(gate158inter0), .b(s_144), .O(gate158inter1));
  and2  gate1557(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1558(.a(s_144), .O(gate158inter3));
  inv1  gate1559(.a(s_145), .O(gate158inter4));
  nand2 gate1560(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1561(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1562(.a(G441), .O(gate158inter7));
  inv1  gate1563(.a(G528), .O(gate158inter8));
  nand2 gate1564(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1565(.a(s_145), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1566(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1567(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1568(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2045(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2046(.a(gate162inter0), .b(s_214), .O(gate162inter1));
  and2  gate2047(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2048(.a(s_214), .O(gate162inter3));
  inv1  gate2049(.a(s_215), .O(gate162inter4));
  nand2 gate2050(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2051(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2052(.a(G453), .O(gate162inter7));
  inv1  gate2053(.a(G534), .O(gate162inter8));
  nand2 gate2054(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2055(.a(s_215), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2056(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2057(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2058(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1891(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1892(.a(gate170inter0), .b(s_192), .O(gate170inter1));
  and2  gate1893(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1894(.a(s_192), .O(gate170inter3));
  inv1  gate1895(.a(s_193), .O(gate170inter4));
  nand2 gate1896(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1897(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1898(.a(G477), .O(gate170inter7));
  inv1  gate1899(.a(G546), .O(gate170inter8));
  nand2 gate1900(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1901(.a(s_193), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1902(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1903(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1904(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1807(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1808(.a(gate172inter0), .b(s_180), .O(gate172inter1));
  and2  gate1809(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1810(.a(s_180), .O(gate172inter3));
  inv1  gate1811(.a(s_181), .O(gate172inter4));
  nand2 gate1812(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1813(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1814(.a(G483), .O(gate172inter7));
  inv1  gate1815(.a(G549), .O(gate172inter8));
  nand2 gate1816(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1817(.a(s_181), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1818(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1819(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1820(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1681(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1682(.a(gate173inter0), .b(s_162), .O(gate173inter1));
  and2  gate1683(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1684(.a(s_162), .O(gate173inter3));
  inv1  gate1685(.a(s_163), .O(gate173inter4));
  nand2 gate1686(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1687(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1688(.a(G486), .O(gate173inter7));
  inv1  gate1689(.a(G552), .O(gate173inter8));
  nand2 gate1690(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1691(.a(s_163), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1692(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1693(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1694(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1051(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1052(.a(gate175inter0), .b(s_72), .O(gate175inter1));
  and2  gate1053(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1054(.a(s_72), .O(gate175inter3));
  inv1  gate1055(.a(s_73), .O(gate175inter4));
  nand2 gate1056(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1057(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1058(.a(G492), .O(gate175inter7));
  inv1  gate1059(.a(G555), .O(gate175inter8));
  nand2 gate1060(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1061(.a(s_73), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1062(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1063(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1064(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1849(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1850(.a(gate176inter0), .b(s_186), .O(gate176inter1));
  and2  gate1851(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1852(.a(s_186), .O(gate176inter3));
  inv1  gate1853(.a(s_187), .O(gate176inter4));
  nand2 gate1854(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1855(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1856(.a(G495), .O(gate176inter7));
  inv1  gate1857(.a(G555), .O(gate176inter8));
  nand2 gate1858(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1859(.a(s_187), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1860(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1861(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1862(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate687(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate688(.a(gate179inter0), .b(s_20), .O(gate179inter1));
  and2  gate689(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate690(.a(s_20), .O(gate179inter3));
  inv1  gate691(.a(s_21), .O(gate179inter4));
  nand2 gate692(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate693(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate694(.a(G504), .O(gate179inter7));
  inv1  gate695(.a(G561), .O(gate179inter8));
  nand2 gate696(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate697(.a(s_21), .b(gate179inter3), .O(gate179inter10));
  nor2  gate698(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate699(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate700(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate869(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate870(.a(gate183inter0), .b(s_46), .O(gate183inter1));
  and2  gate871(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate872(.a(s_46), .O(gate183inter3));
  inv1  gate873(.a(s_47), .O(gate183inter4));
  nand2 gate874(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate875(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate876(.a(G516), .O(gate183inter7));
  inv1  gate877(.a(G567), .O(gate183inter8));
  nand2 gate878(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate879(.a(s_47), .b(gate183inter3), .O(gate183inter10));
  nor2  gate880(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate881(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate882(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1121(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1122(.a(gate191inter0), .b(s_82), .O(gate191inter1));
  and2  gate1123(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1124(.a(s_82), .O(gate191inter3));
  inv1  gate1125(.a(s_83), .O(gate191inter4));
  nand2 gate1126(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1127(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1128(.a(G582), .O(gate191inter7));
  inv1  gate1129(.a(G583), .O(gate191inter8));
  nand2 gate1130(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1131(.a(s_83), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1132(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1133(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1134(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2101(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2102(.a(gate198inter0), .b(s_222), .O(gate198inter1));
  and2  gate2103(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2104(.a(s_222), .O(gate198inter3));
  inv1  gate2105(.a(s_223), .O(gate198inter4));
  nand2 gate2106(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2107(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2108(.a(G596), .O(gate198inter7));
  inv1  gate2109(.a(G597), .O(gate198inter8));
  nand2 gate2110(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2111(.a(s_223), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2112(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2113(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2114(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1723(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1724(.a(gate200inter0), .b(s_168), .O(gate200inter1));
  and2  gate1725(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1726(.a(s_168), .O(gate200inter3));
  inv1  gate1727(.a(s_169), .O(gate200inter4));
  nand2 gate1728(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1729(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1730(.a(G600), .O(gate200inter7));
  inv1  gate1731(.a(G601), .O(gate200inter8));
  nand2 gate1732(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1733(.a(s_169), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1734(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1735(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1736(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate911(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate912(.a(gate201inter0), .b(s_52), .O(gate201inter1));
  and2  gate913(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate914(.a(s_52), .O(gate201inter3));
  inv1  gate915(.a(s_53), .O(gate201inter4));
  nand2 gate916(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate917(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate918(.a(G602), .O(gate201inter7));
  inv1  gate919(.a(G607), .O(gate201inter8));
  nand2 gate920(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate921(.a(s_53), .b(gate201inter3), .O(gate201inter10));
  nor2  gate922(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate923(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate924(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2129(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2130(.a(gate203inter0), .b(s_226), .O(gate203inter1));
  and2  gate2131(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2132(.a(s_226), .O(gate203inter3));
  inv1  gate2133(.a(s_227), .O(gate203inter4));
  nand2 gate2134(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2135(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2136(.a(G602), .O(gate203inter7));
  inv1  gate2137(.a(G612), .O(gate203inter8));
  nand2 gate2138(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2139(.a(s_227), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2140(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2141(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2142(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1261(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1262(.a(gate206inter0), .b(s_102), .O(gate206inter1));
  and2  gate1263(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1264(.a(s_102), .O(gate206inter3));
  inv1  gate1265(.a(s_103), .O(gate206inter4));
  nand2 gate1266(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1267(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1268(.a(G632), .O(gate206inter7));
  inv1  gate1269(.a(G637), .O(gate206inter8));
  nand2 gate1270(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1271(.a(s_103), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1272(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1273(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1274(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1387(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1388(.a(gate210inter0), .b(s_120), .O(gate210inter1));
  and2  gate1389(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1390(.a(s_120), .O(gate210inter3));
  inv1  gate1391(.a(s_121), .O(gate210inter4));
  nand2 gate1392(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1393(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1394(.a(G607), .O(gate210inter7));
  inv1  gate1395(.a(G666), .O(gate210inter8));
  nand2 gate1396(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1397(.a(s_121), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1398(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1399(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1400(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1835(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1836(.a(gate211inter0), .b(s_184), .O(gate211inter1));
  and2  gate1837(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1838(.a(s_184), .O(gate211inter3));
  inv1  gate1839(.a(s_185), .O(gate211inter4));
  nand2 gate1840(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1841(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1842(.a(G612), .O(gate211inter7));
  inv1  gate1843(.a(G669), .O(gate211inter8));
  nand2 gate1844(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1845(.a(s_185), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1846(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1847(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1848(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1401(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1402(.a(gate212inter0), .b(s_122), .O(gate212inter1));
  and2  gate1403(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1404(.a(s_122), .O(gate212inter3));
  inv1  gate1405(.a(s_123), .O(gate212inter4));
  nand2 gate1406(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1407(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1408(.a(G617), .O(gate212inter7));
  inv1  gate1409(.a(G669), .O(gate212inter8));
  nand2 gate1410(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1411(.a(s_123), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1412(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1413(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1414(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate645(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate646(.a(gate218inter0), .b(s_14), .O(gate218inter1));
  and2  gate647(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate648(.a(s_14), .O(gate218inter3));
  inv1  gate649(.a(s_15), .O(gate218inter4));
  nand2 gate650(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate651(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate652(.a(G627), .O(gate218inter7));
  inv1  gate653(.a(G678), .O(gate218inter8));
  nand2 gate654(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate655(.a(s_15), .b(gate218inter3), .O(gate218inter10));
  nor2  gate656(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate657(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate658(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1233(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1234(.a(gate219inter0), .b(s_98), .O(gate219inter1));
  and2  gate1235(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1236(.a(s_98), .O(gate219inter3));
  inv1  gate1237(.a(s_99), .O(gate219inter4));
  nand2 gate1238(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1239(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1240(.a(G632), .O(gate219inter7));
  inv1  gate1241(.a(G681), .O(gate219inter8));
  nand2 gate1242(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1243(.a(s_99), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1244(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1245(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1246(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate659(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate660(.a(gate222inter0), .b(s_16), .O(gate222inter1));
  and2  gate661(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate662(.a(s_16), .O(gate222inter3));
  inv1  gate663(.a(s_17), .O(gate222inter4));
  nand2 gate664(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate665(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate666(.a(G632), .O(gate222inter7));
  inv1  gate667(.a(G684), .O(gate222inter8));
  nand2 gate668(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate669(.a(s_17), .b(gate222inter3), .O(gate222inter10));
  nor2  gate670(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate671(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate672(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate729(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate730(.a(gate225inter0), .b(s_26), .O(gate225inter1));
  and2  gate731(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate732(.a(s_26), .O(gate225inter3));
  inv1  gate733(.a(s_27), .O(gate225inter4));
  nand2 gate734(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate735(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate736(.a(G690), .O(gate225inter7));
  inv1  gate737(.a(G691), .O(gate225inter8));
  nand2 gate738(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate739(.a(s_27), .b(gate225inter3), .O(gate225inter10));
  nor2  gate740(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate741(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate742(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2031(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2032(.a(gate227inter0), .b(s_212), .O(gate227inter1));
  and2  gate2033(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2034(.a(s_212), .O(gate227inter3));
  inv1  gate2035(.a(s_213), .O(gate227inter4));
  nand2 gate2036(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2037(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2038(.a(G694), .O(gate227inter7));
  inv1  gate2039(.a(G695), .O(gate227inter8));
  nand2 gate2040(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2041(.a(s_213), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2042(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2043(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2044(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2115(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2116(.a(gate229inter0), .b(s_224), .O(gate229inter1));
  and2  gate2117(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2118(.a(s_224), .O(gate229inter3));
  inv1  gate2119(.a(s_225), .O(gate229inter4));
  nand2 gate2120(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2121(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2122(.a(G698), .O(gate229inter7));
  inv1  gate2123(.a(G699), .O(gate229inter8));
  nand2 gate2124(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2125(.a(s_225), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2126(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2127(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2128(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1345(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1346(.a(gate235inter0), .b(s_114), .O(gate235inter1));
  and2  gate1347(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1348(.a(s_114), .O(gate235inter3));
  inv1  gate1349(.a(s_115), .O(gate235inter4));
  nand2 gate1350(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1351(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1352(.a(G248), .O(gate235inter7));
  inv1  gate1353(.a(G724), .O(gate235inter8));
  nand2 gate1354(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1355(.a(s_115), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1356(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1357(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1358(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1779(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1780(.a(gate248inter0), .b(s_176), .O(gate248inter1));
  and2  gate1781(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1782(.a(s_176), .O(gate248inter3));
  inv1  gate1783(.a(s_177), .O(gate248inter4));
  nand2 gate1784(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1785(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1786(.a(G727), .O(gate248inter7));
  inv1  gate1787(.a(G739), .O(gate248inter8));
  nand2 gate1788(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1789(.a(s_177), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1790(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1791(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1792(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate617(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate618(.a(gate251inter0), .b(s_10), .O(gate251inter1));
  and2  gate619(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate620(.a(s_10), .O(gate251inter3));
  inv1  gate621(.a(s_11), .O(gate251inter4));
  nand2 gate622(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate623(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate624(.a(G257), .O(gate251inter7));
  inv1  gate625(.a(G745), .O(gate251inter8));
  nand2 gate626(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate627(.a(s_11), .b(gate251inter3), .O(gate251inter10));
  nor2  gate628(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate629(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate630(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1513(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1514(.a(gate255inter0), .b(s_138), .O(gate255inter1));
  and2  gate1515(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1516(.a(s_138), .O(gate255inter3));
  inv1  gate1517(.a(s_139), .O(gate255inter4));
  nand2 gate1518(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1519(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1520(.a(G263), .O(gate255inter7));
  inv1  gate1521(.a(G751), .O(gate255inter8));
  nand2 gate1522(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1523(.a(s_139), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1524(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1525(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1526(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate785(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate786(.a(gate258inter0), .b(s_34), .O(gate258inter1));
  and2  gate787(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate788(.a(s_34), .O(gate258inter3));
  inv1  gate789(.a(s_35), .O(gate258inter4));
  nand2 gate790(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate791(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate792(.a(G756), .O(gate258inter7));
  inv1  gate793(.a(G757), .O(gate258inter8));
  nand2 gate794(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate795(.a(s_35), .b(gate258inter3), .O(gate258inter10));
  nor2  gate796(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate797(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate798(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1751(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1752(.a(gate260inter0), .b(s_172), .O(gate260inter1));
  and2  gate1753(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1754(.a(s_172), .O(gate260inter3));
  inv1  gate1755(.a(s_173), .O(gate260inter4));
  nand2 gate1756(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1757(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1758(.a(G760), .O(gate260inter7));
  inv1  gate1759(.a(G761), .O(gate260inter8));
  nand2 gate1760(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1761(.a(s_173), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1762(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1763(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1764(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1933(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1934(.a(gate264inter0), .b(s_198), .O(gate264inter1));
  and2  gate1935(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1936(.a(s_198), .O(gate264inter3));
  inv1  gate1937(.a(s_199), .O(gate264inter4));
  nand2 gate1938(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1939(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1940(.a(G768), .O(gate264inter7));
  inv1  gate1941(.a(G769), .O(gate264inter8));
  nand2 gate1942(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1943(.a(s_199), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1944(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1945(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1946(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1905(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1906(.a(gate267inter0), .b(s_194), .O(gate267inter1));
  and2  gate1907(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1908(.a(s_194), .O(gate267inter3));
  inv1  gate1909(.a(s_195), .O(gate267inter4));
  nand2 gate1910(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1911(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1912(.a(G648), .O(gate267inter7));
  inv1  gate1913(.a(G776), .O(gate267inter8));
  nand2 gate1914(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1915(.a(s_195), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1916(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1917(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1918(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate547(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate548(.a(gate270inter0), .b(s_0), .O(gate270inter1));
  and2  gate549(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate550(.a(s_0), .O(gate270inter3));
  inv1  gate551(.a(s_1), .O(gate270inter4));
  nand2 gate552(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate553(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate554(.a(G657), .O(gate270inter7));
  inv1  gate555(.a(G785), .O(gate270inter8));
  nand2 gate556(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate557(.a(s_1), .b(gate270inter3), .O(gate270inter10));
  nor2  gate558(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate559(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate560(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2143(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2144(.a(gate273inter0), .b(s_228), .O(gate273inter1));
  and2  gate2145(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2146(.a(s_228), .O(gate273inter3));
  inv1  gate2147(.a(s_229), .O(gate273inter4));
  nand2 gate2148(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2149(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2150(.a(G642), .O(gate273inter7));
  inv1  gate2151(.a(G794), .O(gate273inter8));
  nand2 gate2152(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2153(.a(s_229), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2154(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2155(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2156(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1191(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1192(.a(gate274inter0), .b(s_92), .O(gate274inter1));
  and2  gate1193(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1194(.a(s_92), .O(gate274inter3));
  inv1  gate1195(.a(s_93), .O(gate274inter4));
  nand2 gate1196(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1197(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1198(.a(G770), .O(gate274inter7));
  inv1  gate1199(.a(G794), .O(gate274inter8));
  nand2 gate1200(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1201(.a(s_93), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1202(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1203(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1204(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate575(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate576(.a(gate280inter0), .b(s_4), .O(gate280inter1));
  and2  gate577(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate578(.a(s_4), .O(gate280inter3));
  inv1  gate579(.a(s_5), .O(gate280inter4));
  nand2 gate580(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate581(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate582(.a(G779), .O(gate280inter7));
  inv1  gate583(.a(G803), .O(gate280inter8));
  nand2 gate584(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate585(.a(s_5), .b(gate280inter3), .O(gate280inter10));
  nor2  gate586(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate587(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate588(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1737(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1738(.a(gate283inter0), .b(s_170), .O(gate283inter1));
  and2  gate1739(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1740(.a(s_170), .O(gate283inter3));
  inv1  gate1741(.a(s_171), .O(gate283inter4));
  nand2 gate1742(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1743(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1744(.a(G657), .O(gate283inter7));
  inv1  gate1745(.a(G809), .O(gate283inter8));
  nand2 gate1746(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1747(.a(s_171), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1748(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1749(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1750(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1037(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1038(.a(gate288inter0), .b(s_70), .O(gate288inter1));
  and2  gate1039(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1040(.a(s_70), .O(gate288inter3));
  inv1  gate1041(.a(s_71), .O(gate288inter4));
  nand2 gate1042(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1043(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1044(.a(G791), .O(gate288inter7));
  inv1  gate1045(.a(G815), .O(gate288inter8));
  nand2 gate1046(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1047(.a(s_71), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1048(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1049(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1050(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1135(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1136(.a(gate289inter0), .b(s_84), .O(gate289inter1));
  and2  gate1137(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1138(.a(s_84), .O(gate289inter3));
  inv1  gate1139(.a(s_85), .O(gate289inter4));
  nand2 gate1140(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1141(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1142(.a(G818), .O(gate289inter7));
  inv1  gate1143(.a(G819), .O(gate289inter8));
  nand2 gate1144(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1145(.a(s_85), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1146(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1147(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1148(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1583(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1584(.a(gate290inter0), .b(s_148), .O(gate290inter1));
  and2  gate1585(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1586(.a(s_148), .O(gate290inter3));
  inv1  gate1587(.a(s_149), .O(gate290inter4));
  nand2 gate1588(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1589(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1590(.a(G820), .O(gate290inter7));
  inv1  gate1591(.a(G821), .O(gate290inter8));
  nand2 gate1592(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1593(.a(s_149), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1594(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1595(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1596(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1653(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1654(.a(gate293inter0), .b(s_158), .O(gate293inter1));
  and2  gate1655(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1656(.a(s_158), .O(gate293inter3));
  inv1  gate1657(.a(s_159), .O(gate293inter4));
  nand2 gate1658(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1659(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1660(.a(G828), .O(gate293inter7));
  inv1  gate1661(.a(G829), .O(gate293inter8));
  nand2 gate1662(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1663(.a(s_159), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1664(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1665(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1666(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1177(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1178(.a(gate401inter0), .b(s_90), .O(gate401inter1));
  and2  gate1179(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1180(.a(s_90), .O(gate401inter3));
  inv1  gate1181(.a(s_91), .O(gate401inter4));
  nand2 gate1182(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1183(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1184(.a(G15), .O(gate401inter7));
  inv1  gate1185(.a(G1078), .O(gate401inter8));
  nand2 gate1186(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1187(.a(s_91), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1188(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1189(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1190(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate981(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate982(.a(gate419inter0), .b(s_62), .O(gate419inter1));
  and2  gate983(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate984(.a(s_62), .O(gate419inter3));
  inv1  gate985(.a(s_63), .O(gate419inter4));
  nand2 gate986(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate987(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate988(.a(G1), .O(gate419inter7));
  inv1  gate989(.a(G1132), .O(gate419inter8));
  nand2 gate990(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate991(.a(s_63), .b(gate419inter3), .O(gate419inter10));
  nor2  gate992(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate993(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate994(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2157(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2158(.a(gate420inter0), .b(s_230), .O(gate420inter1));
  and2  gate2159(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2160(.a(s_230), .O(gate420inter3));
  inv1  gate2161(.a(s_231), .O(gate420inter4));
  nand2 gate2162(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2163(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2164(.a(G1036), .O(gate420inter7));
  inv1  gate2165(.a(G1132), .O(gate420inter8));
  nand2 gate2166(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2167(.a(s_231), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2168(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2169(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2170(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1499(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1500(.a(gate421inter0), .b(s_136), .O(gate421inter1));
  and2  gate1501(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1502(.a(s_136), .O(gate421inter3));
  inv1  gate1503(.a(s_137), .O(gate421inter4));
  nand2 gate1504(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1505(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1506(.a(G2), .O(gate421inter7));
  inv1  gate1507(.a(G1135), .O(gate421inter8));
  nand2 gate1508(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1509(.a(s_137), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1510(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1511(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1512(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate771(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate772(.a(gate422inter0), .b(s_32), .O(gate422inter1));
  and2  gate773(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate774(.a(s_32), .O(gate422inter3));
  inv1  gate775(.a(s_33), .O(gate422inter4));
  nand2 gate776(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate777(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate778(.a(G1039), .O(gate422inter7));
  inv1  gate779(.a(G1135), .O(gate422inter8));
  nand2 gate780(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate781(.a(s_33), .b(gate422inter3), .O(gate422inter10));
  nor2  gate782(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate783(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate784(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2003(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2004(.a(gate428inter0), .b(s_208), .O(gate428inter1));
  and2  gate2005(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2006(.a(s_208), .O(gate428inter3));
  inv1  gate2007(.a(s_209), .O(gate428inter4));
  nand2 gate2008(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2009(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2010(.a(G1048), .O(gate428inter7));
  inv1  gate2011(.a(G1144), .O(gate428inter8));
  nand2 gate2012(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2013(.a(s_209), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2014(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2015(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2016(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1247(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1248(.a(gate434inter0), .b(s_100), .O(gate434inter1));
  and2  gate1249(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1250(.a(s_100), .O(gate434inter3));
  inv1  gate1251(.a(s_101), .O(gate434inter4));
  nand2 gate1252(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1253(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1254(.a(G1057), .O(gate434inter7));
  inv1  gate1255(.a(G1153), .O(gate434inter8));
  nand2 gate1256(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1257(.a(s_101), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1258(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1259(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1260(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1989(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1990(.a(gate436inter0), .b(s_206), .O(gate436inter1));
  and2  gate1991(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1992(.a(s_206), .O(gate436inter3));
  inv1  gate1993(.a(s_207), .O(gate436inter4));
  nand2 gate1994(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1995(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1996(.a(G1060), .O(gate436inter7));
  inv1  gate1997(.a(G1156), .O(gate436inter8));
  nand2 gate1998(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1999(.a(s_207), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2000(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2001(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2002(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1275(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1276(.a(gate439inter0), .b(s_104), .O(gate439inter1));
  and2  gate1277(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1278(.a(s_104), .O(gate439inter3));
  inv1  gate1279(.a(s_105), .O(gate439inter4));
  nand2 gate1280(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1281(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1282(.a(G11), .O(gate439inter7));
  inv1  gate1283(.a(G1162), .O(gate439inter8));
  nand2 gate1284(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1285(.a(s_105), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1286(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1287(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1288(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1821(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1822(.a(gate441inter0), .b(s_182), .O(gate441inter1));
  and2  gate1823(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1824(.a(s_182), .O(gate441inter3));
  inv1  gate1825(.a(s_183), .O(gate441inter4));
  nand2 gate1826(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1827(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1828(.a(G12), .O(gate441inter7));
  inv1  gate1829(.a(G1165), .O(gate441inter8));
  nand2 gate1830(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1831(.a(s_183), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1832(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1833(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1834(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1163(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1164(.a(gate447inter0), .b(s_88), .O(gate447inter1));
  and2  gate1165(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1166(.a(s_88), .O(gate447inter3));
  inv1  gate1167(.a(s_89), .O(gate447inter4));
  nand2 gate1168(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1169(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1170(.a(G15), .O(gate447inter7));
  inv1  gate1171(.a(G1174), .O(gate447inter8));
  nand2 gate1172(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1173(.a(s_89), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1174(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1175(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1176(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1023(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1024(.a(gate451inter0), .b(s_68), .O(gate451inter1));
  and2  gate1025(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1026(.a(s_68), .O(gate451inter3));
  inv1  gate1027(.a(s_69), .O(gate451inter4));
  nand2 gate1028(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1029(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1030(.a(G17), .O(gate451inter7));
  inv1  gate1031(.a(G1180), .O(gate451inter8));
  nand2 gate1032(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1033(.a(s_69), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1034(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1035(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1036(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1107(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1108(.a(gate454inter0), .b(s_80), .O(gate454inter1));
  and2  gate1109(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1110(.a(s_80), .O(gate454inter3));
  inv1  gate1111(.a(s_81), .O(gate454inter4));
  nand2 gate1112(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1113(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1114(.a(G1087), .O(gate454inter7));
  inv1  gate1115(.a(G1183), .O(gate454inter8));
  nand2 gate1116(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1117(.a(s_81), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1118(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1119(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1120(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1695(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1696(.a(gate456inter0), .b(s_164), .O(gate456inter1));
  and2  gate1697(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1698(.a(s_164), .O(gate456inter3));
  inv1  gate1699(.a(s_165), .O(gate456inter4));
  nand2 gate1700(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1701(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1702(.a(G1090), .O(gate456inter7));
  inv1  gate1703(.a(G1186), .O(gate456inter8));
  nand2 gate1704(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1705(.a(s_165), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1706(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1707(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1708(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1205(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1206(.a(gate457inter0), .b(s_94), .O(gate457inter1));
  and2  gate1207(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1208(.a(s_94), .O(gate457inter3));
  inv1  gate1209(.a(s_95), .O(gate457inter4));
  nand2 gate1210(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1211(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1212(.a(G20), .O(gate457inter7));
  inv1  gate1213(.a(G1189), .O(gate457inter8));
  nand2 gate1214(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1215(.a(s_95), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1216(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1217(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1218(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1485(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1486(.a(gate458inter0), .b(s_134), .O(gate458inter1));
  and2  gate1487(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1488(.a(s_134), .O(gate458inter3));
  inv1  gate1489(.a(s_135), .O(gate458inter4));
  nand2 gate1490(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1491(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1492(.a(G1093), .O(gate458inter7));
  inv1  gate1493(.a(G1189), .O(gate458inter8));
  nand2 gate1494(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1495(.a(s_135), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1496(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1497(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1498(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2017(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2018(.a(gate463inter0), .b(s_210), .O(gate463inter1));
  and2  gate2019(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2020(.a(s_210), .O(gate463inter3));
  inv1  gate2021(.a(s_211), .O(gate463inter4));
  nand2 gate2022(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2023(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2024(.a(G23), .O(gate463inter7));
  inv1  gate2025(.a(G1198), .O(gate463inter8));
  nand2 gate2026(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2027(.a(s_211), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2028(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2029(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2030(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1597(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1598(.a(gate468inter0), .b(s_150), .O(gate468inter1));
  and2  gate1599(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1600(.a(s_150), .O(gate468inter3));
  inv1  gate1601(.a(s_151), .O(gate468inter4));
  nand2 gate1602(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1603(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1604(.a(G1108), .O(gate468inter7));
  inv1  gate1605(.a(G1204), .O(gate468inter8));
  nand2 gate1606(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1607(.a(s_151), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1608(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1609(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1610(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate953(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate954(.a(gate469inter0), .b(s_58), .O(gate469inter1));
  and2  gate955(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate956(.a(s_58), .O(gate469inter3));
  inv1  gate957(.a(s_59), .O(gate469inter4));
  nand2 gate958(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate959(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate960(.a(G26), .O(gate469inter7));
  inv1  gate961(.a(G1207), .O(gate469inter8));
  nand2 gate962(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate963(.a(s_59), .b(gate469inter3), .O(gate469inter10));
  nor2  gate964(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate965(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate966(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1961(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1962(.a(gate476inter0), .b(s_202), .O(gate476inter1));
  and2  gate1963(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1964(.a(s_202), .O(gate476inter3));
  inv1  gate1965(.a(s_203), .O(gate476inter4));
  nand2 gate1966(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1967(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1968(.a(G1120), .O(gate476inter7));
  inv1  gate1969(.a(G1216), .O(gate476inter8));
  nand2 gate1970(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1971(.a(s_203), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1972(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1973(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1974(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1149(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1150(.a(gate481inter0), .b(s_86), .O(gate481inter1));
  and2  gate1151(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1152(.a(s_86), .O(gate481inter3));
  inv1  gate1153(.a(s_87), .O(gate481inter4));
  nand2 gate1154(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1155(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1156(.a(G32), .O(gate481inter7));
  inv1  gate1157(.a(G1225), .O(gate481inter8));
  nand2 gate1158(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1159(.a(s_87), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1160(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1161(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1162(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1373(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1374(.a(gate483inter0), .b(s_118), .O(gate483inter1));
  and2  gate1375(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1376(.a(s_118), .O(gate483inter3));
  inv1  gate1377(.a(s_119), .O(gate483inter4));
  nand2 gate1378(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1379(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1380(.a(G1228), .O(gate483inter7));
  inv1  gate1381(.a(G1229), .O(gate483inter8));
  nand2 gate1382(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1383(.a(s_119), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1384(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1385(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1386(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2059(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2060(.a(gate486inter0), .b(s_216), .O(gate486inter1));
  and2  gate2061(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2062(.a(s_216), .O(gate486inter3));
  inv1  gate2063(.a(s_217), .O(gate486inter4));
  nand2 gate2064(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2065(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2066(.a(G1234), .O(gate486inter7));
  inv1  gate2067(.a(G1235), .O(gate486inter8));
  nand2 gate2068(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2069(.a(s_217), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2070(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2071(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2072(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1667(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1668(.a(gate487inter0), .b(s_160), .O(gate487inter1));
  and2  gate1669(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1670(.a(s_160), .O(gate487inter3));
  inv1  gate1671(.a(s_161), .O(gate487inter4));
  nand2 gate1672(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1673(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1674(.a(G1236), .O(gate487inter7));
  inv1  gate1675(.a(G1237), .O(gate487inter8));
  nand2 gate1676(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1677(.a(s_161), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1678(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1679(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1680(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate631(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate632(.a(gate488inter0), .b(s_12), .O(gate488inter1));
  and2  gate633(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate634(.a(s_12), .O(gate488inter3));
  inv1  gate635(.a(s_13), .O(gate488inter4));
  nand2 gate636(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate637(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate638(.a(G1238), .O(gate488inter7));
  inv1  gate639(.a(G1239), .O(gate488inter8));
  nand2 gate640(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate641(.a(s_13), .b(gate488inter3), .O(gate488inter10));
  nor2  gate642(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate643(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate644(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate855(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate856(.a(gate490inter0), .b(s_44), .O(gate490inter1));
  and2  gate857(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate858(.a(s_44), .O(gate490inter3));
  inv1  gate859(.a(s_45), .O(gate490inter4));
  nand2 gate860(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate861(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate862(.a(G1242), .O(gate490inter7));
  inv1  gate863(.a(G1243), .O(gate490inter8));
  nand2 gate864(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate865(.a(s_45), .b(gate490inter3), .O(gate490inter10));
  nor2  gate866(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate867(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate868(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1079(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1080(.a(gate494inter0), .b(s_76), .O(gate494inter1));
  and2  gate1081(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1082(.a(s_76), .O(gate494inter3));
  inv1  gate1083(.a(s_77), .O(gate494inter4));
  nand2 gate1084(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1085(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1086(.a(G1250), .O(gate494inter7));
  inv1  gate1087(.a(G1251), .O(gate494inter8));
  nand2 gate1088(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1089(.a(s_77), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1090(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1091(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1092(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1541(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1542(.a(gate496inter0), .b(s_142), .O(gate496inter1));
  and2  gate1543(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1544(.a(s_142), .O(gate496inter3));
  inv1  gate1545(.a(s_143), .O(gate496inter4));
  nand2 gate1546(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1547(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1548(.a(G1254), .O(gate496inter7));
  inv1  gate1549(.a(G1255), .O(gate496inter8));
  nand2 gate1550(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1551(.a(s_143), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1552(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1553(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1554(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1009(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1010(.a(gate497inter0), .b(s_66), .O(gate497inter1));
  and2  gate1011(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1012(.a(s_66), .O(gate497inter3));
  inv1  gate1013(.a(s_67), .O(gate497inter4));
  nand2 gate1014(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1015(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1016(.a(G1256), .O(gate497inter7));
  inv1  gate1017(.a(G1257), .O(gate497inter8));
  nand2 gate1018(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1019(.a(s_67), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1020(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1021(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1022(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1569(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1570(.a(gate499inter0), .b(s_146), .O(gate499inter1));
  and2  gate1571(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1572(.a(s_146), .O(gate499inter3));
  inv1  gate1573(.a(s_147), .O(gate499inter4));
  nand2 gate1574(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1575(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1576(.a(G1260), .O(gate499inter7));
  inv1  gate1577(.a(G1261), .O(gate499inter8));
  nand2 gate1578(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1579(.a(s_147), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1580(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1581(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1582(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate603(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate604(.a(gate501inter0), .b(s_8), .O(gate501inter1));
  and2  gate605(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate606(.a(s_8), .O(gate501inter3));
  inv1  gate607(.a(s_9), .O(gate501inter4));
  nand2 gate608(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate609(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate610(.a(G1264), .O(gate501inter7));
  inv1  gate611(.a(G1265), .O(gate501inter8));
  nand2 gate612(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate613(.a(s_9), .b(gate501inter3), .O(gate501inter10));
  nor2  gate614(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate615(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate616(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate561(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate562(.a(gate503inter0), .b(s_2), .O(gate503inter1));
  and2  gate563(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate564(.a(s_2), .O(gate503inter3));
  inv1  gate565(.a(s_3), .O(gate503inter4));
  nand2 gate566(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate567(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate568(.a(G1268), .O(gate503inter7));
  inv1  gate569(.a(G1269), .O(gate503inter8));
  nand2 gate570(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate571(.a(s_3), .b(gate503inter3), .O(gate503inter10));
  nor2  gate572(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate573(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate574(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1317(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1318(.a(gate504inter0), .b(s_110), .O(gate504inter1));
  and2  gate1319(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1320(.a(s_110), .O(gate504inter3));
  inv1  gate1321(.a(s_111), .O(gate504inter4));
  nand2 gate1322(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1323(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1324(.a(G1270), .O(gate504inter7));
  inv1  gate1325(.a(G1271), .O(gate504inter8));
  nand2 gate1326(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1327(.a(s_111), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1328(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1329(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1330(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1303(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1304(.a(gate505inter0), .b(s_108), .O(gate505inter1));
  and2  gate1305(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1306(.a(s_108), .O(gate505inter3));
  inv1  gate1307(.a(s_109), .O(gate505inter4));
  nand2 gate1308(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1309(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1310(.a(G1272), .O(gate505inter7));
  inv1  gate1311(.a(G1273), .O(gate505inter8));
  nand2 gate1312(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1313(.a(s_109), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1314(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1315(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1316(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1877(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1878(.a(gate511inter0), .b(s_190), .O(gate511inter1));
  and2  gate1879(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1880(.a(s_190), .O(gate511inter3));
  inv1  gate1881(.a(s_191), .O(gate511inter4));
  nand2 gate1882(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1883(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1884(.a(G1284), .O(gate511inter7));
  inv1  gate1885(.a(G1285), .O(gate511inter8));
  nand2 gate1886(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1887(.a(s_191), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1888(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1889(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1890(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule