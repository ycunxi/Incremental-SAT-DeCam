module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
input s_382,s_383;//RE__ALLOW(00,01,10,11);
input s_384,s_385;//RE__ALLOW(00,01,10,11);
input s_386,s_387;//RE__ALLOW(00,01,10,11);
input s_388,s_389;//RE__ALLOW(00,01,10,11);
input s_390,s_391;//RE__ALLOW(00,01,10,11);
input s_392,s_393;//RE__ALLOW(00,01,10,11);
input s_394,s_395;//RE__ALLOW(00,01,10,11);
input s_396,s_397;//RE__ALLOW(00,01,10,11);
input s_398,s_399;//RE__ALLOW(00,01,10,11);
input s_400,s_401;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate995(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate996(.a(gate9inter0), .b(s_64), .O(gate9inter1));
  and2  gate997(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate998(.a(s_64), .O(gate9inter3));
  inv1  gate999(.a(s_65), .O(gate9inter4));
  nand2 gate1000(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1001(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1002(.a(G1), .O(gate9inter7));
  inv1  gate1003(.a(G2), .O(gate9inter8));
  nand2 gate1004(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1005(.a(s_65), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1006(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1007(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1008(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2829(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2830(.a(gate15inter0), .b(s_326), .O(gate15inter1));
  and2  gate2831(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2832(.a(s_326), .O(gate15inter3));
  inv1  gate2833(.a(s_327), .O(gate15inter4));
  nand2 gate2834(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2835(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2836(.a(G13), .O(gate15inter7));
  inv1  gate2837(.a(G14), .O(gate15inter8));
  nand2 gate2838(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2839(.a(s_327), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2840(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2841(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2842(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2619(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2620(.a(gate21inter0), .b(s_296), .O(gate21inter1));
  and2  gate2621(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2622(.a(s_296), .O(gate21inter3));
  inv1  gate2623(.a(s_297), .O(gate21inter4));
  nand2 gate2624(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2625(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2626(.a(G25), .O(gate21inter7));
  inv1  gate2627(.a(G26), .O(gate21inter8));
  nand2 gate2628(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2629(.a(s_297), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2630(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2631(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2632(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate3179(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate3180(.a(gate25inter0), .b(s_376), .O(gate25inter1));
  and2  gate3181(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate3182(.a(s_376), .O(gate25inter3));
  inv1  gate3183(.a(s_377), .O(gate25inter4));
  nand2 gate3184(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate3185(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate3186(.a(G1), .O(gate25inter7));
  inv1  gate3187(.a(G5), .O(gate25inter8));
  nand2 gate3188(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate3189(.a(s_377), .b(gate25inter3), .O(gate25inter10));
  nor2  gate3190(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate3191(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate3192(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2577(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2578(.a(gate29inter0), .b(s_290), .O(gate29inter1));
  and2  gate2579(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2580(.a(s_290), .O(gate29inter3));
  inv1  gate2581(.a(s_291), .O(gate29inter4));
  nand2 gate2582(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2583(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2584(.a(G3), .O(gate29inter7));
  inv1  gate2585(.a(G7), .O(gate29inter8));
  nand2 gate2586(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2587(.a(s_291), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2588(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2589(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2590(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2941(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2942(.a(gate31inter0), .b(s_342), .O(gate31inter1));
  and2  gate2943(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2944(.a(s_342), .O(gate31inter3));
  inv1  gate2945(.a(s_343), .O(gate31inter4));
  nand2 gate2946(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2947(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2948(.a(G4), .O(gate31inter7));
  inv1  gate2949(.a(G8), .O(gate31inter8));
  nand2 gate2950(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2951(.a(s_343), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2952(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2953(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2954(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2003(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2004(.a(gate34inter0), .b(s_208), .O(gate34inter1));
  and2  gate2005(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2006(.a(s_208), .O(gate34inter3));
  inv1  gate2007(.a(s_209), .O(gate34inter4));
  nand2 gate2008(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2009(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2010(.a(G25), .O(gate34inter7));
  inv1  gate2011(.a(G29), .O(gate34inter8));
  nand2 gate2012(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2013(.a(s_209), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2014(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2015(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2016(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1219(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1220(.a(gate35inter0), .b(s_96), .O(gate35inter1));
  and2  gate1221(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1222(.a(s_96), .O(gate35inter3));
  inv1  gate1223(.a(s_97), .O(gate35inter4));
  nand2 gate1224(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1225(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1226(.a(G18), .O(gate35inter7));
  inv1  gate1227(.a(G22), .O(gate35inter8));
  nand2 gate1228(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1229(.a(s_97), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1230(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1231(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1232(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1303(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1304(.a(gate36inter0), .b(s_108), .O(gate36inter1));
  and2  gate1305(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1306(.a(s_108), .O(gate36inter3));
  inv1  gate1307(.a(s_109), .O(gate36inter4));
  nand2 gate1308(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1309(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1310(.a(G26), .O(gate36inter7));
  inv1  gate1311(.a(G30), .O(gate36inter8));
  nand2 gate1312(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1313(.a(s_109), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1314(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1315(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1316(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2465(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2466(.a(gate40inter0), .b(s_274), .O(gate40inter1));
  and2  gate2467(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2468(.a(s_274), .O(gate40inter3));
  inv1  gate2469(.a(s_275), .O(gate40inter4));
  nand2 gate2470(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2471(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2472(.a(G28), .O(gate40inter7));
  inv1  gate2473(.a(G32), .O(gate40inter8));
  nand2 gate2474(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2475(.a(s_275), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2476(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2477(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2478(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate3053(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate3054(.a(gate46inter0), .b(s_358), .O(gate46inter1));
  and2  gate3055(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate3056(.a(s_358), .O(gate46inter3));
  inv1  gate3057(.a(s_359), .O(gate46inter4));
  nand2 gate3058(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate3059(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate3060(.a(G6), .O(gate46inter7));
  inv1  gate3061(.a(G272), .O(gate46inter8));
  nand2 gate3062(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate3063(.a(s_359), .b(gate46inter3), .O(gate46inter10));
  nor2  gate3064(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate3065(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate3066(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1289(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1290(.a(gate48inter0), .b(s_106), .O(gate48inter1));
  and2  gate1291(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1292(.a(s_106), .O(gate48inter3));
  inv1  gate1293(.a(s_107), .O(gate48inter4));
  nand2 gate1294(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1295(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1296(.a(G8), .O(gate48inter7));
  inv1  gate1297(.a(G275), .O(gate48inter8));
  nand2 gate1298(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1299(.a(s_107), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1300(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1301(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1302(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate3095(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate3096(.a(gate50inter0), .b(s_364), .O(gate50inter1));
  and2  gate3097(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate3098(.a(s_364), .O(gate50inter3));
  inv1  gate3099(.a(s_365), .O(gate50inter4));
  nand2 gate3100(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate3101(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate3102(.a(G10), .O(gate50inter7));
  inv1  gate3103(.a(G278), .O(gate50inter8));
  nand2 gate3104(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate3105(.a(s_365), .b(gate50inter3), .O(gate50inter10));
  nor2  gate3106(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate3107(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate3108(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2171(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2172(.a(gate51inter0), .b(s_232), .O(gate51inter1));
  and2  gate2173(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2174(.a(s_232), .O(gate51inter3));
  inv1  gate2175(.a(s_233), .O(gate51inter4));
  nand2 gate2176(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2177(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2178(.a(G11), .O(gate51inter7));
  inv1  gate2179(.a(G281), .O(gate51inter8));
  nand2 gate2180(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2181(.a(s_233), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2182(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2183(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2184(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1681(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1682(.a(gate52inter0), .b(s_162), .O(gate52inter1));
  and2  gate1683(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1684(.a(s_162), .O(gate52inter3));
  inv1  gate1685(.a(s_163), .O(gate52inter4));
  nand2 gate1686(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1687(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1688(.a(G12), .O(gate52inter7));
  inv1  gate1689(.a(G281), .O(gate52inter8));
  nand2 gate1690(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1691(.a(s_163), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1692(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1693(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1694(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2255(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2256(.a(gate54inter0), .b(s_244), .O(gate54inter1));
  and2  gate2257(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2258(.a(s_244), .O(gate54inter3));
  inv1  gate2259(.a(s_245), .O(gate54inter4));
  nand2 gate2260(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2261(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2262(.a(G14), .O(gate54inter7));
  inv1  gate2263(.a(G284), .O(gate54inter8));
  nand2 gate2264(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2265(.a(s_245), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2266(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2267(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2268(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2857(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2858(.a(gate56inter0), .b(s_330), .O(gate56inter1));
  and2  gate2859(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2860(.a(s_330), .O(gate56inter3));
  inv1  gate2861(.a(s_331), .O(gate56inter4));
  nand2 gate2862(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2863(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2864(.a(G16), .O(gate56inter7));
  inv1  gate2865(.a(G287), .O(gate56inter8));
  nand2 gate2866(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2867(.a(s_331), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2868(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2869(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2870(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1583(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1584(.a(gate57inter0), .b(s_148), .O(gate57inter1));
  and2  gate1585(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1586(.a(s_148), .O(gate57inter3));
  inv1  gate1587(.a(s_149), .O(gate57inter4));
  nand2 gate1588(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1589(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1590(.a(G17), .O(gate57inter7));
  inv1  gate1591(.a(G290), .O(gate57inter8));
  nand2 gate1592(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1593(.a(s_149), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1594(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1595(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1596(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2479(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2480(.a(gate59inter0), .b(s_276), .O(gate59inter1));
  and2  gate2481(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2482(.a(s_276), .O(gate59inter3));
  inv1  gate2483(.a(s_277), .O(gate59inter4));
  nand2 gate2484(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2485(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2486(.a(G19), .O(gate59inter7));
  inv1  gate2487(.a(G293), .O(gate59inter8));
  nand2 gate2488(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2489(.a(s_277), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2490(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2491(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2492(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate561(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate562(.a(gate61inter0), .b(s_2), .O(gate61inter1));
  and2  gate563(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate564(.a(s_2), .O(gate61inter3));
  inv1  gate565(.a(s_3), .O(gate61inter4));
  nand2 gate566(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate567(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate568(.a(G21), .O(gate61inter7));
  inv1  gate569(.a(G296), .O(gate61inter8));
  nand2 gate570(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate571(.a(s_3), .b(gate61inter3), .O(gate61inter10));
  nor2  gate572(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate573(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate574(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1835(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1836(.a(gate63inter0), .b(s_184), .O(gate63inter1));
  and2  gate1837(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1838(.a(s_184), .O(gate63inter3));
  inv1  gate1839(.a(s_185), .O(gate63inter4));
  nand2 gate1840(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1841(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1842(.a(G23), .O(gate63inter7));
  inv1  gate1843(.a(G299), .O(gate63inter8));
  nand2 gate1844(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1845(.a(s_185), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1846(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1847(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1848(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1933(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1934(.a(gate64inter0), .b(s_198), .O(gate64inter1));
  and2  gate1935(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1936(.a(s_198), .O(gate64inter3));
  inv1  gate1937(.a(s_199), .O(gate64inter4));
  nand2 gate1938(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1939(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1940(.a(G24), .O(gate64inter7));
  inv1  gate1941(.a(G299), .O(gate64inter8));
  nand2 gate1942(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1943(.a(s_199), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1944(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1945(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1946(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2899(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2900(.a(gate66inter0), .b(s_336), .O(gate66inter1));
  and2  gate2901(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2902(.a(s_336), .O(gate66inter3));
  inv1  gate2903(.a(s_337), .O(gate66inter4));
  nand2 gate2904(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2905(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2906(.a(G26), .O(gate66inter7));
  inv1  gate2907(.a(G302), .O(gate66inter8));
  nand2 gate2908(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2909(.a(s_337), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2910(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2911(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2912(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate2199(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2200(.a(gate67inter0), .b(s_236), .O(gate67inter1));
  and2  gate2201(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2202(.a(s_236), .O(gate67inter3));
  inv1  gate2203(.a(s_237), .O(gate67inter4));
  nand2 gate2204(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2205(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2206(.a(G27), .O(gate67inter7));
  inv1  gate2207(.a(G305), .O(gate67inter8));
  nand2 gate2208(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2209(.a(s_237), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2210(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2211(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2212(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2129(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2130(.a(gate70inter0), .b(s_226), .O(gate70inter1));
  and2  gate2131(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2132(.a(s_226), .O(gate70inter3));
  inv1  gate2133(.a(s_227), .O(gate70inter4));
  nand2 gate2134(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2135(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2136(.a(G30), .O(gate70inter7));
  inv1  gate2137(.a(G308), .O(gate70inter8));
  nand2 gate2138(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2139(.a(s_227), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2140(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2141(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2142(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1695(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1696(.a(gate74inter0), .b(s_164), .O(gate74inter1));
  and2  gate1697(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1698(.a(s_164), .O(gate74inter3));
  inv1  gate1699(.a(s_165), .O(gate74inter4));
  nand2 gate1700(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1701(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1702(.a(G5), .O(gate74inter7));
  inv1  gate1703(.a(G314), .O(gate74inter8));
  nand2 gate1704(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1705(.a(s_165), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1706(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1707(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1708(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate785(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate786(.a(gate75inter0), .b(s_34), .O(gate75inter1));
  and2  gate787(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate788(.a(s_34), .O(gate75inter3));
  inv1  gate789(.a(s_35), .O(gate75inter4));
  nand2 gate790(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate791(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate792(.a(G9), .O(gate75inter7));
  inv1  gate793(.a(G317), .O(gate75inter8));
  nand2 gate794(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate795(.a(s_35), .b(gate75inter3), .O(gate75inter10));
  nor2  gate796(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate797(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate798(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate3109(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate3110(.a(gate77inter0), .b(s_366), .O(gate77inter1));
  and2  gate3111(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate3112(.a(s_366), .O(gate77inter3));
  inv1  gate3113(.a(s_367), .O(gate77inter4));
  nand2 gate3114(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate3115(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate3116(.a(G2), .O(gate77inter7));
  inv1  gate3117(.a(G320), .O(gate77inter8));
  nand2 gate3118(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate3119(.a(s_367), .b(gate77inter3), .O(gate77inter10));
  nor2  gate3120(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate3121(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate3122(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2787(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2788(.a(gate79inter0), .b(s_320), .O(gate79inter1));
  and2  gate2789(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2790(.a(s_320), .O(gate79inter3));
  inv1  gate2791(.a(s_321), .O(gate79inter4));
  nand2 gate2792(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2793(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2794(.a(G10), .O(gate79inter7));
  inv1  gate2795(.a(G323), .O(gate79inter8));
  nand2 gate2796(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2797(.a(s_321), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2798(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2799(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2800(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate617(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate618(.a(gate81inter0), .b(s_10), .O(gate81inter1));
  and2  gate619(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate620(.a(s_10), .O(gate81inter3));
  inv1  gate621(.a(s_11), .O(gate81inter4));
  nand2 gate622(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate623(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate624(.a(G3), .O(gate81inter7));
  inv1  gate625(.a(G326), .O(gate81inter8));
  nand2 gate626(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate627(.a(s_11), .b(gate81inter3), .O(gate81inter10));
  nor2  gate628(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate629(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate630(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2409(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2410(.a(gate88inter0), .b(s_266), .O(gate88inter1));
  and2  gate2411(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2412(.a(s_266), .O(gate88inter3));
  inv1  gate2413(.a(s_267), .O(gate88inter4));
  nand2 gate2414(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2415(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2416(.a(G16), .O(gate88inter7));
  inv1  gate2417(.a(G335), .O(gate88inter8));
  nand2 gate2418(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2419(.a(s_267), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2420(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2421(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2422(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate3039(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate3040(.a(gate89inter0), .b(s_356), .O(gate89inter1));
  and2  gate3041(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate3042(.a(s_356), .O(gate89inter3));
  inv1  gate3043(.a(s_357), .O(gate89inter4));
  nand2 gate3044(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate3045(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate3046(.a(G17), .O(gate89inter7));
  inv1  gate3047(.a(G338), .O(gate89inter8));
  nand2 gate3048(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate3049(.a(s_357), .b(gate89inter3), .O(gate89inter10));
  nor2  gate3050(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate3051(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate3052(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate631(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate632(.a(gate100inter0), .b(s_12), .O(gate100inter1));
  and2  gate633(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate634(.a(s_12), .O(gate100inter3));
  inv1  gate635(.a(s_13), .O(gate100inter4));
  nand2 gate636(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate637(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate638(.a(G31), .O(gate100inter7));
  inv1  gate639(.a(G353), .O(gate100inter8));
  nand2 gate640(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate641(.a(s_13), .b(gate100inter3), .O(gate100inter10));
  nor2  gate642(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate643(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate644(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1331(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1332(.a(gate101inter0), .b(s_112), .O(gate101inter1));
  and2  gate1333(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1334(.a(s_112), .O(gate101inter3));
  inv1  gate1335(.a(s_113), .O(gate101inter4));
  nand2 gate1336(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1337(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1338(.a(G20), .O(gate101inter7));
  inv1  gate1339(.a(G356), .O(gate101inter8));
  nand2 gate1340(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1341(.a(s_113), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1342(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1343(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1344(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate3333(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate3334(.a(gate103inter0), .b(s_398), .O(gate103inter1));
  and2  gate3335(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate3336(.a(s_398), .O(gate103inter3));
  inv1  gate3337(.a(s_399), .O(gate103inter4));
  nand2 gate3338(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate3339(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate3340(.a(G28), .O(gate103inter7));
  inv1  gate3341(.a(G359), .O(gate103inter8));
  nand2 gate3342(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate3343(.a(s_399), .b(gate103inter3), .O(gate103inter10));
  nor2  gate3344(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate3345(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate3346(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1429(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1430(.a(gate104inter0), .b(s_126), .O(gate104inter1));
  and2  gate1431(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1432(.a(s_126), .O(gate104inter3));
  inv1  gate1433(.a(s_127), .O(gate104inter4));
  nand2 gate1434(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1435(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1436(.a(G32), .O(gate104inter7));
  inv1  gate1437(.a(G359), .O(gate104inter8));
  nand2 gate1438(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1439(.a(s_127), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1440(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1441(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1442(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate3263(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate3264(.a(gate106inter0), .b(s_388), .O(gate106inter1));
  and2  gate3265(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate3266(.a(s_388), .O(gate106inter3));
  inv1  gate3267(.a(s_389), .O(gate106inter4));
  nand2 gate3268(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate3269(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate3270(.a(G364), .O(gate106inter7));
  inv1  gate3271(.a(G365), .O(gate106inter8));
  nand2 gate3272(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate3273(.a(s_389), .b(gate106inter3), .O(gate106inter10));
  nor2  gate3274(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate3275(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate3276(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2661(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2662(.a(gate112inter0), .b(s_302), .O(gate112inter1));
  and2  gate2663(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2664(.a(s_302), .O(gate112inter3));
  inv1  gate2665(.a(s_303), .O(gate112inter4));
  nand2 gate2666(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2667(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2668(.a(G376), .O(gate112inter7));
  inv1  gate2669(.a(G377), .O(gate112inter8));
  nand2 gate2670(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2671(.a(s_303), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2672(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2673(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2674(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate3235(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate3236(.a(gate115inter0), .b(s_384), .O(gate115inter1));
  and2  gate3237(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate3238(.a(s_384), .O(gate115inter3));
  inv1  gate3239(.a(s_385), .O(gate115inter4));
  nand2 gate3240(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate3241(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate3242(.a(G382), .O(gate115inter7));
  inv1  gate3243(.a(G383), .O(gate115inter8));
  nand2 gate3244(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate3245(.a(s_385), .b(gate115inter3), .O(gate115inter10));
  nor2  gate3246(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate3247(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate3248(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2241(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2242(.a(gate117inter0), .b(s_242), .O(gate117inter1));
  and2  gate2243(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2244(.a(s_242), .O(gate117inter3));
  inv1  gate2245(.a(s_243), .O(gate117inter4));
  nand2 gate2246(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2247(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2248(.a(G386), .O(gate117inter7));
  inv1  gate2249(.a(G387), .O(gate117inter8));
  nand2 gate2250(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2251(.a(s_243), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2252(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2253(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2254(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1317(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1318(.a(gate123inter0), .b(s_110), .O(gate123inter1));
  and2  gate1319(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1320(.a(s_110), .O(gate123inter3));
  inv1  gate1321(.a(s_111), .O(gate123inter4));
  nand2 gate1322(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1323(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1324(.a(G398), .O(gate123inter7));
  inv1  gate1325(.a(G399), .O(gate123inter8));
  nand2 gate1326(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1327(.a(s_111), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1328(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1329(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1330(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate2773(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2774(.a(gate124inter0), .b(s_318), .O(gate124inter1));
  and2  gate2775(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2776(.a(s_318), .O(gate124inter3));
  inv1  gate2777(.a(s_319), .O(gate124inter4));
  nand2 gate2778(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2779(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2780(.a(G400), .O(gate124inter7));
  inv1  gate2781(.a(G401), .O(gate124inter8));
  nand2 gate2782(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2783(.a(s_319), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2784(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2785(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2786(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1779(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1780(.a(gate125inter0), .b(s_176), .O(gate125inter1));
  and2  gate1781(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1782(.a(s_176), .O(gate125inter3));
  inv1  gate1783(.a(s_177), .O(gate125inter4));
  nand2 gate1784(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1785(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1786(.a(G402), .O(gate125inter7));
  inv1  gate1787(.a(G403), .O(gate125inter8));
  nand2 gate1788(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1789(.a(s_177), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1790(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1791(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1792(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate939(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate940(.a(gate126inter0), .b(s_56), .O(gate126inter1));
  and2  gate941(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate942(.a(s_56), .O(gate126inter3));
  inv1  gate943(.a(s_57), .O(gate126inter4));
  nand2 gate944(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate945(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate946(.a(G404), .O(gate126inter7));
  inv1  gate947(.a(G405), .O(gate126inter8));
  nand2 gate948(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate949(.a(s_57), .b(gate126inter3), .O(gate126inter10));
  nor2  gate950(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate951(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate952(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1891(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1892(.a(gate127inter0), .b(s_192), .O(gate127inter1));
  and2  gate1893(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1894(.a(s_192), .O(gate127inter3));
  inv1  gate1895(.a(s_193), .O(gate127inter4));
  nand2 gate1896(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1897(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1898(.a(G406), .O(gate127inter7));
  inv1  gate1899(.a(G407), .O(gate127inter8));
  nand2 gate1900(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1901(.a(s_193), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1902(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1903(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1904(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1121(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1122(.a(gate128inter0), .b(s_82), .O(gate128inter1));
  and2  gate1123(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1124(.a(s_82), .O(gate128inter3));
  inv1  gate1125(.a(s_83), .O(gate128inter4));
  nand2 gate1126(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1127(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1128(.a(G408), .O(gate128inter7));
  inv1  gate1129(.a(G409), .O(gate128inter8));
  nand2 gate1130(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1131(.a(s_83), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1132(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1133(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1134(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate3221(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate3222(.a(gate130inter0), .b(s_382), .O(gate130inter1));
  and2  gate3223(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate3224(.a(s_382), .O(gate130inter3));
  inv1  gate3225(.a(s_383), .O(gate130inter4));
  nand2 gate3226(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate3227(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate3228(.a(G412), .O(gate130inter7));
  inv1  gate3229(.a(G413), .O(gate130inter8));
  nand2 gate3230(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate3231(.a(s_383), .b(gate130inter3), .O(gate130inter10));
  nor2  gate3232(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate3233(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate3234(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2955(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2956(.a(gate135inter0), .b(s_344), .O(gate135inter1));
  and2  gate2957(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2958(.a(s_344), .O(gate135inter3));
  inv1  gate2959(.a(s_345), .O(gate135inter4));
  nand2 gate2960(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2961(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2962(.a(G422), .O(gate135inter7));
  inv1  gate2963(.a(G423), .O(gate135inter8));
  nand2 gate2964(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2965(.a(s_345), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2966(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2967(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2968(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1373(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1374(.a(gate136inter0), .b(s_118), .O(gate136inter1));
  and2  gate1375(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1376(.a(s_118), .O(gate136inter3));
  inv1  gate1377(.a(s_119), .O(gate136inter4));
  nand2 gate1378(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1379(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1380(.a(G424), .O(gate136inter7));
  inv1  gate1381(.a(G425), .O(gate136inter8));
  nand2 gate1382(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1383(.a(s_119), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1384(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1385(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1386(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2101(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2102(.a(gate137inter0), .b(s_222), .O(gate137inter1));
  and2  gate2103(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2104(.a(s_222), .O(gate137inter3));
  inv1  gate2105(.a(s_223), .O(gate137inter4));
  nand2 gate2106(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2107(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2108(.a(G426), .O(gate137inter7));
  inv1  gate2109(.a(G429), .O(gate137inter8));
  nand2 gate2110(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2111(.a(s_223), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2112(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2113(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2114(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate3347(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate3348(.a(gate138inter0), .b(s_400), .O(gate138inter1));
  and2  gate3349(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate3350(.a(s_400), .O(gate138inter3));
  inv1  gate3351(.a(s_401), .O(gate138inter4));
  nand2 gate3352(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate3353(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate3354(.a(G432), .O(gate138inter7));
  inv1  gate3355(.a(G435), .O(gate138inter8));
  nand2 gate3356(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate3357(.a(s_401), .b(gate138inter3), .O(gate138inter10));
  nor2  gate3358(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate3359(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate3360(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1975(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1976(.a(gate140inter0), .b(s_204), .O(gate140inter1));
  and2  gate1977(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1978(.a(s_204), .O(gate140inter3));
  inv1  gate1979(.a(s_205), .O(gate140inter4));
  nand2 gate1980(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1981(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1982(.a(G444), .O(gate140inter7));
  inv1  gate1983(.a(G447), .O(gate140inter8));
  nand2 gate1984(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1985(.a(s_205), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1986(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1987(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1988(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2437(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2438(.a(gate143inter0), .b(s_270), .O(gate143inter1));
  and2  gate2439(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2440(.a(s_270), .O(gate143inter3));
  inv1  gate2441(.a(s_271), .O(gate143inter4));
  nand2 gate2442(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2443(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2444(.a(G462), .O(gate143inter7));
  inv1  gate2445(.a(G465), .O(gate143inter8));
  nand2 gate2446(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2447(.a(s_271), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2448(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2449(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2450(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2675(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2676(.a(gate146inter0), .b(s_304), .O(gate146inter1));
  and2  gate2677(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2678(.a(s_304), .O(gate146inter3));
  inv1  gate2679(.a(s_305), .O(gate146inter4));
  nand2 gate2680(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2681(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2682(.a(G480), .O(gate146inter7));
  inv1  gate2683(.a(G483), .O(gate146inter8));
  nand2 gate2684(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2685(.a(s_305), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2686(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2687(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2688(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1597(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1598(.a(gate148inter0), .b(s_150), .O(gate148inter1));
  and2  gate1599(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1600(.a(s_150), .O(gate148inter3));
  inv1  gate1601(.a(s_151), .O(gate148inter4));
  nand2 gate1602(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1603(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1604(.a(G492), .O(gate148inter7));
  inv1  gate1605(.a(G495), .O(gate148inter8));
  nand2 gate1606(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1607(.a(s_151), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1608(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1609(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1610(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2647(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2648(.a(gate153inter0), .b(s_300), .O(gate153inter1));
  and2  gate2649(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2650(.a(s_300), .O(gate153inter3));
  inv1  gate2651(.a(s_301), .O(gate153inter4));
  nand2 gate2652(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2653(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2654(.a(G426), .O(gate153inter7));
  inv1  gate2655(.a(G522), .O(gate153inter8));
  nand2 gate2656(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2657(.a(s_301), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2658(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2659(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2660(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2563(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2564(.a(gate155inter0), .b(s_288), .O(gate155inter1));
  and2  gate2565(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2566(.a(s_288), .O(gate155inter3));
  inv1  gate2567(.a(s_289), .O(gate155inter4));
  nand2 gate2568(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2569(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2570(.a(G432), .O(gate155inter7));
  inv1  gate2571(.a(G525), .O(gate155inter8));
  nand2 gate2572(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2573(.a(s_289), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2574(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2575(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2576(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2815(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2816(.a(gate157inter0), .b(s_324), .O(gate157inter1));
  and2  gate2817(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2818(.a(s_324), .O(gate157inter3));
  inv1  gate2819(.a(s_325), .O(gate157inter4));
  nand2 gate2820(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2821(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2822(.a(G438), .O(gate157inter7));
  inv1  gate2823(.a(G528), .O(gate157inter8));
  nand2 gate2824(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2825(.a(s_325), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2826(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2827(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2828(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2367(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2368(.a(gate158inter0), .b(s_260), .O(gate158inter1));
  and2  gate2369(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2370(.a(s_260), .O(gate158inter3));
  inv1  gate2371(.a(s_261), .O(gate158inter4));
  nand2 gate2372(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2373(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2374(.a(G441), .O(gate158inter7));
  inv1  gate2375(.a(G528), .O(gate158inter8));
  nand2 gate2376(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2377(.a(s_261), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2378(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2379(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2380(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1653(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1654(.a(gate159inter0), .b(s_158), .O(gate159inter1));
  and2  gate1655(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1656(.a(s_158), .O(gate159inter3));
  inv1  gate1657(.a(s_159), .O(gate159inter4));
  nand2 gate1658(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1659(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1660(.a(G444), .O(gate159inter7));
  inv1  gate1661(.a(G531), .O(gate159inter8));
  nand2 gate1662(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1663(.a(s_159), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1664(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1665(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1666(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate911(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate912(.a(gate160inter0), .b(s_52), .O(gate160inter1));
  and2  gate913(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate914(.a(s_52), .O(gate160inter3));
  inv1  gate915(.a(s_53), .O(gate160inter4));
  nand2 gate916(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate917(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate918(.a(G447), .O(gate160inter7));
  inv1  gate919(.a(G531), .O(gate160inter8));
  nand2 gate920(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate921(.a(s_53), .b(gate160inter3), .O(gate160inter10));
  nor2  gate922(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate923(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate924(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1261(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1262(.a(gate162inter0), .b(s_102), .O(gate162inter1));
  and2  gate1263(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1264(.a(s_102), .O(gate162inter3));
  inv1  gate1265(.a(s_103), .O(gate162inter4));
  nand2 gate1266(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1267(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1268(.a(G453), .O(gate162inter7));
  inv1  gate1269(.a(G534), .O(gate162inter8));
  nand2 gate1270(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1271(.a(s_103), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1272(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1273(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1274(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2087(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2088(.a(gate163inter0), .b(s_220), .O(gate163inter1));
  and2  gate2089(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2090(.a(s_220), .O(gate163inter3));
  inv1  gate2091(.a(s_221), .O(gate163inter4));
  nand2 gate2092(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2093(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2094(.a(G456), .O(gate163inter7));
  inv1  gate2095(.a(G537), .O(gate163inter8));
  nand2 gate2096(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2097(.a(s_221), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2098(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2099(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2100(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1709(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1710(.a(gate169inter0), .b(s_166), .O(gate169inter1));
  and2  gate1711(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1712(.a(s_166), .O(gate169inter3));
  inv1  gate1713(.a(s_167), .O(gate169inter4));
  nand2 gate1714(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1715(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1716(.a(G474), .O(gate169inter7));
  inv1  gate1717(.a(G546), .O(gate169inter8));
  nand2 gate1718(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1719(.a(s_167), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1720(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1721(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1722(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2045(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2046(.a(gate173inter0), .b(s_214), .O(gate173inter1));
  and2  gate2047(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2048(.a(s_214), .O(gate173inter3));
  inv1  gate2049(.a(s_215), .O(gate173inter4));
  nand2 gate2050(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2051(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2052(.a(G486), .O(gate173inter7));
  inv1  gate2053(.a(G552), .O(gate173inter8));
  nand2 gate2054(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2055(.a(s_215), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2056(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2057(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2058(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2535(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2536(.a(gate176inter0), .b(s_284), .O(gate176inter1));
  and2  gate2537(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2538(.a(s_284), .O(gate176inter3));
  inv1  gate2539(.a(s_285), .O(gate176inter4));
  nand2 gate2540(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2541(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2542(.a(G495), .O(gate176inter7));
  inv1  gate2543(.a(G555), .O(gate176inter8));
  nand2 gate2544(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2545(.a(s_285), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2546(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2547(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2548(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1093(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1094(.a(gate178inter0), .b(s_78), .O(gate178inter1));
  and2  gate1095(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1096(.a(s_78), .O(gate178inter3));
  inv1  gate1097(.a(s_79), .O(gate178inter4));
  nand2 gate1098(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1099(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1100(.a(G501), .O(gate178inter7));
  inv1  gate1101(.a(G558), .O(gate178inter8));
  nand2 gate1102(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1103(.a(s_79), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1104(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1105(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1106(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate715(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate716(.a(gate179inter0), .b(s_24), .O(gate179inter1));
  and2  gate717(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate718(.a(s_24), .O(gate179inter3));
  inv1  gate719(.a(s_25), .O(gate179inter4));
  nand2 gate720(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate721(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate722(.a(G504), .O(gate179inter7));
  inv1  gate723(.a(G561), .O(gate179inter8));
  nand2 gate724(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate725(.a(s_25), .b(gate179inter3), .O(gate179inter10));
  nor2  gate726(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate727(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate728(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2017(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2018(.a(gate181inter0), .b(s_210), .O(gate181inter1));
  and2  gate2019(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2020(.a(s_210), .O(gate181inter3));
  inv1  gate2021(.a(s_211), .O(gate181inter4));
  nand2 gate2022(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2023(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2024(.a(G510), .O(gate181inter7));
  inv1  gate2025(.a(G564), .O(gate181inter8));
  nand2 gate2026(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2027(.a(s_211), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2028(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2029(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2030(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1247(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1248(.a(gate184inter0), .b(s_100), .O(gate184inter1));
  and2  gate1249(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1250(.a(s_100), .O(gate184inter3));
  inv1  gate1251(.a(s_101), .O(gate184inter4));
  nand2 gate1252(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1253(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1254(.a(G519), .O(gate184inter7));
  inv1  gate1255(.a(G567), .O(gate184inter8));
  nand2 gate1256(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1257(.a(s_101), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1258(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1259(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1260(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate3305(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate3306(.a(gate187inter0), .b(s_394), .O(gate187inter1));
  and2  gate3307(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate3308(.a(s_394), .O(gate187inter3));
  inv1  gate3309(.a(s_395), .O(gate187inter4));
  nand2 gate3310(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate3311(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate3312(.a(G574), .O(gate187inter7));
  inv1  gate3313(.a(G575), .O(gate187inter8));
  nand2 gate3314(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate3315(.a(s_395), .b(gate187inter3), .O(gate187inter10));
  nor2  gate3316(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate3317(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate3318(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1541(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1542(.a(gate188inter0), .b(s_142), .O(gate188inter1));
  and2  gate1543(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1544(.a(s_142), .O(gate188inter3));
  inv1  gate1545(.a(s_143), .O(gate188inter4));
  nand2 gate1546(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1547(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1548(.a(G576), .O(gate188inter7));
  inv1  gate1549(.a(G577), .O(gate188inter8));
  nand2 gate1550(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1551(.a(s_143), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1552(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1553(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1554(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2983(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2984(.a(gate189inter0), .b(s_348), .O(gate189inter1));
  and2  gate2985(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2986(.a(s_348), .O(gate189inter3));
  inv1  gate2987(.a(s_349), .O(gate189inter4));
  nand2 gate2988(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2989(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2990(.a(G578), .O(gate189inter7));
  inv1  gate2991(.a(G579), .O(gate189inter8));
  nand2 gate2992(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2993(.a(s_349), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2994(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2995(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2996(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1821(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1822(.a(gate191inter0), .b(s_182), .O(gate191inter1));
  and2  gate1823(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1824(.a(s_182), .O(gate191inter3));
  inv1  gate1825(.a(s_183), .O(gate191inter4));
  nand2 gate1826(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1827(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1828(.a(G582), .O(gate191inter7));
  inv1  gate1829(.a(G583), .O(gate191inter8));
  nand2 gate1830(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1831(.a(s_183), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1832(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1833(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1834(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1345(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1346(.a(gate194inter0), .b(s_114), .O(gate194inter1));
  and2  gate1347(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1348(.a(s_114), .O(gate194inter3));
  inv1  gate1349(.a(s_115), .O(gate194inter4));
  nand2 gate1350(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1351(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1352(.a(G588), .O(gate194inter7));
  inv1  gate1353(.a(G589), .O(gate194inter8));
  nand2 gate1354(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1355(.a(s_115), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1356(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1357(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1358(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2073(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2074(.a(gate195inter0), .b(s_218), .O(gate195inter1));
  and2  gate2075(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2076(.a(s_218), .O(gate195inter3));
  inv1  gate2077(.a(s_219), .O(gate195inter4));
  nand2 gate2078(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2079(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2080(.a(G590), .O(gate195inter7));
  inv1  gate2081(.a(G591), .O(gate195inter8));
  nand2 gate2082(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2083(.a(s_219), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2084(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2085(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2086(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate589(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate590(.a(gate197inter0), .b(s_6), .O(gate197inter1));
  and2  gate591(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate592(.a(s_6), .O(gate197inter3));
  inv1  gate593(.a(s_7), .O(gate197inter4));
  nand2 gate594(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate595(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate596(.a(G594), .O(gate197inter7));
  inv1  gate597(.a(G595), .O(gate197inter8));
  nand2 gate598(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate599(.a(s_7), .b(gate197inter3), .O(gate197inter10));
  nor2  gate600(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate601(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate602(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate3011(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate3012(.a(gate202inter0), .b(s_352), .O(gate202inter1));
  and2  gate3013(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate3014(.a(s_352), .O(gate202inter3));
  inv1  gate3015(.a(s_353), .O(gate202inter4));
  nand2 gate3016(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate3017(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate3018(.a(G612), .O(gate202inter7));
  inv1  gate3019(.a(G617), .O(gate202inter8));
  nand2 gate3020(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate3021(.a(s_353), .b(gate202inter3), .O(gate202inter10));
  nor2  gate3022(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate3023(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate3024(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate925(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate926(.a(gate204inter0), .b(s_54), .O(gate204inter1));
  and2  gate927(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate928(.a(s_54), .O(gate204inter3));
  inv1  gate929(.a(s_55), .O(gate204inter4));
  nand2 gate930(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate931(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate932(.a(G607), .O(gate204inter7));
  inv1  gate933(.a(G617), .O(gate204inter8));
  nand2 gate934(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate935(.a(s_55), .b(gate204inter3), .O(gate204inter10));
  nor2  gate936(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate937(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate938(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate2997(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2998(.a(gate205inter0), .b(s_350), .O(gate205inter1));
  and2  gate2999(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate3000(.a(s_350), .O(gate205inter3));
  inv1  gate3001(.a(s_351), .O(gate205inter4));
  nand2 gate3002(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate3003(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate3004(.a(G622), .O(gate205inter7));
  inv1  gate3005(.a(G627), .O(gate205inter8));
  nand2 gate3006(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate3007(.a(s_351), .b(gate205inter3), .O(gate205inter10));
  nor2  gate3008(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate3009(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate3010(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2423(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2424(.a(gate206inter0), .b(s_268), .O(gate206inter1));
  and2  gate2425(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2426(.a(s_268), .O(gate206inter3));
  inv1  gate2427(.a(s_269), .O(gate206inter4));
  nand2 gate2428(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2429(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2430(.a(G632), .O(gate206inter7));
  inv1  gate2431(.a(G637), .O(gate206inter8));
  nand2 gate2432(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2433(.a(s_269), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2434(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2435(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2436(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2381(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2382(.a(gate207inter0), .b(s_262), .O(gate207inter1));
  and2  gate2383(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2384(.a(s_262), .O(gate207inter3));
  inv1  gate2385(.a(s_263), .O(gate207inter4));
  nand2 gate2386(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2387(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2388(.a(G622), .O(gate207inter7));
  inv1  gate2389(.a(G632), .O(gate207inter8));
  nand2 gate2390(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2391(.a(s_263), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2392(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2393(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2394(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1163(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1164(.a(gate208inter0), .b(s_88), .O(gate208inter1));
  and2  gate1165(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1166(.a(s_88), .O(gate208inter3));
  inv1  gate1167(.a(s_89), .O(gate208inter4));
  nand2 gate1168(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1169(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1170(.a(G627), .O(gate208inter7));
  inv1  gate1171(.a(G637), .O(gate208inter8));
  nand2 gate1172(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1173(.a(s_89), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1174(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1175(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1176(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1569(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1570(.a(gate210inter0), .b(s_146), .O(gate210inter1));
  and2  gate1571(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1572(.a(s_146), .O(gate210inter3));
  inv1  gate1573(.a(s_147), .O(gate210inter4));
  nand2 gate1574(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1575(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1576(.a(G607), .O(gate210inter7));
  inv1  gate1577(.a(G666), .O(gate210inter8));
  nand2 gate1578(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1579(.a(s_147), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1580(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1581(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1582(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1919(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1920(.a(gate212inter0), .b(s_196), .O(gate212inter1));
  and2  gate1921(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1922(.a(s_196), .O(gate212inter3));
  inv1  gate1923(.a(s_197), .O(gate212inter4));
  nand2 gate1924(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1925(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1926(.a(G617), .O(gate212inter7));
  inv1  gate1927(.a(G669), .O(gate212inter8));
  nand2 gate1928(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1929(.a(s_197), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1930(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1931(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1932(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1275(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1276(.a(gate214inter0), .b(s_104), .O(gate214inter1));
  and2  gate1277(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1278(.a(s_104), .O(gate214inter3));
  inv1  gate1279(.a(s_105), .O(gate214inter4));
  nand2 gate1280(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1281(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1282(.a(G612), .O(gate214inter7));
  inv1  gate1283(.a(G672), .O(gate214inter8));
  nand2 gate1284(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1285(.a(s_105), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1286(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1287(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1288(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate981(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate982(.a(gate215inter0), .b(s_62), .O(gate215inter1));
  and2  gate983(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate984(.a(s_62), .O(gate215inter3));
  inv1  gate985(.a(s_63), .O(gate215inter4));
  nand2 gate986(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate987(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate988(.a(G607), .O(gate215inter7));
  inv1  gate989(.a(G675), .O(gate215inter8));
  nand2 gate990(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate991(.a(s_63), .b(gate215inter3), .O(gate215inter10));
  nor2  gate992(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate993(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate994(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate2717(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2718(.a(gate216inter0), .b(s_310), .O(gate216inter1));
  and2  gate2719(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2720(.a(s_310), .O(gate216inter3));
  inv1  gate2721(.a(s_311), .O(gate216inter4));
  nand2 gate2722(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2723(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2724(.a(G617), .O(gate216inter7));
  inv1  gate2725(.a(G675), .O(gate216inter8));
  nand2 gate2726(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2727(.a(s_311), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2728(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2729(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2730(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1457(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1458(.a(gate217inter0), .b(s_130), .O(gate217inter1));
  and2  gate1459(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1460(.a(s_130), .O(gate217inter3));
  inv1  gate1461(.a(s_131), .O(gate217inter4));
  nand2 gate1462(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1463(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1464(.a(G622), .O(gate217inter7));
  inv1  gate1465(.a(G678), .O(gate217inter8));
  nand2 gate1466(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1467(.a(s_131), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1468(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1469(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1470(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1723(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1724(.a(gate218inter0), .b(s_168), .O(gate218inter1));
  and2  gate1725(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1726(.a(s_168), .O(gate218inter3));
  inv1  gate1727(.a(s_169), .O(gate218inter4));
  nand2 gate1728(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1729(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1730(.a(G627), .O(gate218inter7));
  inv1  gate1731(.a(G678), .O(gate218inter8));
  nand2 gate1732(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1733(.a(s_169), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1734(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1735(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1736(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate3165(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate3166(.a(gate220inter0), .b(s_374), .O(gate220inter1));
  and2  gate3167(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate3168(.a(s_374), .O(gate220inter3));
  inv1  gate3169(.a(s_375), .O(gate220inter4));
  nand2 gate3170(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate3171(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate3172(.a(G637), .O(gate220inter7));
  inv1  gate3173(.a(G681), .O(gate220inter8));
  nand2 gate3174(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate3175(.a(s_375), .b(gate220inter3), .O(gate220inter10));
  nor2  gate3176(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate3177(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate3178(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1135(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1136(.a(gate221inter0), .b(s_84), .O(gate221inter1));
  and2  gate1137(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1138(.a(s_84), .O(gate221inter3));
  inv1  gate1139(.a(s_85), .O(gate221inter4));
  nand2 gate1140(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1141(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1142(.a(G622), .O(gate221inter7));
  inv1  gate1143(.a(G684), .O(gate221inter8));
  nand2 gate1144(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1145(.a(s_85), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1146(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1147(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1148(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1387(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1388(.a(gate222inter0), .b(s_120), .O(gate222inter1));
  and2  gate1389(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1390(.a(s_120), .O(gate222inter3));
  inv1  gate1391(.a(s_121), .O(gate222inter4));
  nand2 gate1392(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1393(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1394(.a(G632), .O(gate222inter7));
  inv1  gate1395(.a(G684), .O(gate222inter8));
  nand2 gate1396(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1397(.a(s_121), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1398(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1399(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1400(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2115(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2116(.a(gate224inter0), .b(s_224), .O(gate224inter1));
  and2  gate2117(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2118(.a(s_224), .O(gate224inter3));
  inv1  gate2119(.a(s_225), .O(gate224inter4));
  nand2 gate2120(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2121(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2122(.a(G637), .O(gate224inter7));
  inv1  gate2123(.a(G687), .O(gate224inter8));
  nand2 gate2124(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2125(.a(s_225), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2126(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2127(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2128(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1359(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1360(.a(gate226inter0), .b(s_116), .O(gate226inter1));
  and2  gate1361(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1362(.a(s_116), .O(gate226inter3));
  inv1  gate1363(.a(s_117), .O(gate226inter4));
  nand2 gate1364(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1365(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1366(.a(G692), .O(gate226inter7));
  inv1  gate1367(.a(G693), .O(gate226inter8));
  nand2 gate1368(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1369(.a(s_117), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1370(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1371(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1372(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate2605(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2606(.a(gate227inter0), .b(s_294), .O(gate227inter1));
  and2  gate2607(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2608(.a(s_294), .O(gate227inter3));
  inv1  gate2609(.a(s_295), .O(gate227inter4));
  nand2 gate2610(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2611(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2612(.a(G694), .O(gate227inter7));
  inv1  gate2613(.a(G695), .O(gate227inter8));
  nand2 gate2614(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2615(.a(s_295), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2616(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2617(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2618(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate841(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate842(.a(gate228inter0), .b(s_42), .O(gate228inter1));
  and2  gate843(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate844(.a(s_42), .O(gate228inter3));
  inv1  gate845(.a(s_43), .O(gate228inter4));
  nand2 gate846(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate847(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate848(.a(G696), .O(gate228inter7));
  inv1  gate849(.a(G697), .O(gate228inter8));
  nand2 gate850(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate851(.a(s_43), .b(gate228inter3), .O(gate228inter10));
  nor2  gate852(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate853(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate854(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1863(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1864(.a(gate229inter0), .b(s_188), .O(gate229inter1));
  and2  gate1865(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1866(.a(s_188), .O(gate229inter3));
  inv1  gate1867(.a(s_189), .O(gate229inter4));
  nand2 gate1868(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1869(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1870(.a(G698), .O(gate229inter7));
  inv1  gate1871(.a(G699), .O(gate229inter8));
  nand2 gate1872(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1873(.a(s_189), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1874(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1875(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1876(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate967(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate968(.a(gate233inter0), .b(s_60), .O(gate233inter1));
  and2  gate969(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate970(.a(s_60), .O(gate233inter3));
  inv1  gate971(.a(s_61), .O(gate233inter4));
  nand2 gate972(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate973(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate974(.a(G242), .O(gate233inter7));
  inv1  gate975(.a(G718), .O(gate233inter8));
  nand2 gate976(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate977(.a(s_61), .b(gate233inter3), .O(gate233inter10));
  nor2  gate978(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate979(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate980(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate813(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate814(.a(gate238inter0), .b(s_38), .O(gate238inter1));
  and2  gate815(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate816(.a(s_38), .O(gate238inter3));
  inv1  gate817(.a(s_39), .O(gate238inter4));
  nand2 gate818(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate819(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate820(.a(G257), .O(gate238inter7));
  inv1  gate821(.a(G709), .O(gate238inter8));
  nand2 gate822(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate823(.a(s_39), .b(gate238inter3), .O(gate238inter10));
  nor2  gate824(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate825(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate826(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1401(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1402(.a(gate240inter0), .b(s_122), .O(gate240inter1));
  and2  gate1403(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1404(.a(s_122), .O(gate240inter3));
  inv1  gate1405(.a(s_123), .O(gate240inter4));
  nand2 gate1406(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1407(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1408(.a(G263), .O(gate240inter7));
  inv1  gate1409(.a(G715), .O(gate240inter8));
  nand2 gate1410(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1411(.a(s_123), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1412(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1413(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1414(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1471(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1472(.a(gate242inter0), .b(s_132), .O(gate242inter1));
  and2  gate1473(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1474(.a(s_132), .O(gate242inter3));
  inv1  gate1475(.a(s_133), .O(gate242inter4));
  nand2 gate1476(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1477(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1478(.a(G718), .O(gate242inter7));
  inv1  gate1479(.a(G730), .O(gate242inter8));
  nand2 gate1480(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1481(.a(s_133), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1482(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1483(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1484(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate2297(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2298(.a(gate243inter0), .b(s_250), .O(gate243inter1));
  and2  gate2299(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2300(.a(s_250), .O(gate243inter3));
  inv1  gate2301(.a(s_251), .O(gate243inter4));
  nand2 gate2302(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2303(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2304(.a(G245), .O(gate243inter7));
  inv1  gate2305(.a(G733), .O(gate243inter8));
  nand2 gate2306(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2307(.a(s_251), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2308(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2309(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2310(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate757(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate758(.a(gate244inter0), .b(s_30), .O(gate244inter1));
  and2  gate759(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate760(.a(s_30), .O(gate244inter3));
  inv1  gate761(.a(s_31), .O(gate244inter4));
  nand2 gate762(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate763(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate764(.a(G721), .O(gate244inter7));
  inv1  gate765(.a(G733), .O(gate244inter8));
  nand2 gate766(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate767(.a(s_31), .b(gate244inter3), .O(gate244inter10));
  nor2  gate768(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate769(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate770(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1989(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1990(.a(gate245inter0), .b(s_206), .O(gate245inter1));
  and2  gate1991(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1992(.a(s_206), .O(gate245inter3));
  inv1  gate1993(.a(s_207), .O(gate245inter4));
  nand2 gate1994(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1995(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1996(.a(G248), .O(gate245inter7));
  inv1  gate1997(.a(G736), .O(gate245inter8));
  nand2 gate1998(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1999(.a(s_207), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2000(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2001(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2002(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate3081(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate3082(.a(gate248inter0), .b(s_362), .O(gate248inter1));
  and2  gate3083(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate3084(.a(s_362), .O(gate248inter3));
  inv1  gate3085(.a(s_363), .O(gate248inter4));
  nand2 gate3086(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate3087(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate3088(.a(G727), .O(gate248inter7));
  inv1  gate3089(.a(G739), .O(gate248inter8));
  nand2 gate3090(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate3091(.a(s_363), .b(gate248inter3), .O(gate248inter10));
  nor2  gate3092(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate3093(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate3094(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1737(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1738(.a(gate249inter0), .b(s_170), .O(gate249inter1));
  and2  gate1739(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1740(.a(s_170), .O(gate249inter3));
  inv1  gate1741(.a(s_171), .O(gate249inter4));
  nand2 gate1742(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1743(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1744(.a(G254), .O(gate249inter7));
  inv1  gate1745(.a(G742), .O(gate249inter8));
  nand2 gate1746(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1747(.a(s_171), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1748(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1749(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1750(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2927(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2928(.a(gate252inter0), .b(s_340), .O(gate252inter1));
  and2  gate2929(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2930(.a(s_340), .O(gate252inter3));
  inv1  gate2931(.a(s_341), .O(gate252inter4));
  nand2 gate2932(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2933(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2934(.a(G709), .O(gate252inter7));
  inv1  gate2935(.a(G745), .O(gate252inter8));
  nand2 gate2936(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2937(.a(s_341), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2938(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2939(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2940(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1191(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1192(.a(gate254inter0), .b(s_92), .O(gate254inter1));
  and2  gate1193(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1194(.a(s_92), .O(gate254inter3));
  inv1  gate1195(.a(s_93), .O(gate254inter4));
  nand2 gate1196(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1197(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1198(.a(G712), .O(gate254inter7));
  inv1  gate1199(.a(G748), .O(gate254inter8));
  nand2 gate1200(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1201(.a(s_93), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1202(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1203(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1204(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1177(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1178(.a(gate255inter0), .b(s_90), .O(gate255inter1));
  and2  gate1179(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1180(.a(s_90), .O(gate255inter3));
  inv1  gate1181(.a(s_91), .O(gate255inter4));
  nand2 gate1182(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1183(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1184(.a(G263), .O(gate255inter7));
  inv1  gate1185(.a(G751), .O(gate255inter8));
  nand2 gate1186(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1187(.a(s_91), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1188(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1189(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1190(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1765(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1766(.a(gate259inter0), .b(s_174), .O(gate259inter1));
  and2  gate1767(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1768(.a(s_174), .O(gate259inter3));
  inv1  gate1769(.a(s_175), .O(gate259inter4));
  nand2 gate1770(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1771(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1772(.a(G758), .O(gate259inter7));
  inv1  gate1773(.a(G759), .O(gate259inter8));
  nand2 gate1774(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1775(.a(s_175), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1776(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1777(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1778(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1947(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1948(.a(gate260inter0), .b(s_200), .O(gate260inter1));
  and2  gate1949(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1950(.a(s_200), .O(gate260inter3));
  inv1  gate1951(.a(s_201), .O(gate260inter4));
  nand2 gate1952(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1953(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1954(.a(G760), .O(gate260inter7));
  inv1  gate1955(.a(G761), .O(gate260inter8));
  nand2 gate1956(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1957(.a(s_201), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1958(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1959(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1960(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate3025(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate3026(.a(gate261inter0), .b(s_354), .O(gate261inter1));
  and2  gate3027(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate3028(.a(s_354), .O(gate261inter3));
  inv1  gate3029(.a(s_355), .O(gate261inter4));
  nand2 gate3030(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate3031(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate3032(.a(G762), .O(gate261inter7));
  inv1  gate3033(.a(G763), .O(gate261inter8));
  nand2 gate3034(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate3035(.a(s_355), .b(gate261inter3), .O(gate261inter10));
  nor2  gate3036(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate3037(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate3038(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate3137(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate3138(.a(gate262inter0), .b(s_370), .O(gate262inter1));
  and2  gate3139(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate3140(.a(s_370), .O(gate262inter3));
  inv1  gate3141(.a(s_371), .O(gate262inter4));
  nand2 gate3142(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate3143(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate3144(.a(G764), .O(gate262inter7));
  inv1  gate3145(.a(G765), .O(gate262inter8));
  nand2 gate3146(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate3147(.a(s_371), .b(gate262inter3), .O(gate262inter10));
  nor2  gate3148(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate3149(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate3150(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate869(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate870(.a(gate263inter0), .b(s_46), .O(gate263inter1));
  and2  gate871(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate872(.a(s_46), .O(gate263inter3));
  inv1  gate873(.a(s_47), .O(gate263inter4));
  nand2 gate874(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate875(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate876(.a(G766), .O(gate263inter7));
  inv1  gate877(.a(G767), .O(gate263inter8));
  nand2 gate878(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate879(.a(s_47), .b(gate263inter3), .O(gate263inter10));
  nor2  gate880(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate881(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate882(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1807(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1808(.a(gate264inter0), .b(s_180), .O(gate264inter1));
  and2  gate1809(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1810(.a(s_180), .O(gate264inter3));
  inv1  gate1811(.a(s_181), .O(gate264inter4));
  nand2 gate1812(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1813(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1814(.a(G768), .O(gate264inter7));
  inv1  gate1815(.a(G769), .O(gate264inter8));
  nand2 gate1816(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1817(.a(s_181), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1818(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1819(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1820(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1485(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1486(.a(gate265inter0), .b(s_134), .O(gate265inter1));
  and2  gate1487(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1488(.a(s_134), .O(gate265inter3));
  inv1  gate1489(.a(s_135), .O(gate265inter4));
  nand2 gate1490(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1491(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1492(.a(G642), .O(gate265inter7));
  inv1  gate1493(.a(G770), .O(gate265inter8));
  nand2 gate1494(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1495(.a(s_135), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1496(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1497(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1498(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1877(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1878(.a(gate266inter0), .b(s_190), .O(gate266inter1));
  and2  gate1879(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1880(.a(s_190), .O(gate266inter3));
  inv1  gate1881(.a(s_191), .O(gate266inter4));
  nand2 gate1882(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1883(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1884(.a(G645), .O(gate266inter7));
  inv1  gate1885(.a(G773), .O(gate266inter8));
  nand2 gate1886(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1887(.a(s_191), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1888(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1889(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1890(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1513(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1514(.a(gate269inter0), .b(s_138), .O(gate269inter1));
  and2  gate1515(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1516(.a(s_138), .O(gate269inter3));
  inv1  gate1517(.a(s_139), .O(gate269inter4));
  nand2 gate1518(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1519(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1520(.a(G654), .O(gate269inter7));
  inv1  gate1521(.a(G782), .O(gate269inter8));
  nand2 gate1522(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1523(.a(s_139), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1524(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1525(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1526(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate883(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate884(.a(gate270inter0), .b(s_48), .O(gate270inter1));
  and2  gate885(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate886(.a(s_48), .O(gate270inter3));
  inv1  gate887(.a(s_49), .O(gate270inter4));
  nand2 gate888(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate889(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate890(.a(G657), .O(gate270inter7));
  inv1  gate891(.a(G785), .O(gate270inter8));
  nand2 gate892(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate893(.a(s_49), .b(gate270inter3), .O(gate270inter10));
  nor2  gate894(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate895(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate896(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate687(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate688(.a(gate271inter0), .b(s_20), .O(gate271inter1));
  and2  gate689(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate690(.a(s_20), .O(gate271inter3));
  inv1  gate691(.a(s_21), .O(gate271inter4));
  nand2 gate692(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate693(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate694(.a(G660), .O(gate271inter7));
  inv1  gate695(.a(G788), .O(gate271inter8));
  nand2 gate696(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate697(.a(s_21), .b(gate271inter3), .O(gate271inter10));
  nor2  gate698(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate699(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate700(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2311(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2312(.a(gate273inter0), .b(s_252), .O(gate273inter1));
  and2  gate2313(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2314(.a(s_252), .O(gate273inter3));
  inv1  gate2315(.a(s_253), .O(gate273inter4));
  nand2 gate2316(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2317(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2318(.a(G642), .O(gate273inter7));
  inv1  gate2319(.a(G794), .O(gate273inter8));
  nand2 gate2320(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2321(.a(s_253), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2322(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2323(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2324(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2689(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2690(.a(gate278inter0), .b(s_306), .O(gate278inter1));
  and2  gate2691(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2692(.a(s_306), .O(gate278inter3));
  inv1  gate2693(.a(s_307), .O(gate278inter4));
  nand2 gate2694(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2695(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2696(.a(G776), .O(gate278inter7));
  inv1  gate2697(.a(G800), .O(gate278inter8));
  nand2 gate2698(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2699(.a(s_307), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2700(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2701(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2702(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate2143(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2144(.a(gate279inter0), .b(s_228), .O(gate279inter1));
  and2  gate2145(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2146(.a(s_228), .O(gate279inter3));
  inv1  gate2147(.a(s_229), .O(gate279inter4));
  nand2 gate2148(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2149(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2150(.a(G651), .O(gate279inter7));
  inv1  gate2151(.a(G803), .O(gate279inter8));
  nand2 gate2152(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2153(.a(s_229), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2154(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2155(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2156(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate2633(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2634(.a(gate280inter0), .b(s_298), .O(gate280inter1));
  and2  gate2635(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2636(.a(s_298), .O(gate280inter3));
  inv1  gate2637(.a(s_299), .O(gate280inter4));
  nand2 gate2638(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2639(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2640(.a(G779), .O(gate280inter7));
  inv1  gate2641(.a(G803), .O(gate280inter8));
  nand2 gate2642(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2643(.a(s_299), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2644(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2645(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2646(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1009(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1010(.a(gate281inter0), .b(s_66), .O(gate281inter1));
  and2  gate1011(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1012(.a(s_66), .O(gate281inter3));
  inv1  gate1013(.a(s_67), .O(gate281inter4));
  nand2 gate1014(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1015(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1016(.a(G654), .O(gate281inter7));
  inv1  gate1017(.a(G806), .O(gate281inter8));
  nand2 gate1018(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1019(.a(s_67), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1020(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1021(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1022(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate729(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate730(.a(gate282inter0), .b(s_26), .O(gate282inter1));
  and2  gate731(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate732(.a(s_26), .O(gate282inter3));
  inv1  gate733(.a(s_27), .O(gate282inter4));
  nand2 gate734(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate735(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate736(.a(G782), .O(gate282inter7));
  inv1  gate737(.a(G806), .O(gate282inter8));
  nand2 gate738(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate739(.a(s_27), .b(gate282inter3), .O(gate282inter10));
  nor2  gate740(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate741(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate742(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate575(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate576(.a(gate283inter0), .b(s_4), .O(gate283inter1));
  and2  gate577(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate578(.a(s_4), .O(gate283inter3));
  inv1  gate579(.a(s_5), .O(gate283inter4));
  nand2 gate580(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate581(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate582(.a(G657), .O(gate283inter7));
  inv1  gate583(.a(G809), .O(gate283inter8));
  nand2 gate584(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate585(.a(s_5), .b(gate283inter3), .O(gate283inter10));
  nor2  gate586(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate587(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate588(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate701(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate702(.a(gate284inter0), .b(s_22), .O(gate284inter1));
  and2  gate703(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate704(.a(s_22), .O(gate284inter3));
  inv1  gate705(.a(s_23), .O(gate284inter4));
  nand2 gate706(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate707(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate708(.a(G785), .O(gate284inter7));
  inv1  gate709(.a(G809), .O(gate284inter8));
  nand2 gate710(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate711(.a(s_23), .b(gate284inter3), .O(gate284inter10));
  nor2  gate712(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate713(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate714(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1415(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1416(.a(gate289inter0), .b(s_124), .O(gate289inter1));
  and2  gate1417(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1418(.a(s_124), .O(gate289inter3));
  inv1  gate1419(.a(s_125), .O(gate289inter4));
  nand2 gate1420(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1421(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1422(.a(G818), .O(gate289inter7));
  inv1  gate1423(.a(G819), .O(gate289inter8));
  nand2 gate1424(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1425(.a(s_125), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1426(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1427(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1428(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1849(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1850(.a(gate291inter0), .b(s_186), .O(gate291inter1));
  and2  gate1851(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1852(.a(s_186), .O(gate291inter3));
  inv1  gate1853(.a(s_187), .O(gate291inter4));
  nand2 gate1854(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1855(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1856(.a(G822), .O(gate291inter7));
  inv1  gate1857(.a(G823), .O(gate291inter8));
  nand2 gate1858(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1859(.a(s_187), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1860(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1861(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1862(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate953(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate954(.a(gate292inter0), .b(s_58), .O(gate292inter1));
  and2  gate955(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate956(.a(s_58), .O(gate292inter3));
  inv1  gate957(.a(s_59), .O(gate292inter4));
  nand2 gate958(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate959(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate960(.a(G824), .O(gate292inter7));
  inv1  gate961(.a(G825), .O(gate292inter8));
  nand2 gate962(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate963(.a(s_59), .b(gate292inter3), .O(gate292inter10));
  nor2  gate964(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate965(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate966(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1527(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1528(.a(gate293inter0), .b(s_140), .O(gate293inter1));
  and2  gate1529(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1530(.a(s_140), .O(gate293inter3));
  inv1  gate1531(.a(s_141), .O(gate293inter4));
  nand2 gate1532(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1533(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1534(.a(G828), .O(gate293inter7));
  inv1  gate1535(.a(G829), .O(gate293inter8));
  nand2 gate1536(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1537(.a(s_141), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1538(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1539(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1540(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate3067(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate3068(.a(gate294inter0), .b(s_360), .O(gate294inter1));
  and2  gate3069(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate3070(.a(s_360), .O(gate294inter3));
  inv1  gate3071(.a(s_361), .O(gate294inter4));
  nand2 gate3072(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate3073(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate3074(.a(G832), .O(gate294inter7));
  inv1  gate3075(.a(G833), .O(gate294inter8));
  nand2 gate3076(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate3077(.a(s_361), .b(gate294inter3), .O(gate294inter10));
  nor2  gate3078(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate3079(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate3080(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1639(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1640(.a(gate296inter0), .b(s_156), .O(gate296inter1));
  and2  gate1641(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1642(.a(s_156), .O(gate296inter3));
  inv1  gate1643(.a(s_157), .O(gate296inter4));
  nand2 gate1644(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1645(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1646(.a(G826), .O(gate296inter7));
  inv1  gate1647(.a(G827), .O(gate296inter8));
  nand2 gate1648(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1649(.a(s_157), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1650(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1651(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1652(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2031(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2032(.a(gate387inter0), .b(s_212), .O(gate387inter1));
  and2  gate2033(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2034(.a(s_212), .O(gate387inter3));
  inv1  gate2035(.a(s_213), .O(gate387inter4));
  nand2 gate2036(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2037(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2038(.a(G1), .O(gate387inter7));
  inv1  gate2039(.a(G1036), .O(gate387inter8));
  nand2 gate2040(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2041(.a(s_213), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2042(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2043(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2044(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1037(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1038(.a(gate390inter0), .b(s_70), .O(gate390inter1));
  and2  gate1039(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1040(.a(s_70), .O(gate390inter3));
  inv1  gate1041(.a(s_71), .O(gate390inter4));
  nand2 gate1042(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1043(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1044(.a(G4), .O(gate390inter7));
  inv1  gate1045(.a(G1045), .O(gate390inter8));
  nand2 gate1046(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1047(.a(s_71), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1048(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1049(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1050(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1205(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1206(.a(gate396inter0), .b(s_94), .O(gate396inter1));
  and2  gate1207(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1208(.a(s_94), .O(gate396inter3));
  inv1  gate1209(.a(s_95), .O(gate396inter4));
  nand2 gate1210(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1211(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1212(.a(G10), .O(gate396inter7));
  inv1  gate1213(.a(G1063), .O(gate396inter8));
  nand2 gate1214(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1215(.a(s_95), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1216(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1217(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1218(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1961(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1962(.a(gate397inter0), .b(s_202), .O(gate397inter1));
  and2  gate1963(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1964(.a(s_202), .O(gate397inter3));
  inv1  gate1965(.a(s_203), .O(gate397inter4));
  nand2 gate1966(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1967(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1968(.a(G11), .O(gate397inter7));
  inv1  gate1969(.a(G1066), .O(gate397inter8));
  nand2 gate1970(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1971(.a(s_203), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1972(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1973(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1974(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate2969(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2970(.a(gate399inter0), .b(s_346), .O(gate399inter1));
  and2  gate2971(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2972(.a(s_346), .O(gate399inter3));
  inv1  gate2973(.a(s_347), .O(gate399inter4));
  nand2 gate2974(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2975(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2976(.a(G13), .O(gate399inter7));
  inv1  gate2977(.a(G1072), .O(gate399inter8));
  nand2 gate2978(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2979(.a(s_347), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2980(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2981(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2982(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate743(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate744(.a(gate401inter0), .b(s_28), .O(gate401inter1));
  and2  gate745(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate746(.a(s_28), .O(gate401inter3));
  inv1  gate747(.a(s_29), .O(gate401inter4));
  nand2 gate748(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate749(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate750(.a(G15), .O(gate401inter7));
  inv1  gate751(.a(G1078), .O(gate401inter8));
  nand2 gate752(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate753(.a(s_29), .b(gate401inter3), .O(gate401inter10));
  nor2  gate754(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate755(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate756(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate2059(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2060(.a(gate405inter0), .b(s_216), .O(gate405inter1));
  and2  gate2061(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2062(.a(s_216), .O(gate405inter3));
  inv1  gate2063(.a(s_217), .O(gate405inter4));
  nand2 gate2064(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2065(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2066(.a(G19), .O(gate405inter7));
  inv1  gate2067(.a(G1090), .O(gate405inter8));
  nand2 gate2068(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2069(.a(s_217), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2070(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2071(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2072(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2339(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2340(.a(gate406inter0), .b(s_256), .O(gate406inter1));
  and2  gate2341(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2342(.a(s_256), .O(gate406inter3));
  inv1  gate2343(.a(s_257), .O(gate406inter4));
  nand2 gate2344(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2345(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2346(.a(G20), .O(gate406inter7));
  inv1  gate2347(.a(G1093), .O(gate406inter8));
  nand2 gate2348(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2349(.a(s_257), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2350(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2351(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2352(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate3249(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate3250(.a(gate407inter0), .b(s_386), .O(gate407inter1));
  and2  gate3251(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate3252(.a(s_386), .O(gate407inter3));
  inv1  gate3253(.a(s_387), .O(gate407inter4));
  nand2 gate3254(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate3255(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate3256(.a(G21), .O(gate407inter7));
  inv1  gate3257(.a(G1096), .O(gate407inter8));
  nand2 gate3258(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate3259(.a(s_387), .b(gate407inter3), .O(gate407inter10));
  nor2  gate3260(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate3261(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate3262(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate2913(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2914(.a(gate408inter0), .b(s_338), .O(gate408inter1));
  and2  gate2915(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2916(.a(s_338), .O(gate408inter3));
  inv1  gate2917(.a(s_339), .O(gate408inter4));
  nand2 gate2918(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2919(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2920(.a(G22), .O(gate408inter7));
  inv1  gate2921(.a(G1099), .O(gate408inter8));
  nand2 gate2922(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2923(.a(s_339), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2924(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2925(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2926(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate3123(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate3124(.a(gate413inter0), .b(s_368), .O(gate413inter1));
  and2  gate3125(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate3126(.a(s_368), .O(gate413inter3));
  inv1  gate3127(.a(s_369), .O(gate413inter4));
  nand2 gate3128(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate3129(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate3130(.a(G27), .O(gate413inter7));
  inv1  gate3131(.a(G1114), .O(gate413inter8));
  nand2 gate3132(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate3133(.a(s_369), .b(gate413inter3), .O(gate413inter10));
  nor2  gate3134(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate3135(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate3136(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2843(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2844(.a(gate414inter0), .b(s_328), .O(gate414inter1));
  and2  gate2845(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2846(.a(s_328), .O(gate414inter3));
  inv1  gate2847(.a(s_329), .O(gate414inter4));
  nand2 gate2848(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2849(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2850(.a(G28), .O(gate414inter7));
  inv1  gate2851(.a(G1117), .O(gate414inter8));
  nand2 gate2852(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2853(.a(s_329), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2854(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2855(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2856(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1107(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1108(.a(gate415inter0), .b(s_80), .O(gate415inter1));
  and2  gate1109(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1110(.a(s_80), .O(gate415inter3));
  inv1  gate1111(.a(s_81), .O(gate415inter4));
  nand2 gate1112(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1113(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1114(.a(G29), .O(gate415inter7));
  inv1  gate1115(.a(G1120), .O(gate415inter8));
  nand2 gate1116(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1117(.a(s_81), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1118(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1119(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1120(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate2493(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2494(.a(gate416inter0), .b(s_278), .O(gate416inter1));
  and2  gate2495(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2496(.a(s_278), .O(gate416inter3));
  inv1  gate2497(.a(s_279), .O(gate416inter4));
  nand2 gate2498(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2499(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2500(.a(G30), .O(gate416inter7));
  inv1  gate2501(.a(G1123), .O(gate416inter8));
  nand2 gate2502(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2503(.a(s_279), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2504(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2505(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2506(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2227(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2228(.a(gate420inter0), .b(s_240), .O(gate420inter1));
  and2  gate2229(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2230(.a(s_240), .O(gate420inter3));
  inv1  gate2231(.a(s_241), .O(gate420inter4));
  nand2 gate2232(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2233(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2234(.a(G1036), .O(gate420inter7));
  inv1  gate2235(.a(G1132), .O(gate420inter8));
  nand2 gate2236(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2237(.a(s_241), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2238(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2239(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2240(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate645(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate646(.a(gate423inter0), .b(s_14), .O(gate423inter1));
  and2  gate647(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate648(.a(s_14), .O(gate423inter3));
  inv1  gate649(.a(s_15), .O(gate423inter4));
  nand2 gate650(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate651(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate652(.a(G3), .O(gate423inter7));
  inv1  gate653(.a(G1138), .O(gate423inter8));
  nand2 gate654(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate655(.a(s_15), .b(gate423inter3), .O(gate423inter10));
  nor2  gate656(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate657(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate658(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate799(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate800(.a(gate424inter0), .b(s_36), .O(gate424inter1));
  and2  gate801(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate802(.a(s_36), .O(gate424inter3));
  inv1  gate803(.a(s_37), .O(gate424inter4));
  nand2 gate804(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate805(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate806(.a(G1042), .O(gate424inter7));
  inv1  gate807(.a(G1138), .O(gate424inter8));
  nand2 gate808(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate809(.a(s_37), .b(gate424inter3), .O(gate424inter10));
  nor2  gate810(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate811(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate812(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate3319(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate3320(.a(gate425inter0), .b(s_396), .O(gate425inter1));
  and2  gate3321(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate3322(.a(s_396), .O(gate425inter3));
  inv1  gate3323(.a(s_397), .O(gate425inter4));
  nand2 gate3324(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate3325(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate3326(.a(G4), .O(gate425inter7));
  inv1  gate3327(.a(G1141), .O(gate425inter8));
  nand2 gate3328(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate3329(.a(s_397), .b(gate425inter3), .O(gate425inter10));
  nor2  gate3330(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate3331(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate3332(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2731(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2732(.a(gate426inter0), .b(s_312), .O(gate426inter1));
  and2  gate2733(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2734(.a(s_312), .O(gate426inter3));
  inv1  gate2735(.a(s_313), .O(gate426inter4));
  nand2 gate2736(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2737(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2738(.a(G1045), .O(gate426inter7));
  inv1  gate2739(.a(G1141), .O(gate426inter8));
  nand2 gate2740(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2741(.a(s_313), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2742(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2743(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2744(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1751(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1752(.a(gate429inter0), .b(s_172), .O(gate429inter1));
  and2  gate1753(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1754(.a(s_172), .O(gate429inter3));
  inv1  gate1755(.a(s_173), .O(gate429inter4));
  nand2 gate1756(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1757(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1758(.a(G6), .O(gate429inter7));
  inv1  gate1759(.a(G1147), .O(gate429inter8));
  nand2 gate1760(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1761(.a(s_173), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1762(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1763(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1764(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2283(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2284(.a(gate431inter0), .b(s_248), .O(gate431inter1));
  and2  gate2285(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2286(.a(s_248), .O(gate431inter3));
  inv1  gate2287(.a(s_249), .O(gate431inter4));
  nand2 gate2288(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2289(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2290(.a(G7), .O(gate431inter7));
  inv1  gate2291(.a(G1150), .O(gate431inter8));
  nand2 gate2292(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2293(.a(s_249), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2294(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2295(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2296(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1023(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1024(.a(gate432inter0), .b(s_68), .O(gate432inter1));
  and2  gate1025(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1026(.a(s_68), .O(gate432inter3));
  inv1  gate1027(.a(s_69), .O(gate432inter4));
  nand2 gate1028(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1029(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1030(.a(G1054), .O(gate432inter7));
  inv1  gate1031(.a(G1150), .O(gate432inter8));
  nand2 gate1032(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1033(.a(s_69), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1034(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1035(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1036(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate673(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate674(.a(gate434inter0), .b(s_18), .O(gate434inter1));
  and2  gate675(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate676(.a(s_18), .O(gate434inter3));
  inv1  gate677(.a(s_19), .O(gate434inter4));
  nand2 gate678(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate679(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate680(.a(G1057), .O(gate434inter7));
  inv1  gate681(.a(G1153), .O(gate434inter8));
  nand2 gate682(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate683(.a(s_19), .b(gate434inter3), .O(gate434inter10));
  nor2  gate684(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate685(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate686(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2745(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2746(.a(gate435inter0), .b(s_314), .O(gate435inter1));
  and2  gate2747(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2748(.a(s_314), .O(gate435inter3));
  inv1  gate2749(.a(s_315), .O(gate435inter4));
  nand2 gate2750(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2751(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2752(.a(G9), .O(gate435inter7));
  inv1  gate2753(.a(G1156), .O(gate435inter8));
  nand2 gate2754(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2755(.a(s_315), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2756(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2757(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2758(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate827(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate828(.a(gate436inter0), .b(s_40), .O(gate436inter1));
  and2  gate829(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate830(.a(s_40), .O(gate436inter3));
  inv1  gate831(.a(s_41), .O(gate436inter4));
  nand2 gate832(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate833(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate834(.a(G1060), .O(gate436inter7));
  inv1  gate835(.a(G1156), .O(gate436inter8));
  nand2 gate836(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate837(.a(s_41), .b(gate436inter3), .O(gate436inter10));
  nor2  gate838(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate839(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate840(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2353(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2354(.a(gate439inter0), .b(s_258), .O(gate439inter1));
  and2  gate2355(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2356(.a(s_258), .O(gate439inter3));
  inv1  gate2357(.a(s_259), .O(gate439inter4));
  nand2 gate2358(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2359(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2360(.a(G11), .O(gate439inter7));
  inv1  gate2361(.a(G1162), .O(gate439inter8));
  nand2 gate2362(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2363(.a(s_259), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2364(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2365(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2366(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2325(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2326(.a(gate441inter0), .b(s_254), .O(gate441inter1));
  and2  gate2327(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2328(.a(s_254), .O(gate441inter3));
  inv1  gate2329(.a(s_255), .O(gate441inter4));
  nand2 gate2330(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2331(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2332(.a(G12), .O(gate441inter7));
  inv1  gate2333(.a(G1165), .O(gate441inter8));
  nand2 gate2334(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2335(.a(s_255), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2336(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2337(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2338(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2801(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2802(.a(gate444inter0), .b(s_322), .O(gate444inter1));
  and2  gate2803(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2804(.a(s_322), .O(gate444inter3));
  inv1  gate2805(.a(s_323), .O(gate444inter4));
  nand2 gate2806(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2807(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2808(.a(G1072), .O(gate444inter7));
  inv1  gate2809(.a(G1168), .O(gate444inter8));
  nand2 gate2810(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2811(.a(s_323), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2812(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2813(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2814(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2871(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2872(.a(gate446inter0), .b(s_332), .O(gate446inter1));
  and2  gate2873(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2874(.a(s_332), .O(gate446inter3));
  inv1  gate2875(.a(s_333), .O(gate446inter4));
  nand2 gate2876(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2877(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2878(.a(G1075), .O(gate446inter7));
  inv1  gate2879(.a(G1171), .O(gate446inter8));
  nand2 gate2880(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2881(.a(s_333), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2882(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2883(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2884(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2591(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2592(.a(gate447inter0), .b(s_292), .O(gate447inter1));
  and2  gate2593(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2594(.a(s_292), .O(gate447inter3));
  inv1  gate2595(.a(s_293), .O(gate447inter4));
  nand2 gate2596(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2597(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2598(.a(G15), .O(gate447inter7));
  inv1  gate2599(.a(G1174), .O(gate447inter8));
  nand2 gate2600(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2601(.a(s_293), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2602(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2603(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2604(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate3193(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate3194(.a(gate448inter0), .b(s_378), .O(gate448inter1));
  and2  gate3195(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate3196(.a(s_378), .O(gate448inter3));
  inv1  gate3197(.a(s_379), .O(gate448inter4));
  nand2 gate3198(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate3199(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate3200(.a(G1078), .O(gate448inter7));
  inv1  gate3201(.a(G1174), .O(gate448inter8));
  nand2 gate3202(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate3203(.a(s_379), .b(gate448inter3), .O(gate448inter10));
  nor2  gate3204(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate3205(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate3206(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate3151(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate3152(.a(gate450inter0), .b(s_372), .O(gate450inter1));
  and2  gate3153(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate3154(.a(s_372), .O(gate450inter3));
  inv1  gate3155(.a(s_373), .O(gate450inter4));
  nand2 gate3156(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate3157(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate3158(.a(G1081), .O(gate450inter7));
  inv1  gate3159(.a(G1177), .O(gate450inter8));
  nand2 gate3160(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate3161(.a(s_373), .b(gate450inter3), .O(gate450inter10));
  nor2  gate3162(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate3163(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate3164(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2703(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2704(.a(gate452inter0), .b(s_308), .O(gate452inter1));
  and2  gate2705(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2706(.a(s_308), .O(gate452inter3));
  inv1  gate2707(.a(s_309), .O(gate452inter4));
  nand2 gate2708(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2709(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2710(.a(G1084), .O(gate452inter7));
  inv1  gate2711(.a(G1180), .O(gate452inter8));
  nand2 gate2712(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2713(.a(s_309), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2714(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2715(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2716(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate855(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate856(.a(gate456inter0), .b(s_44), .O(gate456inter1));
  and2  gate857(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate858(.a(s_44), .O(gate456inter3));
  inv1  gate859(.a(s_45), .O(gate456inter4));
  nand2 gate860(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate861(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate862(.a(G1090), .O(gate456inter7));
  inv1  gate863(.a(G1186), .O(gate456inter8));
  nand2 gate864(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate865(.a(s_45), .b(gate456inter3), .O(gate456inter10));
  nor2  gate866(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate867(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate868(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate897(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate898(.a(gate459inter0), .b(s_50), .O(gate459inter1));
  and2  gate899(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate900(.a(s_50), .O(gate459inter3));
  inv1  gate901(.a(s_51), .O(gate459inter4));
  nand2 gate902(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate903(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate904(.a(G21), .O(gate459inter7));
  inv1  gate905(.a(G1192), .O(gate459inter8));
  nand2 gate906(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate907(.a(s_51), .b(gate459inter3), .O(gate459inter10));
  nor2  gate908(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate909(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate910(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2451(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2452(.a(gate464inter0), .b(s_272), .O(gate464inter1));
  and2  gate2453(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2454(.a(s_272), .O(gate464inter3));
  inv1  gate2455(.a(s_273), .O(gate464inter4));
  nand2 gate2456(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2457(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2458(.a(G1102), .O(gate464inter7));
  inv1  gate2459(.a(G1198), .O(gate464inter8));
  nand2 gate2460(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2461(.a(s_273), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2462(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2463(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2464(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2269(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2270(.a(gate466inter0), .b(s_246), .O(gate466inter1));
  and2  gate2271(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2272(.a(s_246), .O(gate466inter3));
  inv1  gate2273(.a(s_247), .O(gate466inter4));
  nand2 gate2274(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2275(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2276(.a(G1105), .O(gate466inter7));
  inv1  gate2277(.a(G1201), .O(gate466inter8));
  nand2 gate2278(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2279(.a(s_247), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2280(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2281(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2282(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate603(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate604(.a(gate468inter0), .b(s_8), .O(gate468inter1));
  and2  gate605(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate606(.a(s_8), .O(gate468inter3));
  inv1  gate607(.a(s_9), .O(gate468inter4));
  nand2 gate608(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate609(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate610(.a(G1108), .O(gate468inter7));
  inv1  gate611(.a(G1204), .O(gate468inter8));
  nand2 gate612(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate613(.a(s_9), .b(gate468inter3), .O(gate468inter10));
  nor2  gate614(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate615(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate616(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate1149(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1150(.a(gate469inter0), .b(s_86), .O(gate469inter1));
  and2  gate1151(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1152(.a(s_86), .O(gate469inter3));
  inv1  gate1153(.a(s_87), .O(gate469inter4));
  nand2 gate1154(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1155(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1156(.a(G26), .O(gate469inter7));
  inv1  gate1157(.a(G1207), .O(gate469inter8));
  nand2 gate1158(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1159(.a(s_87), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1160(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1161(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1162(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2157(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2158(.a(gate470inter0), .b(s_230), .O(gate470inter1));
  and2  gate2159(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2160(.a(s_230), .O(gate470inter3));
  inv1  gate2161(.a(s_231), .O(gate470inter4));
  nand2 gate2162(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2163(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2164(.a(G1111), .O(gate470inter7));
  inv1  gate2165(.a(G1207), .O(gate470inter8));
  nand2 gate2166(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2167(.a(s_231), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2168(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2169(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2170(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1443(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1444(.a(gate472inter0), .b(s_128), .O(gate472inter1));
  and2  gate1445(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1446(.a(s_128), .O(gate472inter3));
  inv1  gate1447(.a(s_129), .O(gate472inter4));
  nand2 gate1448(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1449(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1450(.a(G1114), .O(gate472inter7));
  inv1  gate1451(.a(G1210), .O(gate472inter8));
  nand2 gate1452(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1453(.a(s_129), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1454(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1455(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1456(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1233(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1234(.a(gate474inter0), .b(s_98), .O(gate474inter1));
  and2  gate1235(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1236(.a(s_98), .O(gate474inter3));
  inv1  gate1237(.a(s_99), .O(gate474inter4));
  nand2 gate1238(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1239(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1240(.a(G1117), .O(gate474inter7));
  inv1  gate1241(.a(G1213), .O(gate474inter8));
  nand2 gate1242(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1243(.a(s_99), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1244(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1245(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1246(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2549(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2550(.a(gate477inter0), .b(s_286), .O(gate477inter1));
  and2  gate2551(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2552(.a(s_286), .O(gate477inter3));
  inv1  gate2553(.a(s_287), .O(gate477inter4));
  nand2 gate2554(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2555(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2556(.a(G30), .O(gate477inter7));
  inv1  gate2557(.a(G1219), .O(gate477inter8));
  nand2 gate2558(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2559(.a(s_287), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2560(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2561(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2562(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2213(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2214(.a(gate478inter0), .b(s_238), .O(gate478inter1));
  and2  gate2215(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2216(.a(s_238), .O(gate478inter3));
  inv1  gate2217(.a(s_239), .O(gate478inter4));
  nand2 gate2218(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2219(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2220(.a(G1123), .O(gate478inter7));
  inv1  gate2221(.a(G1219), .O(gate478inter8));
  nand2 gate2222(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2223(.a(s_239), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2224(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2225(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2226(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2395(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2396(.a(gate479inter0), .b(s_264), .O(gate479inter1));
  and2  gate2397(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2398(.a(s_264), .O(gate479inter3));
  inv1  gate2399(.a(s_265), .O(gate479inter4));
  nand2 gate2400(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2401(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2402(.a(G31), .O(gate479inter7));
  inv1  gate2403(.a(G1222), .O(gate479inter8));
  nand2 gate2404(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2405(.a(s_265), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2406(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2407(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2408(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1905(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1906(.a(gate482inter0), .b(s_194), .O(gate482inter1));
  and2  gate1907(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1908(.a(s_194), .O(gate482inter3));
  inv1  gate1909(.a(s_195), .O(gate482inter4));
  nand2 gate1910(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1911(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1912(.a(G1129), .O(gate482inter7));
  inv1  gate1913(.a(G1225), .O(gate482inter8));
  nand2 gate1914(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1915(.a(s_195), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1916(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1917(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1918(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1555(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1556(.a(gate484inter0), .b(s_144), .O(gate484inter1));
  and2  gate1557(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1558(.a(s_144), .O(gate484inter3));
  inv1  gate1559(.a(s_145), .O(gate484inter4));
  nand2 gate1560(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1561(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1562(.a(G1230), .O(gate484inter7));
  inv1  gate1563(.a(G1231), .O(gate484inter8));
  nand2 gate1564(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1565(.a(s_145), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1566(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1567(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1568(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2185(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2186(.a(gate485inter0), .b(s_234), .O(gate485inter1));
  and2  gate2187(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2188(.a(s_234), .O(gate485inter3));
  inv1  gate2189(.a(s_235), .O(gate485inter4));
  nand2 gate2190(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2191(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2192(.a(G1232), .O(gate485inter7));
  inv1  gate2193(.a(G1233), .O(gate485inter8));
  nand2 gate2194(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2195(.a(s_235), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2196(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2197(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2198(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate2885(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2886(.a(gate486inter0), .b(s_334), .O(gate486inter1));
  and2  gate2887(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2888(.a(s_334), .O(gate486inter3));
  inv1  gate2889(.a(s_335), .O(gate486inter4));
  nand2 gate2890(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2891(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2892(.a(G1234), .O(gate486inter7));
  inv1  gate2893(.a(G1235), .O(gate486inter8));
  nand2 gate2894(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2895(.a(s_335), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2896(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2897(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2898(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1625(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1626(.a(gate488inter0), .b(s_154), .O(gate488inter1));
  and2  gate1627(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1628(.a(s_154), .O(gate488inter3));
  inv1  gate1629(.a(s_155), .O(gate488inter4));
  nand2 gate1630(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1631(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1632(.a(G1238), .O(gate488inter7));
  inv1  gate1633(.a(G1239), .O(gate488inter8));
  nand2 gate1634(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1635(.a(s_155), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1636(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1637(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1638(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate3291(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate3292(.a(gate490inter0), .b(s_392), .O(gate490inter1));
  and2  gate3293(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate3294(.a(s_392), .O(gate490inter3));
  inv1  gate3295(.a(s_393), .O(gate490inter4));
  nand2 gate3296(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate3297(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate3298(.a(G1242), .O(gate490inter7));
  inv1  gate3299(.a(G1243), .O(gate490inter8));
  nand2 gate3300(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate3301(.a(s_393), .b(gate490inter3), .O(gate490inter10));
  nor2  gate3302(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate3303(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate3304(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1611(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1612(.a(gate491inter0), .b(s_152), .O(gate491inter1));
  and2  gate1613(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1614(.a(s_152), .O(gate491inter3));
  inv1  gate1615(.a(s_153), .O(gate491inter4));
  nand2 gate1616(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1617(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1618(.a(G1244), .O(gate491inter7));
  inv1  gate1619(.a(G1245), .O(gate491inter8));
  nand2 gate1620(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1621(.a(s_153), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1622(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1623(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1624(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1065(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1066(.a(gate492inter0), .b(s_74), .O(gate492inter1));
  and2  gate1067(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1068(.a(s_74), .O(gate492inter3));
  inv1  gate1069(.a(s_75), .O(gate492inter4));
  nand2 gate1070(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1071(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1072(.a(G1246), .O(gate492inter7));
  inv1  gate1073(.a(G1247), .O(gate492inter8));
  nand2 gate1074(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1075(.a(s_75), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1076(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1077(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1078(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1079(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1080(.a(gate494inter0), .b(s_76), .O(gate494inter1));
  and2  gate1081(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1082(.a(s_76), .O(gate494inter3));
  inv1  gate1083(.a(s_77), .O(gate494inter4));
  nand2 gate1084(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1085(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1086(.a(G1250), .O(gate494inter7));
  inv1  gate1087(.a(G1251), .O(gate494inter8));
  nand2 gate1088(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1089(.a(s_77), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1090(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1091(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1092(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate659(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate660(.a(gate495inter0), .b(s_16), .O(gate495inter1));
  and2  gate661(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate662(.a(s_16), .O(gate495inter3));
  inv1  gate663(.a(s_17), .O(gate495inter4));
  nand2 gate664(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate665(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate666(.a(G1252), .O(gate495inter7));
  inv1  gate667(.a(G1253), .O(gate495inter8));
  nand2 gate668(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate669(.a(s_17), .b(gate495inter3), .O(gate495inter10));
  nor2  gate670(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate671(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate672(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate547(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate548(.a(gate498inter0), .b(s_0), .O(gate498inter1));
  and2  gate549(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate550(.a(s_0), .O(gate498inter3));
  inv1  gate551(.a(s_1), .O(gate498inter4));
  nand2 gate552(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate553(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate554(.a(G1258), .O(gate498inter7));
  inv1  gate555(.a(G1259), .O(gate498inter8));
  nand2 gate556(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate557(.a(s_1), .b(gate498inter3), .O(gate498inter10));
  nor2  gate558(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate559(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate560(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1793(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1794(.a(gate501inter0), .b(s_178), .O(gate501inter1));
  and2  gate1795(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1796(.a(s_178), .O(gate501inter3));
  inv1  gate1797(.a(s_179), .O(gate501inter4));
  nand2 gate1798(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1799(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1800(.a(G1264), .O(gate501inter7));
  inv1  gate1801(.a(G1265), .O(gate501inter8));
  nand2 gate1802(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1803(.a(s_179), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1804(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1805(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1806(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2507(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2508(.a(gate502inter0), .b(s_280), .O(gate502inter1));
  and2  gate2509(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2510(.a(s_280), .O(gate502inter3));
  inv1  gate2511(.a(s_281), .O(gate502inter4));
  nand2 gate2512(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2513(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2514(.a(G1266), .O(gate502inter7));
  inv1  gate2515(.a(G1267), .O(gate502inter8));
  nand2 gate2516(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2517(.a(s_281), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2518(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2519(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2520(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2521(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2522(.a(gate503inter0), .b(s_282), .O(gate503inter1));
  and2  gate2523(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2524(.a(s_282), .O(gate503inter3));
  inv1  gate2525(.a(s_283), .O(gate503inter4));
  nand2 gate2526(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2527(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2528(.a(G1268), .O(gate503inter7));
  inv1  gate2529(.a(G1269), .O(gate503inter8));
  nand2 gate2530(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2531(.a(s_283), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2532(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2533(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2534(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2759(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2760(.a(gate505inter0), .b(s_316), .O(gate505inter1));
  and2  gate2761(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2762(.a(s_316), .O(gate505inter3));
  inv1  gate2763(.a(s_317), .O(gate505inter4));
  nand2 gate2764(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2765(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2766(.a(G1272), .O(gate505inter7));
  inv1  gate2767(.a(G1273), .O(gate505inter8));
  nand2 gate2768(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2769(.a(s_317), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2770(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2771(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2772(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate3207(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate3208(.a(gate506inter0), .b(s_380), .O(gate506inter1));
  and2  gate3209(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate3210(.a(s_380), .O(gate506inter3));
  inv1  gate3211(.a(s_381), .O(gate506inter4));
  nand2 gate3212(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate3213(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate3214(.a(G1274), .O(gate506inter7));
  inv1  gate3215(.a(G1275), .O(gate506inter8));
  nand2 gate3216(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate3217(.a(s_381), .b(gate506inter3), .O(gate506inter10));
  nor2  gate3218(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate3219(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate3220(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1499(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1500(.a(gate507inter0), .b(s_136), .O(gate507inter1));
  and2  gate1501(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1502(.a(s_136), .O(gate507inter3));
  inv1  gate1503(.a(s_137), .O(gate507inter4));
  nand2 gate1504(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1505(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1506(.a(G1276), .O(gate507inter7));
  inv1  gate1507(.a(G1277), .O(gate507inter8));
  nand2 gate1508(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1509(.a(s_137), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1510(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1511(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1512(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1667(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1668(.a(gate508inter0), .b(s_160), .O(gate508inter1));
  and2  gate1669(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1670(.a(s_160), .O(gate508inter3));
  inv1  gate1671(.a(s_161), .O(gate508inter4));
  nand2 gate1672(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1673(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1674(.a(G1278), .O(gate508inter7));
  inv1  gate1675(.a(G1279), .O(gate508inter8));
  nand2 gate1676(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1677(.a(s_161), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1678(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1679(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1680(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1051(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1052(.a(gate509inter0), .b(s_72), .O(gate509inter1));
  and2  gate1053(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1054(.a(s_72), .O(gate509inter3));
  inv1  gate1055(.a(s_73), .O(gate509inter4));
  nand2 gate1056(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1057(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1058(.a(G1280), .O(gate509inter7));
  inv1  gate1059(.a(G1281), .O(gate509inter8));
  nand2 gate1060(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1061(.a(s_73), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1062(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1063(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1064(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate771(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate772(.a(gate510inter0), .b(s_32), .O(gate510inter1));
  and2  gate773(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate774(.a(s_32), .O(gate510inter3));
  inv1  gate775(.a(s_33), .O(gate510inter4));
  nand2 gate776(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate777(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate778(.a(G1282), .O(gate510inter7));
  inv1  gate779(.a(G1283), .O(gate510inter8));
  nand2 gate780(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate781(.a(s_33), .b(gate510inter3), .O(gate510inter10));
  nor2  gate782(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate783(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate784(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate3277(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate3278(.a(gate514inter0), .b(s_390), .O(gate514inter1));
  and2  gate3279(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate3280(.a(s_390), .O(gate514inter3));
  inv1  gate3281(.a(s_391), .O(gate514inter4));
  nand2 gate3282(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate3283(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate3284(.a(G1290), .O(gate514inter7));
  inv1  gate3285(.a(G1291), .O(gate514inter8));
  nand2 gate3286(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate3287(.a(s_391), .b(gate514inter3), .O(gate514inter10));
  nor2  gate3288(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate3289(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate3290(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule