module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2101(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2102(.a(gate15inter0), .b(s_222), .O(gate15inter1));
  and2  gate2103(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2104(.a(s_222), .O(gate15inter3));
  inv1  gate2105(.a(s_223), .O(gate15inter4));
  nand2 gate2106(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2107(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2108(.a(G13), .O(gate15inter7));
  inv1  gate2109(.a(G14), .O(gate15inter8));
  nand2 gate2110(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2111(.a(s_223), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2112(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2113(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2114(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1121(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1122(.a(gate26inter0), .b(s_82), .O(gate26inter1));
  and2  gate1123(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1124(.a(s_82), .O(gate26inter3));
  inv1  gate1125(.a(s_83), .O(gate26inter4));
  nand2 gate1126(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1127(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1128(.a(G9), .O(gate26inter7));
  inv1  gate1129(.a(G13), .O(gate26inter8));
  nand2 gate1130(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1131(.a(s_83), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1132(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1133(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1134(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1387(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1388(.a(gate32inter0), .b(s_120), .O(gate32inter1));
  and2  gate1389(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1390(.a(s_120), .O(gate32inter3));
  inv1  gate1391(.a(s_121), .O(gate32inter4));
  nand2 gate1392(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1393(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1394(.a(G12), .O(gate32inter7));
  inv1  gate1395(.a(G16), .O(gate32inter8));
  nand2 gate1396(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1397(.a(s_121), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1398(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1399(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1400(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1989(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1990(.a(gate33inter0), .b(s_206), .O(gate33inter1));
  and2  gate1991(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1992(.a(s_206), .O(gate33inter3));
  inv1  gate1993(.a(s_207), .O(gate33inter4));
  nand2 gate1994(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1995(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1996(.a(G17), .O(gate33inter7));
  inv1  gate1997(.a(G21), .O(gate33inter8));
  nand2 gate1998(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1999(.a(s_207), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2000(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2001(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2002(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1793(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1794(.a(gate35inter0), .b(s_178), .O(gate35inter1));
  and2  gate1795(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1796(.a(s_178), .O(gate35inter3));
  inv1  gate1797(.a(s_179), .O(gate35inter4));
  nand2 gate1798(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1799(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1800(.a(G18), .O(gate35inter7));
  inv1  gate1801(.a(G22), .O(gate35inter8));
  nand2 gate1802(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1803(.a(s_179), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1804(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1805(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1806(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1009(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1010(.a(gate37inter0), .b(s_66), .O(gate37inter1));
  and2  gate1011(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1012(.a(s_66), .O(gate37inter3));
  inv1  gate1013(.a(s_67), .O(gate37inter4));
  nand2 gate1014(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1015(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1016(.a(G19), .O(gate37inter7));
  inv1  gate1017(.a(G23), .O(gate37inter8));
  nand2 gate1018(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1019(.a(s_67), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1020(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1021(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1022(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate925(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate926(.a(gate40inter0), .b(s_54), .O(gate40inter1));
  and2  gate927(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate928(.a(s_54), .O(gate40inter3));
  inv1  gate929(.a(s_55), .O(gate40inter4));
  nand2 gate930(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate931(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate932(.a(G28), .O(gate40inter7));
  inv1  gate933(.a(G32), .O(gate40inter8));
  nand2 gate934(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate935(.a(s_55), .b(gate40inter3), .O(gate40inter10));
  nor2  gate936(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate937(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate938(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate911(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate912(.a(gate46inter0), .b(s_52), .O(gate46inter1));
  and2  gate913(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate914(.a(s_52), .O(gate46inter3));
  inv1  gate915(.a(s_53), .O(gate46inter4));
  nand2 gate916(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate917(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate918(.a(G6), .O(gate46inter7));
  inv1  gate919(.a(G272), .O(gate46inter8));
  nand2 gate920(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate921(.a(s_53), .b(gate46inter3), .O(gate46inter10));
  nor2  gate922(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate923(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate924(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate743(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate744(.a(gate54inter0), .b(s_28), .O(gate54inter1));
  and2  gate745(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate746(.a(s_28), .O(gate54inter3));
  inv1  gate747(.a(s_29), .O(gate54inter4));
  nand2 gate748(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate749(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate750(.a(G14), .O(gate54inter7));
  inv1  gate751(.a(G284), .O(gate54inter8));
  nand2 gate752(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate753(.a(s_29), .b(gate54inter3), .O(gate54inter10));
  nor2  gate754(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate755(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate756(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate827(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate828(.a(gate57inter0), .b(s_40), .O(gate57inter1));
  and2  gate829(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate830(.a(s_40), .O(gate57inter3));
  inv1  gate831(.a(s_41), .O(gate57inter4));
  nand2 gate832(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate833(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate834(.a(G17), .O(gate57inter7));
  inv1  gate835(.a(G290), .O(gate57inter8));
  nand2 gate836(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate837(.a(s_41), .b(gate57inter3), .O(gate57inter10));
  nor2  gate838(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate839(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate840(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1247(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1248(.a(gate63inter0), .b(s_100), .O(gate63inter1));
  and2  gate1249(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1250(.a(s_100), .O(gate63inter3));
  inv1  gate1251(.a(s_101), .O(gate63inter4));
  nand2 gate1252(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1253(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1254(.a(G23), .O(gate63inter7));
  inv1  gate1255(.a(G299), .O(gate63inter8));
  nand2 gate1256(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1257(.a(s_101), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1258(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1259(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1260(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1751(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1752(.a(gate66inter0), .b(s_172), .O(gate66inter1));
  and2  gate1753(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1754(.a(s_172), .O(gate66inter3));
  inv1  gate1755(.a(s_173), .O(gate66inter4));
  nand2 gate1756(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1757(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1758(.a(G26), .O(gate66inter7));
  inv1  gate1759(.a(G302), .O(gate66inter8));
  nand2 gate1760(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1761(.a(s_173), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1762(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1763(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1764(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1373(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1374(.a(gate69inter0), .b(s_118), .O(gate69inter1));
  and2  gate1375(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1376(.a(s_118), .O(gate69inter3));
  inv1  gate1377(.a(s_119), .O(gate69inter4));
  nand2 gate1378(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1379(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1380(.a(G29), .O(gate69inter7));
  inv1  gate1381(.a(G308), .O(gate69inter8));
  nand2 gate1382(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1383(.a(s_119), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1384(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1385(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1386(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2073(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2074(.a(gate74inter0), .b(s_218), .O(gate74inter1));
  and2  gate2075(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2076(.a(s_218), .O(gate74inter3));
  inv1  gate2077(.a(s_219), .O(gate74inter4));
  nand2 gate2078(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2079(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2080(.a(G5), .O(gate74inter7));
  inv1  gate2081(.a(G314), .O(gate74inter8));
  nand2 gate2082(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2083(.a(s_219), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2084(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2085(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2086(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2059(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2060(.a(gate79inter0), .b(s_216), .O(gate79inter1));
  and2  gate2061(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2062(.a(s_216), .O(gate79inter3));
  inv1  gate2063(.a(s_217), .O(gate79inter4));
  nand2 gate2064(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2065(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2066(.a(G10), .O(gate79inter7));
  inv1  gate2067(.a(G323), .O(gate79inter8));
  nand2 gate2068(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2069(.a(s_217), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2070(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2071(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2072(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1821(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1822(.a(gate85inter0), .b(s_182), .O(gate85inter1));
  and2  gate1823(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1824(.a(s_182), .O(gate85inter3));
  inv1  gate1825(.a(s_183), .O(gate85inter4));
  nand2 gate1826(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1827(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1828(.a(G4), .O(gate85inter7));
  inv1  gate1829(.a(G332), .O(gate85inter8));
  nand2 gate1830(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1831(.a(s_183), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1832(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1833(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1834(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate771(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate772(.a(gate87inter0), .b(s_32), .O(gate87inter1));
  and2  gate773(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate774(.a(s_32), .O(gate87inter3));
  inv1  gate775(.a(s_33), .O(gate87inter4));
  nand2 gate776(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate777(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate778(.a(G12), .O(gate87inter7));
  inv1  gate779(.a(G335), .O(gate87inter8));
  nand2 gate780(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate781(.a(s_33), .b(gate87inter3), .O(gate87inter10));
  nor2  gate782(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate783(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate784(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate897(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate898(.a(gate91inter0), .b(s_50), .O(gate91inter1));
  and2  gate899(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate900(.a(s_50), .O(gate91inter3));
  inv1  gate901(.a(s_51), .O(gate91inter4));
  nand2 gate902(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate903(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate904(.a(G25), .O(gate91inter7));
  inv1  gate905(.a(G341), .O(gate91inter8));
  nand2 gate906(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate907(.a(s_51), .b(gate91inter3), .O(gate91inter10));
  nor2  gate908(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate909(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate910(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1023(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1024(.a(gate94inter0), .b(s_68), .O(gate94inter1));
  and2  gate1025(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1026(.a(s_68), .O(gate94inter3));
  inv1  gate1027(.a(s_69), .O(gate94inter4));
  nand2 gate1028(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1029(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1030(.a(G22), .O(gate94inter7));
  inv1  gate1031(.a(G344), .O(gate94inter8));
  nand2 gate1032(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1033(.a(s_69), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1034(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1035(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1036(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1093(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1094(.a(gate95inter0), .b(s_78), .O(gate95inter1));
  and2  gate1095(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1096(.a(s_78), .O(gate95inter3));
  inv1  gate1097(.a(s_79), .O(gate95inter4));
  nand2 gate1098(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1099(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1100(.a(G26), .O(gate95inter7));
  inv1  gate1101(.a(G347), .O(gate95inter8));
  nand2 gate1102(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1103(.a(s_79), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1104(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1105(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1106(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1233(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1234(.a(gate98inter0), .b(s_98), .O(gate98inter1));
  and2  gate1235(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1236(.a(s_98), .O(gate98inter3));
  inv1  gate1237(.a(s_99), .O(gate98inter4));
  nand2 gate1238(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1239(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1240(.a(G23), .O(gate98inter7));
  inv1  gate1241(.a(G350), .O(gate98inter8));
  nand2 gate1242(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1243(.a(s_99), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1244(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1245(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1246(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1555(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1556(.a(gate101inter0), .b(s_144), .O(gate101inter1));
  and2  gate1557(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1558(.a(s_144), .O(gate101inter3));
  inv1  gate1559(.a(s_145), .O(gate101inter4));
  nand2 gate1560(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1561(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1562(.a(G20), .O(gate101inter7));
  inv1  gate1563(.a(G356), .O(gate101inter8));
  nand2 gate1564(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1565(.a(s_145), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1566(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1567(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1568(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate841(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate842(.a(gate102inter0), .b(s_42), .O(gate102inter1));
  and2  gate843(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate844(.a(s_42), .O(gate102inter3));
  inv1  gate845(.a(s_43), .O(gate102inter4));
  nand2 gate846(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate847(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate848(.a(G24), .O(gate102inter7));
  inv1  gate849(.a(G356), .O(gate102inter8));
  nand2 gate850(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate851(.a(s_43), .b(gate102inter3), .O(gate102inter10));
  nor2  gate852(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate853(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate854(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2017(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2018(.a(gate105inter0), .b(s_210), .O(gate105inter1));
  and2  gate2019(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2020(.a(s_210), .O(gate105inter3));
  inv1  gate2021(.a(s_211), .O(gate105inter4));
  nand2 gate2022(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2023(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2024(.a(G362), .O(gate105inter7));
  inv1  gate2025(.a(G363), .O(gate105inter8));
  nand2 gate2026(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2027(.a(s_211), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2028(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2029(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2030(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1765(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1766(.a(gate106inter0), .b(s_174), .O(gate106inter1));
  and2  gate1767(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1768(.a(s_174), .O(gate106inter3));
  inv1  gate1769(.a(s_175), .O(gate106inter4));
  nand2 gate1770(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1771(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1772(.a(G364), .O(gate106inter7));
  inv1  gate1773(.a(G365), .O(gate106inter8));
  nand2 gate1774(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1775(.a(s_175), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1776(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1777(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1778(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1499(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1500(.a(gate108inter0), .b(s_136), .O(gate108inter1));
  and2  gate1501(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1502(.a(s_136), .O(gate108inter3));
  inv1  gate1503(.a(s_137), .O(gate108inter4));
  nand2 gate1504(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1505(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1506(.a(G368), .O(gate108inter7));
  inv1  gate1507(.a(G369), .O(gate108inter8));
  nand2 gate1508(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1509(.a(s_137), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1510(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1511(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1512(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1835(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1836(.a(gate109inter0), .b(s_184), .O(gate109inter1));
  and2  gate1837(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1838(.a(s_184), .O(gate109inter3));
  inv1  gate1839(.a(s_185), .O(gate109inter4));
  nand2 gate1840(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1841(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1842(.a(G370), .O(gate109inter7));
  inv1  gate1843(.a(G371), .O(gate109inter8));
  nand2 gate1844(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1845(.a(s_185), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1846(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1847(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1848(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1359(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1360(.a(gate123inter0), .b(s_116), .O(gate123inter1));
  and2  gate1361(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1362(.a(s_116), .O(gate123inter3));
  inv1  gate1363(.a(s_117), .O(gate123inter4));
  nand2 gate1364(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1365(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1366(.a(G398), .O(gate123inter7));
  inv1  gate1367(.a(G399), .O(gate123inter8));
  nand2 gate1368(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1369(.a(s_117), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1370(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1371(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1372(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1597(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1598(.a(gate124inter0), .b(s_150), .O(gate124inter1));
  and2  gate1599(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1600(.a(s_150), .O(gate124inter3));
  inv1  gate1601(.a(s_151), .O(gate124inter4));
  nand2 gate1602(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1603(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1604(.a(G400), .O(gate124inter7));
  inv1  gate1605(.a(G401), .O(gate124inter8));
  nand2 gate1606(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1607(.a(s_151), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1608(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1609(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1610(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1933(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1934(.a(gate129inter0), .b(s_198), .O(gate129inter1));
  and2  gate1935(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1936(.a(s_198), .O(gate129inter3));
  inv1  gate1937(.a(s_199), .O(gate129inter4));
  nand2 gate1938(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1939(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1940(.a(G410), .O(gate129inter7));
  inv1  gate1941(.a(G411), .O(gate129inter8));
  nand2 gate1942(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1943(.a(s_199), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1944(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1945(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1946(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2031(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2032(.a(gate132inter0), .b(s_212), .O(gate132inter1));
  and2  gate2033(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2034(.a(s_212), .O(gate132inter3));
  inv1  gate2035(.a(s_213), .O(gate132inter4));
  nand2 gate2036(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2037(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2038(.a(G416), .O(gate132inter7));
  inv1  gate2039(.a(G417), .O(gate132inter8));
  nand2 gate2040(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2041(.a(s_213), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2042(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2043(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2044(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate855(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate856(.a(gate133inter0), .b(s_44), .O(gate133inter1));
  and2  gate857(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate858(.a(s_44), .O(gate133inter3));
  inv1  gate859(.a(s_45), .O(gate133inter4));
  nand2 gate860(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate861(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate862(.a(G418), .O(gate133inter7));
  inv1  gate863(.a(G419), .O(gate133inter8));
  nand2 gate864(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate865(.a(s_45), .b(gate133inter3), .O(gate133inter10));
  nor2  gate866(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate867(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate868(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate701(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate702(.a(gate135inter0), .b(s_22), .O(gate135inter1));
  and2  gate703(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate704(.a(s_22), .O(gate135inter3));
  inv1  gate705(.a(s_23), .O(gate135inter4));
  nand2 gate706(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate707(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate708(.a(G422), .O(gate135inter7));
  inv1  gate709(.a(G423), .O(gate135inter8));
  nand2 gate710(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate711(.a(s_23), .b(gate135inter3), .O(gate135inter10));
  nor2  gate712(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate713(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate714(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate2087(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2088(.a(gate136inter0), .b(s_220), .O(gate136inter1));
  and2  gate2089(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2090(.a(s_220), .O(gate136inter3));
  inv1  gate2091(.a(s_221), .O(gate136inter4));
  nand2 gate2092(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2093(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2094(.a(G424), .O(gate136inter7));
  inv1  gate2095(.a(G425), .O(gate136inter8));
  nand2 gate2096(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2097(.a(s_221), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2098(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2099(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2100(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1485(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1486(.a(gate138inter0), .b(s_134), .O(gate138inter1));
  and2  gate1487(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1488(.a(s_134), .O(gate138inter3));
  inv1  gate1489(.a(s_135), .O(gate138inter4));
  nand2 gate1490(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1491(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1492(.a(G432), .O(gate138inter7));
  inv1  gate1493(.a(G435), .O(gate138inter8));
  nand2 gate1494(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1495(.a(s_135), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1496(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1497(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1498(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1107(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1108(.a(gate139inter0), .b(s_80), .O(gate139inter1));
  and2  gate1109(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1110(.a(s_80), .O(gate139inter3));
  inv1  gate1111(.a(s_81), .O(gate139inter4));
  nand2 gate1112(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1113(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1114(.a(G438), .O(gate139inter7));
  inv1  gate1115(.a(G441), .O(gate139inter8));
  nand2 gate1116(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1117(.a(s_81), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1118(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1119(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1120(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1261(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1262(.a(gate144inter0), .b(s_102), .O(gate144inter1));
  and2  gate1263(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1264(.a(s_102), .O(gate144inter3));
  inv1  gate1265(.a(s_103), .O(gate144inter4));
  nand2 gate1266(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1267(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1268(.a(G468), .O(gate144inter7));
  inv1  gate1269(.a(G471), .O(gate144inter8));
  nand2 gate1270(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1271(.a(s_103), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1272(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1273(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1274(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate659(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate660(.a(gate155inter0), .b(s_16), .O(gate155inter1));
  and2  gate661(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate662(.a(s_16), .O(gate155inter3));
  inv1  gate663(.a(s_17), .O(gate155inter4));
  nand2 gate664(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate665(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate666(.a(G432), .O(gate155inter7));
  inv1  gate667(.a(G525), .O(gate155inter8));
  nand2 gate668(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate669(.a(s_17), .b(gate155inter3), .O(gate155inter10));
  nor2  gate670(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate671(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate672(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate995(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate996(.a(gate157inter0), .b(s_64), .O(gate157inter1));
  and2  gate997(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate998(.a(s_64), .O(gate157inter3));
  inv1  gate999(.a(s_65), .O(gate157inter4));
  nand2 gate1000(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1001(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1002(.a(G438), .O(gate157inter7));
  inv1  gate1003(.a(G528), .O(gate157inter8));
  nand2 gate1004(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1005(.a(s_65), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1006(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1007(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1008(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2171(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2172(.a(gate160inter0), .b(s_232), .O(gate160inter1));
  and2  gate2173(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2174(.a(s_232), .O(gate160inter3));
  inv1  gate2175(.a(s_233), .O(gate160inter4));
  nand2 gate2176(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2177(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2178(.a(G447), .O(gate160inter7));
  inv1  gate2179(.a(G531), .O(gate160inter8));
  nand2 gate2180(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2181(.a(s_233), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2182(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2183(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2184(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate939(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate940(.a(gate164inter0), .b(s_56), .O(gate164inter1));
  and2  gate941(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate942(.a(s_56), .O(gate164inter3));
  inv1  gate943(.a(s_57), .O(gate164inter4));
  nand2 gate944(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate945(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate946(.a(G459), .O(gate164inter7));
  inv1  gate947(.a(G537), .O(gate164inter8));
  nand2 gate948(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate949(.a(s_57), .b(gate164inter3), .O(gate164inter10));
  nor2  gate950(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate951(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate952(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate953(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate954(.a(gate165inter0), .b(s_58), .O(gate165inter1));
  and2  gate955(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate956(.a(s_58), .O(gate165inter3));
  inv1  gate957(.a(s_59), .O(gate165inter4));
  nand2 gate958(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate959(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate960(.a(G462), .O(gate165inter7));
  inv1  gate961(.a(G540), .O(gate165inter8));
  nand2 gate962(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate963(.a(s_59), .b(gate165inter3), .O(gate165inter10));
  nor2  gate964(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate965(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate966(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1877(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1878(.a(gate170inter0), .b(s_190), .O(gate170inter1));
  and2  gate1879(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1880(.a(s_190), .O(gate170inter3));
  inv1  gate1881(.a(s_191), .O(gate170inter4));
  nand2 gate1882(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1883(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1884(.a(G477), .O(gate170inter7));
  inv1  gate1885(.a(G546), .O(gate170inter8));
  nand2 gate1886(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1887(.a(s_191), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1888(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1889(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1890(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1709(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1710(.a(gate175inter0), .b(s_166), .O(gate175inter1));
  and2  gate1711(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1712(.a(s_166), .O(gate175inter3));
  inv1  gate1713(.a(s_167), .O(gate175inter4));
  nand2 gate1714(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1715(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1716(.a(G492), .O(gate175inter7));
  inv1  gate1717(.a(G555), .O(gate175inter8));
  nand2 gate1718(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1719(.a(s_167), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1720(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1721(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1722(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1583(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1584(.a(gate178inter0), .b(s_148), .O(gate178inter1));
  and2  gate1585(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1586(.a(s_148), .O(gate178inter3));
  inv1  gate1587(.a(s_149), .O(gate178inter4));
  nand2 gate1588(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1589(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1590(.a(G501), .O(gate178inter7));
  inv1  gate1591(.a(G558), .O(gate178inter8));
  nand2 gate1592(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1593(.a(s_149), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1594(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1595(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1596(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate981(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate982(.a(gate180inter0), .b(s_62), .O(gate180inter1));
  and2  gate983(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate984(.a(s_62), .O(gate180inter3));
  inv1  gate985(.a(s_63), .O(gate180inter4));
  nand2 gate986(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate987(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate988(.a(G507), .O(gate180inter7));
  inv1  gate989(.a(G561), .O(gate180inter8));
  nand2 gate990(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate991(.a(s_63), .b(gate180inter3), .O(gate180inter10));
  nor2  gate992(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate993(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate994(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate547(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate548(.a(gate185inter0), .b(s_0), .O(gate185inter1));
  and2  gate549(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate550(.a(s_0), .O(gate185inter3));
  inv1  gate551(.a(s_1), .O(gate185inter4));
  nand2 gate552(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate553(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate554(.a(G570), .O(gate185inter7));
  inv1  gate555(.a(G571), .O(gate185inter8));
  nand2 gate556(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate557(.a(s_1), .b(gate185inter3), .O(gate185inter10));
  nor2  gate558(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate559(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate560(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1149(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1150(.a(gate186inter0), .b(s_86), .O(gate186inter1));
  and2  gate1151(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1152(.a(s_86), .O(gate186inter3));
  inv1  gate1153(.a(s_87), .O(gate186inter4));
  nand2 gate1154(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1155(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1156(.a(G572), .O(gate186inter7));
  inv1  gate1157(.a(G573), .O(gate186inter8));
  nand2 gate1158(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1159(.a(s_87), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1160(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1161(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1162(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1401(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1402(.a(gate190inter0), .b(s_122), .O(gate190inter1));
  and2  gate1403(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1404(.a(s_122), .O(gate190inter3));
  inv1  gate1405(.a(s_123), .O(gate190inter4));
  nand2 gate1406(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1407(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1408(.a(G580), .O(gate190inter7));
  inv1  gate1409(.a(G581), .O(gate190inter8));
  nand2 gate1410(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1411(.a(s_123), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1412(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1413(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1414(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1177(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1178(.a(gate191inter0), .b(s_90), .O(gate191inter1));
  and2  gate1179(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1180(.a(s_90), .O(gate191inter3));
  inv1  gate1181(.a(s_91), .O(gate191inter4));
  nand2 gate1182(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1183(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1184(.a(G582), .O(gate191inter7));
  inv1  gate1185(.a(G583), .O(gate191inter8));
  nand2 gate1186(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1187(.a(s_91), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1188(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1189(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1190(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1695(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1696(.a(gate194inter0), .b(s_164), .O(gate194inter1));
  and2  gate1697(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1698(.a(s_164), .O(gate194inter3));
  inv1  gate1699(.a(s_165), .O(gate194inter4));
  nand2 gate1700(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1701(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1702(.a(G588), .O(gate194inter7));
  inv1  gate1703(.a(G589), .O(gate194inter8));
  nand2 gate1704(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1705(.a(s_165), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1706(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1707(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1708(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate869(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate870(.a(gate195inter0), .b(s_46), .O(gate195inter1));
  and2  gate871(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate872(.a(s_46), .O(gate195inter3));
  inv1  gate873(.a(s_47), .O(gate195inter4));
  nand2 gate874(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate875(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate876(.a(G590), .O(gate195inter7));
  inv1  gate877(.a(G591), .O(gate195inter8));
  nand2 gate878(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate879(.a(s_47), .b(gate195inter3), .O(gate195inter10));
  nor2  gate880(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate881(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate882(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1457(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1458(.a(gate198inter0), .b(s_130), .O(gate198inter1));
  and2  gate1459(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1460(.a(s_130), .O(gate198inter3));
  inv1  gate1461(.a(s_131), .O(gate198inter4));
  nand2 gate1462(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1463(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1464(.a(G596), .O(gate198inter7));
  inv1  gate1465(.a(G597), .O(gate198inter8));
  nand2 gate1466(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1467(.a(s_131), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1468(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1469(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1470(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2199(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2200(.a(gate202inter0), .b(s_236), .O(gate202inter1));
  and2  gate2201(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2202(.a(s_236), .O(gate202inter3));
  inv1  gate2203(.a(s_237), .O(gate202inter4));
  nand2 gate2204(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2205(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2206(.a(G612), .O(gate202inter7));
  inv1  gate2207(.a(G617), .O(gate202inter8));
  nand2 gate2208(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2209(.a(s_237), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2210(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2211(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2212(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate715(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate716(.a(gate213inter0), .b(s_24), .O(gate213inter1));
  and2  gate717(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate718(.a(s_24), .O(gate213inter3));
  inv1  gate719(.a(s_25), .O(gate213inter4));
  nand2 gate720(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate721(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate722(.a(G602), .O(gate213inter7));
  inv1  gate723(.a(G672), .O(gate213inter8));
  nand2 gate724(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate725(.a(s_25), .b(gate213inter3), .O(gate213inter10));
  nor2  gate726(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate727(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate728(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2185(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2186(.a(gate214inter0), .b(s_234), .O(gate214inter1));
  and2  gate2187(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2188(.a(s_234), .O(gate214inter3));
  inv1  gate2189(.a(s_235), .O(gate214inter4));
  nand2 gate2190(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2191(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2192(.a(G612), .O(gate214inter7));
  inv1  gate2193(.a(G672), .O(gate214inter8));
  nand2 gate2194(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2195(.a(s_235), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2196(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2197(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2198(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1513(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1514(.a(gate219inter0), .b(s_138), .O(gate219inter1));
  and2  gate1515(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1516(.a(s_138), .O(gate219inter3));
  inv1  gate1517(.a(s_139), .O(gate219inter4));
  nand2 gate1518(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1519(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1520(.a(G632), .O(gate219inter7));
  inv1  gate1521(.a(G681), .O(gate219inter8));
  nand2 gate1522(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1523(.a(s_139), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1524(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1525(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1526(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1919(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1920(.a(gate221inter0), .b(s_196), .O(gate221inter1));
  and2  gate1921(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1922(.a(s_196), .O(gate221inter3));
  inv1  gate1923(.a(s_197), .O(gate221inter4));
  nand2 gate1924(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1925(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1926(.a(G622), .O(gate221inter7));
  inv1  gate1927(.a(G684), .O(gate221inter8));
  nand2 gate1928(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1929(.a(s_197), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1930(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1931(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1932(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1975(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1976(.a(gate224inter0), .b(s_204), .O(gate224inter1));
  and2  gate1977(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1978(.a(s_204), .O(gate224inter3));
  inv1  gate1979(.a(s_205), .O(gate224inter4));
  nand2 gate1980(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1981(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1982(.a(G637), .O(gate224inter7));
  inv1  gate1983(.a(G687), .O(gate224inter8));
  nand2 gate1984(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1985(.a(s_205), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1986(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1987(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1988(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1163(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1164(.a(gate228inter0), .b(s_88), .O(gate228inter1));
  and2  gate1165(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1166(.a(s_88), .O(gate228inter3));
  inv1  gate1167(.a(s_89), .O(gate228inter4));
  nand2 gate1168(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1169(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1170(.a(G696), .O(gate228inter7));
  inv1  gate1171(.a(G697), .O(gate228inter8));
  nand2 gate1172(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1173(.a(s_89), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1174(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1175(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1176(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1541(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1542(.a(gate230inter0), .b(s_142), .O(gate230inter1));
  and2  gate1543(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1544(.a(s_142), .O(gate230inter3));
  inv1  gate1545(.a(s_143), .O(gate230inter4));
  nand2 gate1546(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1547(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1548(.a(G700), .O(gate230inter7));
  inv1  gate1549(.a(G701), .O(gate230inter8));
  nand2 gate1550(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1551(.a(s_143), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1552(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1553(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1554(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1569(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1570(.a(gate234inter0), .b(s_146), .O(gate234inter1));
  and2  gate1571(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1572(.a(s_146), .O(gate234inter3));
  inv1  gate1573(.a(s_147), .O(gate234inter4));
  nand2 gate1574(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1575(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1576(.a(G245), .O(gate234inter7));
  inv1  gate1577(.a(G721), .O(gate234inter8));
  nand2 gate1578(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1579(.a(s_147), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1580(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1581(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1582(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1331(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1332(.a(gate235inter0), .b(s_112), .O(gate235inter1));
  and2  gate1333(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1334(.a(s_112), .O(gate235inter3));
  inv1  gate1335(.a(s_113), .O(gate235inter4));
  nand2 gate1336(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1337(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1338(.a(G248), .O(gate235inter7));
  inv1  gate1339(.a(G724), .O(gate235inter8));
  nand2 gate1340(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1341(.a(s_113), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1342(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1343(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1344(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate883(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate884(.a(gate239inter0), .b(s_48), .O(gate239inter1));
  and2  gate885(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate886(.a(s_48), .O(gate239inter3));
  inv1  gate887(.a(s_49), .O(gate239inter4));
  nand2 gate888(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate889(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate890(.a(G260), .O(gate239inter7));
  inv1  gate891(.a(G712), .O(gate239inter8));
  nand2 gate892(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate893(.a(s_49), .b(gate239inter3), .O(gate239inter10));
  nor2  gate894(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate895(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate896(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate631(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate632(.a(gate248inter0), .b(s_12), .O(gate248inter1));
  and2  gate633(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate634(.a(s_12), .O(gate248inter3));
  inv1  gate635(.a(s_13), .O(gate248inter4));
  nand2 gate636(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate637(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate638(.a(G727), .O(gate248inter7));
  inv1  gate639(.a(G739), .O(gate248inter8));
  nand2 gate640(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate641(.a(s_13), .b(gate248inter3), .O(gate248inter10));
  nor2  gate642(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate643(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate644(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1653(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1654(.a(gate250inter0), .b(s_158), .O(gate250inter1));
  and2  gate1655(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1656(.a(s_158), .O(gate250inter3));
  inv1  gate1657(.a(s_159), .O(gate250inter4));
  nand2 gate1658(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1659(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1660(.a(G706), .O(gate250inter7));
  inv1  gate1661(.a(G742), .O(gate250inter8));
  nand2 gate1662(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1663(.a(s_159), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1664(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1665(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1666(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1807(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1808(.a(gate253inter0), .b(s_180), .O(gate253inter1));
  and2  gate1809(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1810(.a(s_180), .O(gate253inter3));
  inv1  gate1811(.a(s_181), .O(gate253inter4));
  nand2 gate1812(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1813(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1814(.a(G260), .O(gate253inter7));
  inv1  gate1815(.a(G748), .O(gate253inter8));
  nand2 gate1816(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1817(.a(s_181), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1818(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1819(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1820(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1779(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1780(.a(gate255inter0), .b(s_176), .O(gate255inter1));
  and2  gate1781(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1782(.a(s_176), .O(gate255inter3));
  inv1  gate1783(.a(s_177), .O(gate255inter4));
  nand2 gate1784(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1785(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1786(.a(G263), .O(gate255inter7));
  inv1  gate1787(.a(G751), .O(gate255inter8));
  nand2 gate1788(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1789(.a(s_177), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1790(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1791(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1792(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1135(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1136(.a(gate261inter0), .b(s_84), .O(gate261inter1));
  and2  gate1137(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1138(.a(s_84), .O(gate261inter3));
  inv1  gate1139(.a(s_85), .O(gate261inter4));
  nand2 gate1140(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1141(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1142(.a(G762), .O(gate261inter7));
  inv1  gate1143(.a(G763), .O(gate261inter8));
  nand2 gate1144(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1145(.a(s_85), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1146(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1147(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1148(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1303(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1304(.a(gate262inter0), .b(s_108), .O(gate262inter1));
  and2  gate1305(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1306(.a(s_108), .O(gate262inter3));
  inv1  gate1307(.a(s_109), .O(gate262inter4));
  nand2 gate1308(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1309(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1310(.a(G764), .O(gate262inter7));
  inv1  gate1311(.a(G765), .O(gate262inter8));
  nand2 gate1312(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1313(.a(s_109), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1314(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1315(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1316(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1611(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1612(.a(gate265inter0), .b(s_152), .O(gate265inter1));
  and2  gate1613(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1614(.a(s_152), .O(gate265inter3));
  inv1  gate1615(.a(s_153), .O(gate265inter4));
  nand2 gate1616(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1617(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1618(.a(G642), .O(gate265inter7));
  inv1  gate1619(.a(G770), .O(gate265inter8));
  nand2 gate1620(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1621(.a(s_153), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1622(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1623(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1624(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate561(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate562(.a(gate266inter0), .b(s_2), .O(gate266inter1));
  and2  gate563(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate564(.a(s_2), .O(gate266inter3));
  inv1  gate565(.a(s_3), .O(gate266inter4));
  nand2 gate566(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate567(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate568(.a(G645), .O(gate266inter7));
  inv1  gate569(.a(G773), .O(gate266inter8));
  nand2 gate570(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate571(.a(s_3), .b(gate266inter3), .O(gate266inter10));
  nor2  gate572(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate573(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate574(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1639(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1640(.a(gate268inter0), .b(s_156), .O(gate268inter1));
  and2  gate1641(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1642(.a(s_156), .O(gate268inter3));
  inv1  gate1643(.a(s_157), .O(gate268inter4));
  nand2 gate1644(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1645(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1646(.a(G651), .O(gate268inter7));
  inv1  gate1647(.a(G779), .O(gate268inter8));
  nand2 gate1648(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1649(.a(s_157), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1650(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1651(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1652(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1961(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1962(.a(gate269inter0), .b(s_202), .O(gate269inter1));
  and2  gate1963(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1964(.a(s_202), .O(gate269inter3));
  inv1  gate1965(.a(s_203), .O(gate269inter4));
  nand2 gate1966(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1967(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1968(.a(G654), .O(gate269inter7));
  inv1  gate1969(.a(G782), .O(gate269inter8));
  nand2 gate1970(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1971(.a(s_203), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1972(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1973(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1974(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate785(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate786(.a(gate271inter0), .b(s_34), .O(gate271inter1));
  and2  gate787(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate788(.a(s_34), .O(gate271inter3));
  inv1  gate789(.a(s_35), .O(gate271inter4));
  nand2 gate790(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate791(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate792(.a(G660), .O(gate271inter7));
  inv1  gate793(.a(G788), .O(gate271inter8));
  nand2 gate794(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate795(.a(s_35), .b(gate271inter3), .O(gate271inter10));
  nor2  gate796(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate797(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate798(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1079(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1080(.a(gate277inter0), .b(s_76), .O(gate277inter1));
  and2  gate1081(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1082(.a(s_76), .O(gate277inter3));
  inv1  gate1083(.a(s_77), .O(gate277inter4));
  nand2 gate1084(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1085(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1086(.a(G648), .O(gate277inter7));
  inv1  gate1087(.a(G800), .O(gate277inter8));
  nand2 gate1088(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1089(.a(s_77), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1090(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1091(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1092(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate575(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate576(.a(gate278inter0), .b(s_4), .O(gate278inter1));
  and2  gate577(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate578(.a(s_4), .O(gate278inter3));
  inv1  gate579(.a(s_5), .O(gate278inter4));
  nand2 gate580(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate581(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate582(.a(G776), .O(gate278inter7));
  inv1  gate583(.a(G800), .O(gate278inter8));
  nand2 gate584(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate585(.a(s_5), .b(gate278inter3), .O(gate278inter10));
  nor2  gate586(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate587(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate588(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1065(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1066(.a(gate279inter0), .b(s_74), .O(gate279inter1));
  and2  gate1067(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1068(.a(s_74), .O(gate279inter3));
  inv1  gate1069(.a(s_75), .O(gate279inter4));
  nand2 gate1070(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1071(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1072(.a(G651), .O(gate279inter7));
  inv1  gate1073(.a(G803), .O(gate279inter8));
  nand2 gate1074(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1075(.a(s_75), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1076(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1077(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1078(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1191(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1192(.a(gate281inter0), .b(s_92), .O(gate281inter1));
  and2  gate1193(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1194(.a(s_92), .O(gate281inter3));
  inv1  gate1195(.a(s_93), .O(gate281inter4));
  nand2 gate1196(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1197(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1198(.a(G654), .O(gate281inter7));
  inv1  gate1199(.a(G806), .O(gate281inter8));
  nand2 gate1200(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1201(.a(s_93), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1202(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1203(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1204(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate673(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate674(.a(gate283inter0), .b(s_18), .O(gate283inter1));
  and2  gate675(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate676(.a(s_18), .O(gate283inter3));
  inv1  gate677(.a(s_19), .O(gate283inter4));
  nand2 gate678(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate679(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate680(.a(G657), .O(gate283inter7));
  inv1  gate681(.a(G809), .O(gate283inter8));
  nand2 gate682(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate683(.a(s_19), .b(gate283inter3), .O(gate283inter10));
  nor2  gate684(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate685(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate686(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1737(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1738(.a(gate287inter0), .b(s_170), .O(gate287inter1));
  and2  gate1739(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1740(.a(s_170), .O(gate287inter3));
  inv1  gate1741(.a(s_171), .O(gate287inter4));
  nand2 gate1742(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1743(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1744(.a(G663), .O(gate287inter7));
  inv1  gate1745(.a(G815), .O(gate287inter8));
  nand2 gate1746(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1747(.a(s_171), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1748(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1749(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1750(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1681(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1682(.a(gate293inter0), .b(s_162), .O(gate293inter1));
  and2  gate1683(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1684(.a(s_162), .O(gate293inter3));
  inv1  gate1685(.a(s_163), .O(gate293inter4));
  nand2 gate1686(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1687(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1688(.a(G828), .O(gate293inter7));
  inv1  gate1689(.a(G829), .O(gate293inter8));
  nand2 gate1690(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1691(.a(s_163), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1692(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1693(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1694(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1051(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1052(.a(gate295inter0), .b(s_72), .O(gate295inter1));
  and2  gate1053(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1054(.a(s_72), .O(gate295inter3));
  inv1  gate1055(.a(s_73), .O(gate295inter4));
  nand2 gate1056(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1057(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1058(.a(G830), .O(gate295inter7));
  inv1  gate1059(.a(G831), .O(gate295inter8));
  nand2 gate1060(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1061(.a(s_73), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1062(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1063(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1064(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1345(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1346(.a(gate391inter0), .b(s_114), .O(gate391inter1));
  and2  gate1347(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1348(.a(s_114), .O(gate391inter3));
  inv1  gate1349(.a(s_115), .O(gate391inter4));
  nand2 gate1350(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1351(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1352(.a(G5), .O(gate391inter7));
  inv1  gate1353(.a(G1048), .O(gate391inter8));
  nand2 gate1354(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1355(.a(s_115), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1356(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1357(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1358(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1625(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1626(.a(gate393inter0), .b(s_154), .O(gate393inter1));
  and2  gate1627(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1628(.a(s_154), .O(gate393inter3));
  inv1  gate1629(.a(s_155), .O(gate393inter4));
  nand2 gate1630(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1631(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1632(.a(G7), .O(gate393inter7));
  inv1  gate1633(.a(G1054), .O(gate393inter8));
  nand2 gate1634(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1635(.a(s_155), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1636(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1637(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1638(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate757(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate758(.a(gate397inter0), .b(s_30), .O(gate397inter1));
  and2  gate759(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate760(.a(s_30), .O(gate397inter3));
  inv1  gate761(.a(s_31), .O(gate397inter4));
  nand2 gate762(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate763(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate764(.a(G11), .O(gate397inter7));
  inv1  gate765(.a(G1066), .O(gate397inter8));
  nand2 gate766(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate767(.a(s_31), .b(gate397inter3), .O(gate397inter10));
  nor2  gate768(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate769(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate770(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2045(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2046(.a(gate400inter0), .b(s_214), .O(gate400inter1));
  and2  gate2047(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2048(.a(s_214), .O(gate400inter3));
  inv1  gate2049(.a(s_215), .O(gate400inter4));
  nand2 gate2050(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2051(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2052(.a(G14), .O(gate400inter7));
  inv1  gate2053(.a(G1075), .O(gate400inter8));
  nand2 gate2054(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2055(.a(s_215), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2056(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2057(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2058(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1205(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1206(.a(gate403inter0), .b(s_94), .O(gate403inter1));
  and2  gate1207(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1208(.a(s_94), .O(gate403inter3));
  inv1  gate1209(.a(s_95), .O(gate403inter4));
  nand2 gate1210(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1211(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1212(.a(G17), .O(gate403inter7));
  inv1  gate1213(.a(G1084), .O(gate403inter8));
  nand2 gate1214(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1215(.a(s_95), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1216(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1217(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1218(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate645(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate646(.a(gate408inter0), .b(s_14), .O(gate408inter1));
  and2  gate647(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate648(.a(s_14), .O(gate408inter3));
  inv1  gate649(.a(s_15), .O(gate408inter4));
  nand2 gate650(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate651(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate652(.a(G22), .O(gate408inter7));
  inv1  gate653(.a(G1099), .O(gate408inter8));
  nand2 gate654(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate655(.a(s_15), .b(gate408inter3), .O(gate408inter10));
  nor2  gate656(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate657(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate658(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2227(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2228(.a(gate410inter0), .b(s_240), .O(gate410inter1));
  and2  gate2229(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2230(.a(s_240), .O(gate410inter3));
  inv1  gate2231(.a(s_241), .O(gate410inter4));
  nand2 gate2232(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2233(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2234(.a(G24), .O(gate410inter7));
  inv1  gate2235(.a(G1105), .O(gate410inter8));
  nand2 gate2236(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2237(.a(s_241), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2238(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2239(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2240(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1289(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1290(.a(gate417inter0), .b(s_106), .O(gate417inter1));
  and2  gate1291(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1292(.a(s_106), .O(gate417inter3));
  inv1  gate1293(.a(s_107), .O(gate417inter4));
  nand2 gate1294(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1295(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1296(.a(G31), .O(gate417inter7));
  inv1  gate1297(.a(G1126), .O(gate417inter8));
  nand2 gate1298(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1299(.a(s_107), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1300(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1301(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1302(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate729(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate730(.a(gate419inter0), .b(s_26), .O(gate419inter1));
  and2  gate731(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate732(.a(s_26), .O(gate419inter3));
  inv1  gate733(.a(s_27), .O(gate419inter4));
  nand2 gate734(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate735(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate736(.a(G1), .O(gate419inter7));
  inv1  gate737(.a(G1132), .O(gate419inter8));
  nand2 gate738(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate739(.a(s_27), .b(gate419inter3), .O(gate419inter10));
  nor2  gate740(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate741(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate742(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2115(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2116(.a(gate422inter0), .b(s_224), .O(gate422inter1));
  and2  gate2117(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2118(.a(s_224), .O(gate422inter3));
  inv1  gate2119(.a(s_225), .O(gate422inter4));
  nand2 gate2120(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2121(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2122(.a(G1039), .O(gate422inter7));
  inv1  gate2123(.a(G1135), .O(gate422inter8));
  nand2 gate2124(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2125(.a(s_225), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2126(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2127(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2128(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate813(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate814(.a(gate427inter0), .b(s_38), .O(gate427inter1));
  and2  gate815(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate816(.a(s_38), .O(gate427inter3));
  inv1  gate817(.a(s_39), .O(gate427inter4));
  nand2 gate818(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate819(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate820(.a(G5), .O(gate427inter7));
  inv1  gate821(.a(G1144), .O(gate427inter8));
  nand2 gate822(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate823(.a(s_39), .b(gate427inter3), .O(gate427inter10));
  nor2  gate824(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate825(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate826(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate967(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate968(.a(gate430inter0), .b(s_60), .O(gate430inter1));
  and2  gate969(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate970(.a(s_60), .O(gate430inter3));
  inv1  gate971(.a(s_61), .O(gate430inter4));
  nand2 gate972(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate973(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate974(.a(G1051), .O(gate430inter7));
  inv1  gate975(.a(G1147), .O(gate430inter8));
  nand2 gate976(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate977(.a(s_61), .b(gate430inter3), .O(gate430inter10));
  nor2  gate978(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate979(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate980(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1443(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1444(.a(gate434inter0), .b(s_128), .O(gate434inter1));
  and2  gate1445(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1446(.a(s_128), .O(gate434inter3));
  inv1  gate1447(.a(s_129), .O(gate434inter4));
  nand2 gate1448(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1449(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1450(.a(G1057), .O(gate434inter7));
  inv1  gate1451(.a(G1153), .O(gate434inter8));
  nand2 gate1452(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1453(.a(s_129), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1454(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1455(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1456(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1905(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1906(.a(gate435inter0), .b(s_194), .O(gate435inter1));
  and2  gate1907(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1908(.a(s_194), .O(gate435inter3));
  inv1  gate1909(.a(s_195), .O(gate435inter4));
  nand2 gate1910(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1911(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1912(.a(G9), .O(gate435inter7));
  inv1  gate1913(.a(G1156), .O(gate435inter8));
  nand2 gate1914(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1915(.a(s_195), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1916(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1917(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1918(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate687(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate688(.a(gate438inter0), .b(s_20), .O(gate438inter1));
  and2  gate689(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate690(.a(s_20), .O(gate438inter3));
  inv1  gate691(.a(s_21), .O(gate438inter4));
  nand2 gate692(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate693(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate694(.a(G1063), .O(gate438inter7));
  inv1  gate695(.a(G1159), .O(gate438inter8));
  nand2 gate696(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate697(.a(s_21), .b(gate438inter3), .O(gate438inter10));
  nor2  gate698(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate699(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate700(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2157(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2158(.a(gate442inter0), .b(s_230), .O(gate442inter1));
  and2  gate2159(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2160(.a(s_230), .O(gate442inter3));
  inv1  gate2161(.a(s_231), .O(gate442inter4));
  nand2 gate2162(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2163(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2164(.a(G1069), .O(gate442inter7));
  inv1  gate2165(.a(G1165), .O(gate442inter8));
  nand2 gate2166(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2167(.a(s_231), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2168(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2169(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2170(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate2129(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2130(.a(gate443inter0), .b(s_226), .O(gate443inter1));
  and2  gate2131(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2132(.a(s_226), .O(gate443inter3));
  inv1  gate2133(.a(s_227), .O(gate443inter4));
  nand2 gate2134(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2135(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2136(.a(G13), .O(gate443inter7));
  inv1  gate2137(.a(G1168), .O(gate443inter8));
  nand2 gate2138(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2139(.a(s_227), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2140(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2141(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2142(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1429(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1430(.a(gate445inter0), .b(s_126), .O(gate445inter1));
  and2  gate1431(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1432(.a(s_126), .O(gate445inter3));
  inv1  gate1433(.a(s_127), .O(gate445inter4));
  nand2 gate1434(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1435(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1436(.a(G14), .O(gate445inter7));
  inv1  gate1437(.a(G1171), .O(gate445inter8));
  nand2 gate1438(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1439(.a(s_127), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1440(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1441(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1442(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1667(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1668(.a(gate449inter0), .b(s_160), .O(gate449inter1));
  and2  gate1669(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1670(.a(s_160), .O(gate449inter3));
  inv1  gate1671(.a(s_161), .O(gate449inter4));
  nand2 gate1672(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1673(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1674(.a(G16), .O(gate449inter7));
  inv1  gate1675(.a(G1177), .O(gate449inter8));
  nand2 gate1676(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1677(.a(s_161), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1678(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1679(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1680(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1891(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1892(.a(gate451inter0), .b(s_192), .O(gate451inter1));
  and2  gate1893(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1894(.a(s_192), .O(gate451inter3));
  inv1  gate1895(.a(s_193), .O(gate451inter4));
  nand2 gate1896(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1897(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1898(.a(G17), .O(gate451inter7));
  inv1  gate1899(.a(G1180), .O(gate451inter8));
  nand2 gate1900(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1901(.a(s_193), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1902(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1903(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1904(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1317(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1318(.a(gate457inter0), .b(s_110), .O(gate457inter1));
  and2  gate1319(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1320(.a(s_110), .O(gate457inter3));
  inv1  gate1321(.a(s_111), .O(gate457inter4));
  nand2 gate1322(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1323(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1324(.a(G20), .O(gate457inter7));
  inv1  gate1325(.a(G1189), .O(gate457inter8));
  nand2 gate1326(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1327(.a(s_111), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1328(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1329(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1330(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1947(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1948(.a(gate462inter0), .b(s_200), .O(gate462inter1));
  and2  gate1949(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1950(.a(s_200), .O(gate462inter3));
  inv1  gate1951(.a(s_201), .O(gate462inter4));
  nand2 gate1952(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1953(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1954(.a(G1099), .O(gate462inter7));
  inv1  gate1955(.a(G1195), .O(gate462inter8));
  nand2 gate1956(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1957(.a(s_201), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1958(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1959(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1960(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1849(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1850(.a(gate465inter0), .b(s_186), .O(gate465inter1));
  and2  gate1851(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1852(.a(s_186), .O(gate465inter3));
  inv1  gate1853(.a(s_187), .O(gate465inter4));
  nand2 gate1854(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1855(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1856(.a(G24), .O(gate465inter7));
  inv1  gate1857(.a(G1201), .O(gate465inter8));
  nand2 gate1858(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1859(.a(s_187), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1860(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1861(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1862(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2143(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2144(.a(gate467inter0), .b(s_228), .O(gate467inter1));
  and2  gate2145(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2146(.a(s_228), .O(gate467inter3));
  inv1  gate2147(.a(s_229), .O(gate467inter4));
  nand2 gate2148(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2149(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2150(.a(G25), .O(gate467inter7));
  inv1  gate2151(.a(G1204), .O(gate467inter8));
  nand2 gate2152(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2153(.a(s_229), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2154(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2155(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2156(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate617(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate618(.a(gate478inter0), .b(s_10), .O(gate478inter1));
  and2  gate619(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate620(.a(s_10), .O(gate478inter3));
  inv1  gate621(.a(s_11), .O(gate478inter4));
  nand2 gate622(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate623(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate624(.a(G1123), .O(gate478inter7));
  inv1  gate625(.a(G1219), .O(gate478inter8));
  nand2 gate626(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate627(.a(s_11), .b(gate478inter3), .O(gate478inter10));
  nor2  gate628(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate629(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate630(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1275(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1276(.a(gate479inter0), .b(s_104), .O(gate479inter1));
  and2  gate1277(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1278(.a(s_104), .O(gate479inter3));
  inv1  gate1279(.a(s_105), .O(gate479inter4));
  nand2 gate1280(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1281(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1282(.a(G31), .O(gate479inter7));
  inv1  gate1283(.a(G1222), .O(gate479inter8));
  nand2 gate1284(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1285(.a(s_105), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1286(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1287(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1288(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1527(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1528(.a(gate480inter0), .b(s_140), .O(gate480inter1));
  and2  gate1529(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1530(.a(s_140), .O(gate480inter3));
  inv1  gate1531(.a(s_141), .O(gate480inter4));
  nand2 gate1532(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1533(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1534(.a(G1126), .O(gate480inter7));
  inv1  gate1535(.a(G1222), .O(gate480inter8));
  nand2 gate1536(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1537(.a(s_141), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1538(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1539(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1540(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2213(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2214(.a(gate482inter0), .b(s_238), .O(gate482inter1));
  and2  gate2215(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2216(.a(s_238), .O(gate482inter3));
  inv1  gate2217(.a(s_239), .O(gate482inter4));
  nand2 gate2218(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2219(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2220(.a(G1129), .O(gate482inter7));
  inv1  gate2221(.a(G1225), .O(gate482inter8));
  nand2 gate2222(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2223(.a(s_239), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2224(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2225(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2226(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate799(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate800(.a(gate483inter0), .b(s_36), .O(gate483inter1));
  and2  gate801(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate802(.a(s_36), .O(gate483inter3));
  inv1  gate803(.a(s_37), .O(gate483inter4));
  nand2 gate804(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate805(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate806(.a(G1228), .O(gate483inter7));
  inv1  gate807(.a(G1229), .O(gate483inter8));
  nand2 gate808(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate809(.a(s_37), .b(gate483inter3), .O(gate483inter10));
  nor2  gate810(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate811(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate812(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1415(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1416(.a(gate485inter0), .b(s_124), .O(gate485inter1));
  and2  gate1417(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1418(.a(s_124), .O(gate485inter3));
  inv1  gate1419(.a(s_125), .O(gate485inter4));
  nand2 gate1420(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1421(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1422(.a(G1232), .O(gate485inter7));
  inv1  gate1423(.a(G1233), .O(gate485inter8));
  nand2 gate1424(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1425(.a(s_125), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1426(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1427(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1428(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate603(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate604(.a(gate486inter0), .b(s_8), .O(gate486inter1));
  and2  gate605(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate606(.a(s_8), .O(gate486inter3));
  inv1  gate607(.a(s_9), .O(gate486inter4));
  nand2 gate608(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate609(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate610(.a(G1234), .O(gate486inter7));
  inv1  gate611(.a(G1235), .O(gate486inter8));
  nand2 gate612(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate613(.a(s_9), .b(gate486inter3), .O(gate486inter10));
  nor2  gate614(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate615(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate616(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1037(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1038(.a(gate487inter0), .b(s_70), .O(gate487inter1));
  and2  gate1039(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1040(.a(s_70), .O(gate487inter3));
  inv1  gate1041(.a(s_71), .O(gate487inter4));
  nand2 gate1042(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1043(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1044(.a(G1236), .O(gate487inter7));
  inv1  gate1045(.a(G1237), .O(gate487inter8));
  nand2 gate1046(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1047(.a(s_71), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1048(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1049(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1050(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1471(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1472(.a(gate494inter0), .b(s_132), .O(gate494inter1));
  and2  gate1473(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1474(.a(s_132), .O(gate494inter3));
  inv1  gate1475(.a(s_133), .O(gate494inter4));
  nand2 gate1476(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1477(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1478(.a(G1250), .O(gate494inter7));
  inv1  gate1479(.a(G1251), .O(gate494inter8));
  nand2 gate1480(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1481(.a(s_133), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1482(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1483(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1484(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1219(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1220(.a(gate501inter0), .b(s_96), .O(gate501inter1));
  and2  gate1221(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1222(.a(s_96), .O(gate501inter3));
  inv1  gate1223(.a(s_97), .O(gate501inter4));
  nand2 gate1224(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1225(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1226(.a(G1264), .O(gate501inter7));
  inv1  gate1227(.a(G1265), .O(gate501inter8));
  nand2 gate1228(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1229(.a(s_97), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1230(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1231(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1232(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2003(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2004(.a(gate502inter0), .b(s_208), .O(gate502inter1));
  and2  gate2005(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2006(.a(s_208), .O(gate502inter3));
  inv1  gate2007(.a(s_209), .O(gate502inter4));
  nand2 gate2008(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2009(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2010(.a(G1266), .O(gate502inter7));
  inv1  gate2011(.a(G1267), .O(gate502inter8));
  nand2 gate2012(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2013(.a(s_209), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2014(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2015(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2016(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate589(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate590(.a(gate509inter0), .b(s_6), .O(gate509inter1));
  and2  gate591(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate592(.a(s_6), .O(gate509inter3));
  inv1  gate593(.a(s_7), .O(gate509inter4));
  nand2 gate594(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate595(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate596(.a(G1280), .O(gate509inter7));
  inv1  gate597(.a(G1281), .O(gate509inter8));
  nand2 gate598(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate599(.a(s_7), .b(gate509inter3), .O(gate509inter10));
  nor2  gate600(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate601(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate602(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1723(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1724(.a(gate511inter0), .b(s_168), .O(gate511inter1));
  and2  gate1725(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1726(.a(s_168), .O(gate511inter3));
  inv1  gate1727(.a(s_169), .O(gate511inter4));
  nand2 gate1728(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1729(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1730(.a(G1284), .O(gate511inter7));
  inv1  gate1731(.a(G1285), .O(gate511inter8));
  nand2 gate1732(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1733(.a(s_169), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1734(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1735(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1736(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1863(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1864(.a(gate514inter0), .b(s_188), .O(gate514inter1));
  and2  gate1865(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1866(.a(s_188), .O(gate514inter3));
  inv1  gate1867(.a(s_189), .O(gate514inter4));
  nand2 gate1868(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1869(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1870(.a(G1290), .O(gate514inter7));
  inv1  gate1871(.a(G1291), .O(gate514inter8));
  nand2 gate1872(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1873(.a(s_189), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1874(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1875(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1876(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule