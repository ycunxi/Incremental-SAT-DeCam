module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1541(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1542(.a(gate10inter0), .b(s_142), .O(gate10inter1));
  and2  gate1543(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1544(.a(s_142), .O(gate10inter3));
  inv1  gate1545(.a(s_143), .O(gate10inter4));
  nand2 gate1546(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1547(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1548(.a(G3), .O(gate10inter7));
  inv1  gate1549(.a(G4), .O(gate10inter8));
  nand2 gate1550(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1551(.a(s_143), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1552(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1553(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1554(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate1919(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1920(.a(gate11inter0), .b(s_196), .O(gate11inter1));
  and2  gate1921(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1922(.a(s_196), .O(gate11inter3));
  inv1  gate1923(.a(s_197), .O(gate11inter4));
  nand2 gate1924(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1925(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1926(.a(G5), .O(gate11inter7));
  inv1  gate1927(.a(G6), .O(gate11inter8));
  nand2 gate1928(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1929(.a(s_197), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1930(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1931(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1932(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1121(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1122(.a(gate13inter0), .b(s_82), .O(gate13inter1));
  and2  gate1123(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1124(.a(s_82), .O(gate13inter3));
  inv1  gate1125(.a(s_83), .O(gate13inter4));
  nand2 gate1126(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1127(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1128(.a(G9), .O(gate13inter7));
  inv1  gate1129(.a(G10), .O(gate13inter8));
  nand2 gate1130(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1131(.a(s_83), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1132(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1133(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1134(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2395(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2396(.a(gate15inter0), .b(s_264), .O(gate15inter1));
  and2  gate2397(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2398(.a(s_264), .O(gate15inter3));
  inv1  gate2399(.a(s_265), .O(gate15inter4));
  nand2 gate2400(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2401(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2402(.a(G13), .O(gate15inter7));
  inv1  gate2403(.a(G14), .O(gate15inter8));
  nand2 gate2404(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2405(.a(s_265), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2406(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2407(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2408(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2031(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2032(.a(gate16inter0), .b(s_212), .O(gate16inter1));
  and2  gate2033(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2034(.a(s_212), .O(gate16inter3));
  inv1  gate2035(.a(s_213), .O(gate16inter4));
  nand2 gate2036(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2037(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2038(.a(G15), .O(gate16inter7));
  inv1  gate2039(.a(G16), .O(gate16inter8));
  nand2 gate2040(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2041(.a(s_213), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2042(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2043(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2044(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate757(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate758(.a(gate21inter0), .b(s_30), .O(gate21inter1));
  and2  gate759(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate760(.a(s_30), .O(gate21inter3));
  inv1  gate761(.a(s_31), .O(gate21inter4));
  nand2 gate762(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate763(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate764(.a(G25), .O(gate21inter7));
  inv1  gate765(.a(G26), .O(gate21inter8));
  nand2 gate766(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate767(.a(s_31), .b(gate21inter3), .O(gate21inter10));
  nor2  gate768(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate769(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate770(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1513(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1514(.a(gate30inter0), .b(s_138), .O(gate30inter1));
  and2  gate1515(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1516(.a(s_138), .O(gate30inter3));
  inv1  gate1517(.a(s_139), .O(gate30inter4));
  nand2 gate1518(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1519(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1520(.a(G11), .O(gate30inter7));
  inv1  gate1521(.a(G15), .O(gate30inter8));
  nand2 gate1522(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1523(.a(s_139), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1524(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1525(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1526(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate925(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate926(.a(gate36inter0), .b(s_54), .O(gate36inter1));
  and2  gate927(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate928(.a(s_54), .O(gate36inter3));
  inv1  gate929(.a(s_55), .O(gate36inter4));
  nand2 gate930(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate931(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate932(.a(G26), .O(gate36inter7));
  inv1  gate933(.a(G30), .O(gate36inter8));
  nand2 gate934(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate935(.a(s_55), .b(gate36inter3), .O(gate36inter10));
  nor2  gate936(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate937(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate938(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate911(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate912(.a(gate40inter0), .b(s_52), .O(gate40inter1));
  and2  gate913(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate914(.a(s_52), .O(gate40inter3));
  inv1  gate915(.a(s_53), .O(gate40inter4));
  nand2 gate916(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate917(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate918(.a(G28), .O(gate40inter7));
  inv1  gate919(.a(G32), .O(gate40inter8));
  nand2 gate920(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate921(.a(s_53), .b(gate40inter3), .O(gate40inter10));
  nor2  gate922(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate923(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate924(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1303(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1304(.a(gate41inter0), .b(s_108), .O(gate41inter1));
  and2  gate1305(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1306(.a(s_108), .O(gate41inter3));
  inv1  gate1307(.a(s_109), .O(gate41inter4));
  nand2 gate1308(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1309(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1310(.a(G1), .O(gate41inter7));
  inv1  gate1311(.a(G266), .O(gate41inter8));
  nand2 gate1312(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1313(.a(s_109), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1314(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1315(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1316(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate645(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate646(.a(gate44inter0), .b(s_14), .O(gate44inter1));
  and2  gate647(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate648(.a(s_14), .O(gate44inter3));
  inv1  gate649(.a(s_15), .O(gate44inter4));
  nand2 gate650(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate651(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate652(.a(G4), .O(gate44inter7));
  inv1  gate653(.a(G269), .O(gate44inter8));
  nand2 gate654(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate655(.a(s_15), .b(gate44inter3), .O(gate44inter10));
  nor2  gate656(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate657(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate658(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1009(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1010(.a(gate50inter0), .b(s_66), .O(gate50inter1));
  and2  gate1011(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1012(.a(s_66), .O(gate50inter3));
  inv1  gate1013(.a(s_67), .O(gate50inter4));
  nand2 gate1014(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1015(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1016(.a(G10), .O(gate50inter7));
  inv1  gate1017(.a(G278), .O(gate50inter8));
  nand2 gate1018(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1019(.a(s_67), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1020(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1021(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1022(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1247(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1248(.a(gate55inter0), .b(s_100), .O(gate55inter1));
  and2  gate1249(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1250(.a(s_100), .O(gate55inter3));
  inv1  gate1251(.a(s_101), .O(gate55inter4));
  nand2 gate1252(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1253(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1254(.a(G15), .O(gate55inter7));
  inv1  gate1255(.a(G287), .O(gate55inter8));
  nand2 gate1256(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1257(.a(s_101), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1258(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1259(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1260(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate743(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate744(.a(gate58inter0), .b(s_28), .O(gate58inter1));
  and2  gate745(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate746(.a(s_28), .O(gate58inter3));
  inv1  gate747(.a(s_29), .O(gate58inter4));
  nand2 gate748(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate749(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate750(.a(G18), .O(gate58inter7));
  inv1  gate751(.a(G290), .O(gate58inter8));
  nand2 gate752(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate753(.a(s_29), .b(gate58inter3), .O(gate58inter10));
  nor2  gate754(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate755(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate756(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1471(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1472(.a(gate60inter0), .b(s_132), .O(gate60inter1));
  and2  gate1473(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1474(.a(s_132), .O(gate60inter3));
  inv1  gate1475(.a(s_133), .O(gate60inter4));
  nand2 gate1476(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1477(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1478(.a(G20), .O(gate60inter7));
  inv1  gate1479(.a(G293), .O(gate60inter8));
  nand2 gate1480(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1481(.a(s_133), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1482(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1483(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1484(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1023(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1024(.a(gate61inter0), .b(s_68), .O(gate61inter1));
  and2  gate1025(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1026(.a(s_68), .O(gate61inter3));
  inv1  gate1027(.a(s_69), .O(gate61inter4));
  nand2 gate1028(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1029(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1030(.a(G21), .O(gate61inter7));
  inv1  gate1031(.a(G296), .O(gate61inter8));
  nand2 gate1032(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1033(.a(s_69), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1034(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1035(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1036(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1443(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1444(.a(gate62inter0), .b(s_128), .O(gate62inter1));
  and2  gate1445(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1446(.a(s_128), .O(gate62inter3));
  inv1  gate1447(.a(s_129), .O(gate62inter4));
  nand2 gate1448(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1449(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1450(.a(G22), .O(gate62inter7));
  inv1  gate1451(.a(G296), .O(gate62inter8));
  nand2 gate1452(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1453(.a(s_129), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1454(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1455(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1456(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2241(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2242(.a(gate71inter0), .b(s_242), .O(gate71inter1));
  and2  gate2243(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2244(.a(s_242), .O(gate71inter3));
  inv1  gate2245(.a(s_243), .O(gate71inter4));
  nand2 gate2246(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2247(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2248(.a(G31), .O(gate71inter7));
  inv1  gate2249(.a(G311), .O(gate71inter8));
  nand2 gate2250(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2251(.a(s_243), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2252(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2253(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2254(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1373(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1374(.a(gate73inter0), .b(s_118), .O(gate73inter1));
  and2  gate1375(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1376(.a(s_118), .O(gate73inter3));
  inv1  gate1377(.a(s_119), .O(gate73inter4));
  nand2 gate1378(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1379(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1380(.a(G1), .O(gate73inter7));
  inv1  gate1381(.a(G314), .O(gate73inter8));
  nand2 gate1382(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1383(.a(s_119), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1384(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1385(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1386(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate785(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate786(.a(gate76inter0), .b(s_34), .O(gate76inter1));
  and2  gate787(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate788(.a(s_34), .O(gate76inter3));
  inv1  gate789(.a(s_35), .O(gate76inter4));
  nand2 gate790(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate791(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate792(.a(G13), .O(gate76inter7));
  inv1  gate793(.a(G317), .O(gate76inter8));
  nand2 gate794(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate795(.a(s_35), .b(gate76inter3), .O(gate76inter10));
  nor2  gate796(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate797(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate798(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1065(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1066(.a(gate77inter0), .b(s_74), .O(gate77inter1));
  and2  gate1067(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1068(.a(s_74), .O(gate77inter3));
  inv1  gate1069(.a(s_75), .O(gate77inter4));
  nand2 gate1070(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1071(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1072(.a(G2), .O(gate77inter7));
  inv1  gate1073(.a(G320), .O(gate77inter8));
  nand2 gate1074(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1075(.a(s_75), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1076(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1077(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1078(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate771(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate772(.a(gate80inter0), .b(s_32), .O(gate80inter1));
  and2  gate773(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate774(.a(s_32), .O(gate80inter3));
  inv1  gate775(.a(s_33), .O(gate80inter4));
  nand2 gate776(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate777(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate778(.a(G14), .O(gate80inter7));
  inv1  gate779(.a(G323), .O(gate80inter8));
  nand2 gate780(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate781(.a(s_33), .b(gate80inter3), .O(gate80inter10));
  nor2  gate782(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate783(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate784(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2087(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2088(.a(gate81inter0), .b(s_220), .O(gate81inter1));
  and2  gate2089(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2090(.a(s_220), .O(gate81inter3));
  inv1  gate2091(.a(s_221), .O(gate81inter4));
  nand2 gate2092(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2093(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2094(.a(G3), .O(gate81inter7));
  inv1  gate2095(.a(G326), .O(gate81inter8));
  nand2 gate2096(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2097(.a(s_221), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2098(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2099(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2100(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1863(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1864(.a(gate86inter0), .b(s_188), .O(gate86inter1));
  and2  gate1865(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1866(.a(s_188), .O(gate86inter3));
  inv1  gate1867(.a(s_189), .O(gate86inter4));
  nand2 gate1868(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1869(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1870(.a(G8), .O(gate86inter7));
  inv1  gate1871(.a(G332), .O(gate86inter8));
  nand2 gate1872(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1873(.a(s_189), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1874(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1875(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1876(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate659(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate660(.a(gate88inter0), .b(s_16), .O(gate88inter1));
  and2  gate661(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate662(.a(s_16), .O(gate88inter3));
  inv1  gate663(.a(s_17), .O(gate88inter4));
  nand2 gate664(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate665(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate666(.a(G16), .O(gate88inter7));
  inv1  gate667(.a(G335), .O(gate88inter8));
  nand2 gate668(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate669(.a(s_17), .b(gate88inter3), .O(gate88inter10));
  nor2  gate670(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate671(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate672(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2045(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2046(.a(gate89inter0), .b(s_214), .O(gate89inter1));
  and2  gate2047(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2048(.a(s_214), .O(gate89inter3));
  inv1  gate2049(.a(s_215), .O(gate89inter4));
  nand2 gate2050(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2051(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2052(.a(G17), .O(gate89inter7));
  inv1  gate2053(.a(G338), .O(gate89inter8));
  nand2 gate2054(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2055(.a(s_215), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2056(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2057(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2058(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2101(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2102(.a(gate94inter0), .b(s_222), .O(gate94inter1));
  and2  gate2103(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2104(.a(s_222), .O(gate94inter3));
  inv1  gate2105(.a(s_223), .O(gate94inter4));
  nand2 gate2106(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2107(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2108(.a(G22), .O(gate94inter7));
  inv1  gate2109(.a(G344), .O(gate94inter8));
  nand2 gate2110(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2111(.a(s_223), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2112(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2113(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2114(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1359(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1360(.a(gate98inter0), .b(s_116), .O(gate98inter1));
  and2  gate1361(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1362(.a(s_116), .O(gate98inter3));
  inv1  gate1363(.a(s_117), .O(gate98inter4));
  nand2 gate1364(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1365(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1366(.a(G23), .O(gate98inter7));
  inv1  gate1367(.a(G350), .O(gate98inter8));
  nand2 gate1368(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1369(.a(s_117), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1370(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1371(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1372(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1261(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1262(.a(gate99inter0), .b(s_102), .O(gate99inter1));
  and2  gate1263(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1264(.a(s_102), .O(gate99inter3));
  inv1  gate1265(.a(s_103), .O(gate99inter4));
  nand2 gate1266(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1267(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1268(.a(G27), .O(gate99inter7));
  inv1  gate1269(.a(G353), .O(gate99inter8));
  nand2 gate1270(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1271(.a(s_103), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1272(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1273(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1274(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1989(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1990(.a(gate100inter0), .b(s_206), .O(gate100inter1));
  and2  gate1991(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1992(.a(s_206), .O(gate100inter3));
  inv1  gate1993(.a(s_207), .O(gate100inter4));
  nand2 gate1994(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1995(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1996(.a(G31), .O(gate100inter7));
  inv1  gate1997(.a(G353), .O(gate100inter8));
  nand2 gate1998(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1999(.a(s_207), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2000(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2001(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2002(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1933(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1934(.a(gate102inter0), .b(s_198), .O(gate102inter1));
  and2  gate1935(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1936(.a(s_198), .O(gate102inter3));
  inv1  gate1937(.a(s_199), .O(gate102inter4));
  nand2 gate1938(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1939(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1940(.a(G24), .O(gate102inter7));
  inv1  gate1941(.a(G356), .O(gate102inter8));
  nand2 gate1942(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1943(.a(s_199), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1944(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1945(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1946(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate575(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate576(.a(gate104inter0), .b(s_4), .O(gate104inter1));
  and2  gate577(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate578(.a(s_4), .O(gate104inter3));
  inv1  gate579(.a(s_5), .O(gate104inter4));
  nand2 gate580(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate581(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate582(.a(G32), .O(gate104inter7));
  inv1  gate583(.a(G359), .O(gate104inter8));
  nand2 gate584(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate585(.a(s_5), .b(gate104inter3), .O(gate104inter10));
  nor2  gate586(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate587(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate588(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1107(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1108(.a(gate107inter0), .b(s_80), .O(gate107inter1));
  and2  gate1109(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1110(.a(s_80), .O(gate107inter3));
  inv1  gate1111(.a(s_81), .O(gate107inter4));
  nand2 gate1112(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1113(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1114(.a(G366), .O(gate107inter7));
  inv1  gate1115(.a(G367), .O(gate107inter8));
  nand2 gate1116(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1117(.a(s_81), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1118(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1119(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1120(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate967(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate968(.a(gate110inter0), .b(s_60), .O(gate110inter1));
  and2  gate969(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate970(.a(s_60), .O(gate110inter3));
  inv1  gate971(.a(s_61), .O(gate110inter4));
  nand2 gate972(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate973(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate974(.a(G372), .O(gate110inter7));
  inv1  gate975(.a(G373), .O(gate110inter8));
  nand2 gate976(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate977(.a(s_61), .b(gate110inter3), .O(gate110inter10));
  nor2  gate978(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate979(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate980(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate827(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate828(.a(gate112inter0), .b(s_40), .O(gate112inter1));
  and2  gate829(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate830(.a(s_40), .O(gate112inter3));
  inv1  gate831(.a(s_41), .O(gate112inter4));
  nand2 gate832(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate833(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate834(.a(G376), .O(gate112inter7));
  inv1  gate835(.a(G377), .O(gate112inter8));
  nand2 gate836(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate837(.a(s_41), .b(gate112inter3), .O(gate112inter10));
  nor2  gate838(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate839(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate840(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1401(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1402(.a(gate115inter0), .b(s_122), .O(gate115inter1));
  and2  gate1403(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1404(.a(s_122), .O(gate115inter3));
  inv1  gate1405(.a(s_123), .O(gate115inter4));
  nand2 gate1406(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1407(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1408(.a(G382), .O(gate115inter7));
  inv1  gate1409(.a(G383), .O(gate115inter8));
  nand2 gate1410(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1411(.a(s_123), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1412(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1413(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1414(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate2199(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2200(.a(gate116inter0), .b(s_236), .O(gate116inter1));
  and2  gate2201(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2202(.a(s_236), .O(gate116inter3));
  inv1  gate2203(.a(s_237), .O(gate116inter4));
  nand2 gate2204(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2205(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2206(.a(G384), .O(gate116inter7));
  inv1  gate2207(.a(G385), .O(gate116inter8));
  nand2 gate2208(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2209(.a(s_237), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2210(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2211(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2212(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1765(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1766(.a(gate123inter0), .b(s_174), .O(gate123inter1));
  and2  gate1767(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1768(.a(s_174), .O(gate123inter3));
  inv1  gate1769(.a(s_175), .O(gate123inter4));
  nand2 gate1770(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1771(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1772(.a(G398), .O(gate123inter7));
  inv1  gate1773(.a(G399), .O(gate123inter8));
  nand2 gate1774(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1775(.a(s_175), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1776(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1777(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1778(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1457(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1458(.a(gate124inter0), .b(s_130), .O(gate124inter1));
  and2  gate1459(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1460(.a(s_130), .O(gate124inter3));
  inv1  gate1461(.a(s_131), .O(gate124inter4));
  nand2 gate1462(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1463(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1464(.a(G400), .O(gate124inter7));
  inv1  gate1465(.a(G401), .O(gate124inter8));
  nand2 gate1466(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1467(.a(s_131), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1468(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1469(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1470(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1779(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1780(.a(gate125inter0), .b(s_176), .O(gate125inter1));
  and2  gate1781(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1782(.a(s_176), .O(gate125inter3));
  inv1  gate1783(.a(s_177), .O(gate125inter4));
  nand2 gate1784(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1785(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1786(.a(G402), .O(gate125inter7));
  inv1  gate1787(.a(G403), .O(gate125inter8));
  nand2 gate1788(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1789(.a(s_177), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1790(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1791(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1792(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2451(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2452(.a(gate127inter0), .b(s_272), .O(gate127inter1));
  and2  gate2453(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2454(.a(s_272), .O(gate127inter3));
  inv1  gate2455(.a(s_273), .O(gate127inter4));
  nand2 gate2456(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2457(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2458(.a(G406), .O(gate127inter7));
  inv1  gate2459(.a(G407), .O(gate127inter8));
  nand2 gate2460(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2461(.a(s_273), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2462(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2463(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2464(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1975(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1976(.a(gate129inter0), .b(s_204), .O(gate129inter1));
  and2  gate1977(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1978(.a(s_204), .O(gate129inter3));
  inv1  gate1979(.a(s_205), .O(gate129inter4));
  nand2 gate1980(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1981(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1982(.a(G410), .O(gate129inter7));
  inv1  gate1983(.a(G411), .O(gate129inter8));
  nand2 gate1984(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1985(.a(s_205), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1986(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1987(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1988(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2129(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2130(.a(gate132inter0), .b(s_226), .O(gate132inter1));
  and2  gate2131(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2132(.a(s_226), .O(gate132inter3));
  inv1  gate2133(.a(s_227), .O(gate132inter4));
  nand2 gate2134(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2135(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2136(.a(G416), .O(gate132inter7));
  inv1  gate2137(.a(G417), .O(gate132inter8));
  nand2 gate2138(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2139(.a(s_227), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2140(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2141(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2142(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2185(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2186(.a(gate140inter0), .b(s_234), .O(gate140inter1));
  and2  gate2187(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2188(.a(s_234), .O(gate140inter3));
  inv1  gate2189(.a(s_235), .O(gate140inter4));
  nand2 gate2190(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2191(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2192(.a(G444), .O(gate140inter7));
  inv1  gate2193(.a(G447), .O(gate140inter8));
  nand2 gate2194(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2195(.a(s_235), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2196(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2197(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2198(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1079(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1080(.a(gate142inter0), .b(s_76), .O(gate142inter1));
  and2  gate1081(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1082(.a(s_76), .O(gate142inter3));
  inv1  gate1083(.a(s_77), .O(gate142inter4));
  nand2 gate1084(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1085(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1086(.a(G456), .O(gate142inter7));
  inv1  gate1087(.a(G459), .O(gate142inter8));
  nand2 gate1088(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1089(.a(s_77), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1090(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1091(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1092(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1639(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1640(.a(gate143inter0), .b(s_156), .O(gate143inter1));
  and2  gate1641(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1642(.a(s_156), .O(gate143inter3));
  inv1  gate1643(.a(s_157), .O(gate143inter4));
  nand2 gate1644(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1645(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1646(.a(G462), .O(gate143inter7));
  inv1  gate1647(.a(G465), .O(gate143inter8));
  nand2 gate1648(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1649(.a(s_157), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1650(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1651(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1652(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate981(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate982(.a(gate146inter0), .b(s_62), .O(gate146inter1));
  and2  gate983(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate984(.a(s_62), .O(gate146inter3));
  inv1  gate985(.a(s_63), .O(gate146inter4));
  nand2 gate986(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate987(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate988(.a(G480), .O(gate146inter7));
  inv1  gate989(.a(G483), .O(gate146inter8));
  nand2 gate990(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate991(.a(s_63), .b(gate146inter3), .O(gate146inter10));
  nor2  gate992(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate993(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate994(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2059(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2060(.a(gate148inter0), .b(s_216), .O(gate148inter1));
  and2  gate2061(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2062(.a(s_216), .O(gate148inter3));
  inv1  gate2063(.a(s_217), .O(gate148inter4));
  nand2 gate2064(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2065(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2066(.a(G492), .O(gate148inter7));
  inv1  gate2067(.a(G495), .O(gate148inter8));
  nand2 gate2068(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2069(.a(s_217), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2070(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2071(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2072(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1611(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1612(.a(gate150inter0), .b(s_152), .O(gate150inter1));
  and2  gate1613(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1614(.a(s_152), .O(gate150inter3));
  inv1  gate1615(.a(s_153), .O(gate150inter4));
  nand2 gate1616(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1617(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1618(.a(G504), .O(gate150inter7));
  inv1  gate1619(.a(G507), .O(gate150inter8));
  nand2 gate1620(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1621(.a(s_153), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1622(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1623(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1624(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1891(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1892(.a(gate152inter0), .b(s_192), .O(gate152inter1));
  and2  gate1893(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1894(.a(s_192), .O(gate152inter3));
  inv1  gate1895(.a(s_193), .O(gate152inter4));
  nand2 gate1896(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1897(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1898(.a(G516), .O(gate152inter7));
  inv1  gate1899(.a(G519), .O(gate152inter8));
  nand2 gate1900(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1901(.a(s_193), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1902(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1903(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1904(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2493(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2494(.a(gate154inter0), .b(s_278), .O(gate154inter1));
  and2  gate2495(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2496(.a(s_278), .O(gate154inter3));
  inv1  gate2497(.a(s_279), .O(gate154inter4));
  nand2 gate2498(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2499(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2500(.a(G429), .O(gate154inter7));
  inv1  gate2501(.a(G522), .O(gate154inter8));
  nand2 gate2502(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2503(.a(s_279), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2504(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2505(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2506(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1135(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1136(.a(gate155inter0), .b(s_84), .O(gate155inter1));
  and2  gate1137(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1138(.a(s_84), .O(gate155inter3));
  inv1  gate1139(.a(s_85), .O(gate155inter4));
  nand2 gate1140(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1141(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1142(.a(G432), .O(gate155inter7));
  inv1  gate1143(.a(G525), .O(gate155inter8));
  nand2 gate1144(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1145(.a(s_85), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1146(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1147(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1148(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2227(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2228(.a(gate156inter0), .b(s_240), .O(gate156inter1));
  and2  gate2229(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2230(.a(s_240), .O(gate156inter3));
  inv1  gate2231(.a(s_241), .O(gate156inter4));
  nand2 gate2232(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2233(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2234(.a(G435), .O(gate156inter7));
  inv1  gate2235(.a(G525), .O(gate156inter8));
  nand2 gate2236(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2237(.a(s_241), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2238(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2239(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2240(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2171(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2172(.a(gate157inter0), .b(s_232), .O(gate157inter1));
  and2  gate2173(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2174(.a(s_232), .O(gate157inter3));
  inv1  gate2175(.a(s_233), .O(gate157inter4));
  nand2 gate2176(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2177(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2178(.a(G438), .O(gate157inter7));
  inv1  gate2179(.a(G528), .O(gate157inter8));
  nand2 gate2180(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2181(.a(s_233), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2182(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2183(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2184(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2339(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2340(.a(gate161inter0), .b(s_256), .O(gate161inter1));
  and2  gate2341(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2342(.a(s_256), .O(gate161inter3));
  inv1  gate2343(.a(s_257), .O(gate161inter4));
  nand2 gate2344(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2345(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2346(.a(G450), .O(gate161inter7));
  inv1  gate2347(.a(G534), .O(gate161inter8));
  nand2 gate2348(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2349(.a(s_257), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2350(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2351(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2352(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2507(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2508(.a(gate166inter0), .b(s_280), .O(gate166inter1));
  and2  gate2509(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2510(.a(s_280), .O(gate166inter3));
  inv1  gate2511(.a(s_281), .O(gate166inter4));
  nand2 gate2512(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2513(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2514(.a(G465), .O(gate166inter7));
  inv1  gate2515(.a(G540), .O(gate166inter8));
  nand2 gate2516(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2517(.a(s_281), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2518(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2519(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2520(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate897(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate898(.a(gate167inter0), .b(s_50), .O(gate167inter1));
  and2  gate899(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate900(.a(s_50), .O(gate167inter3));
  inv1  gate901(.a(s_51), .O(gate167inter4));
  nand2 gate902(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate903(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate904(.a(G468), .O(gate167inter7));
  inv1  gate905(.a(G543), .O(gate167inter8));
  nand2 gate906(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate907(.a(s_51), .b(gate167inter3), .O(gate167inter10));
  nor2  gate908(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate909(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate910(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1317(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1318(.a(gate168inter0), .b(s_110), .O(gate168inter1));
  and2  gate1319(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1320(.a(s_110), .O(gate168inter3));
  inv1  gate1321(.a(s_111), .O(gate168inter4));
  nand2 gate1322(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1323(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1324(.a(G471), .O(gate168inter7));
  inv1  gate1325(.a(G543), .O(gate168inter8));
  nand2 gate1326(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1327(.a(s_111), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1328(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1329(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1330(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1485(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1486(.a(gate171inter0), .b(s_134), .O(gate171inter1));
  and2  gate1487(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1488(.a(s_134), .O(gate171inter3));
  inv1  gate1489(.a(s_135), .O(gate171inter4));
  nand2 gate1490(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1491(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1492(.a(G480), .O(gate171inter7));
  inv1  gate1493(.a(G549), .O(gate171inter8));
  nand2 gate1494(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1495(.a(s_135), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1496(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1497(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1498(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2479(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2480(.a(gate174inter0), .b(s_276), .O(gate174inter1));
  and2  gate2481(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2482(.a(s_276), .O(gate174inter3));
  inv1  gate2483(.a(s_277), .O(gate174inter4));
  nand2 gate2484(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2485(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2486(.a(G489), .O(gate174inter7));
  inv1  gate2487(.a(G552), .O(gate174inter8));
  nand2 gate2488(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2489(.a(s_277), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2490(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2491(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2492(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate729(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate730(.a(gate175inter0), .b(s_26), .O(gate175inter1));
  and2  gate731(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate732(.a(s_26), .O(gate175inter3));
  inv1  gate733(.a(s_27), .O(gate175inter4));
  nand2 gate734(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate735(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate736(.a(G492), .O(gate175inter7));
  inv1  gate737(.a(G555), .O(gate175inter8));
  nand2 gate738(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate739(.a(s_27), .b(gate175inter3), .O(gate175inter10));
  nor2  gate740(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate741(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate742(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1331(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1332(.a(gate178inter0), .b(s_112), .O(gate178inter1));
  and2  gate1333(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1334(.a(s_112), .O(gate178inter3));
  inv1  gate1335(.a(s_113), .O(gate178inter4));
  nand2 gate1336(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1337(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1338(.a(G501), .O(gate178inter7));
  inv1  gate1339(.a(G558), .O(gate178inter8));
  nand2 gate1340(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1341(.a(s_113), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1342(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1343(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1344(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate1625(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1626(.a(gate179inter0), .b(s_154), .O(gate179inter1));
  and2  gate1627(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1628(.a(s_154), .O(gate179inter3));
  inv1  gate1629(.a(s_155), .O(gate179inter4));
  nand2 gate1630(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1631(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1632(.a(G504), .O(gate179inter7));
  inv1  gate1633(.a(G561), .O(gate179inter8));
  nand2 gate1634(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1635(.a(s_155), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1636(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1637(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1638(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1877(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1878(.a(gate180inter0), .b(s_190), .O(gate180inter1));
  and2  gate1879(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1880(.a(s_190), .O(gate180inter3));
  inv1  gate1881(.a(s_191), .O(gate180inter4));
  nand2 gate1882(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1883(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1884(.a(G507), .O(gate180inter7));
  inv1  gate1885(.a(G561), .O(gate180inter8));
  nand2 gate1886(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1887(.a(s_191), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1888(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1889(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1890(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1583(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1584(.a(gate183inter0), .b(s_148), .O(gate183inter1));
  and2  gate1585(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1586(.a(s_148), .O(gate183inter3));
  inv1  gate1587(.a(s_149), .O(gate183inter4));
  nand2 gate1588(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1589(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1590(.a(G516), .O(gate183inter7));
  inv1  gate1591(.a(G567), .O(gate183inter8));
  nand2 gate1592(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1593(.a(s_149), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1594(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1595(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1596(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate603(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate604(.a(gate184inter0), .b(s_8), .O(gate184inter1));
  and2  gate605(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate606(.a(s_8), .O(gate184inter3));
  inv1  gate607(.a(s_9), .O(gate184inter4));
  nand2 gate608(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate609(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate610(.a(G519), .O(gate184inter7));
  inv1  gate611(.a(G567), .O(gate184inter8));
  nand2 gate612(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate613(.a(s_9), .b(gate184inter3), .O(gate184inter10));
  nor2  gate614(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate615(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate616(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1849(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1850(.a(gate190inter0), .b(s_186), .O(gate190inter1));
  and2  gate1851(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1852(.a(s_186), .O(gate190inter3));
  inv1  gate1853(.a(s_187), .O(gate190inter4));
  nand2 gate1854(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1855(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1856(.a(G580), .O(gate190inter7));
  inv1  gate1857(.a(G581), .O(gate190inter8));
  nand2 gate1858(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1859(.a(s_187), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1860(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1861(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1862(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1191(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1192(.a(gate194inter0), .b(s_92), .O(gate194inter1));
  and2  gate1193(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1194(.a(s_92), .O(gate194inter3));
  inv1  gate1195(.a(s_93), .O(gate194inter4));
  nand2 gate1196(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1197(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1198(.a(G588), .O(gate194inter7));
  inv1  gate1199(.a(G589), .O(gate194inter8));
  nand2 gate1200(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1201(.a(s_93), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1202(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1203(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1204(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1653(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1654(.a(gate202inter0), .b(s_158), .O(gate202inter1));
  and2  gate1655(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1656(.a(s_158), .O(gate202inter3));
  inv1  gate1657(.a(s_159), .O(gate202inter4));
  nand2 gate1658(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1659(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1660(.a(G612), .O(gate202inter7));
  inv1  gate1661(.a(G617), .O(gate202inter8));
  nand2 gate1662(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1663(.a(s_159), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1664(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1665(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1666(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1205(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1206(.a(gate203inter0), .b(s_94), .O(gate203inter1));
  and2  gate1207(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1208(.a(s_94), .O(gate203inter3));
  inv1  gate1209(.a(s_95), .O(gate203inter4));
  nand2 gate1210(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1211(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1212(.a(G602), .O(gate203inter7));
  inv1  gate1213(.a(G612), .O(gate203inter8));
  nand2 gate1214(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1215(.a(s_95), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1216(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1217(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1218(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate715(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate716(.a(gate205inter0), .b(s_24), .O(gate205inter1));
  and2  gate717(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate718(.a(s_24), .O(gate205inter3));
  inv1  gate719(.a(s_25), .O(gate205inter4));
  nand2 gate720(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate721(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate722(.a(G622), .O(gate205inter7));
  inv1  gate723(.a(G627), .O(gate205inter8));
  nand2 gate724(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate725(.a(s_25), .b(gate205inter3), .O(gate205inter10));
  nor2  gate726(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate727(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate728(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2073(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2074(.a(gate206inter0), .b(s_218), .O(gate206inter1));
  and2  gate2075(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2076(.a(s_218), .O(gate206inter3));
  inv1  gate2077(.a(s_219), .O(gate206inter4));
  nand2 gate2078(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2079(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2080(.a(G632), .O(gate206inter7));
  inv1  gate2081(.a(G637), .O(gate206inter8));
  nand2 gate2082(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2083(.a(s_219), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2084(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2085(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2086(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate687(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate688(.a(gate208inter0), .b(s_20), .O(gate208inter1));
  and2  gate689(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate690(.a(s_20), .O(gate208inter3));
  inv1  gate691(.a(s_21), .O(gate208inter4));
  nand2 gate692(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate693(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate694(.a(G627), .O(gate208inter7));
  inv1  gate695(.a(G637), .O(gate208inter8));
  nand2 gate696(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate697(.a(s_21), .b(gate208inter3), .O(gate208inter10));
  nor2  gate698(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate699(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate700(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1793(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1794(.a(gate213inter0), .b(s_178), .O(gate213inter1));
  and2  gate1795(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1796(.a(s_178), .O(gate213inter3));
  inv1  gate1797(.a(s_179), .O(gate213inter4));
  nand2 gate1798(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1799(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1800(.a(G602), .O(gate213inter7));
  inv1  gate1801(.a(G672), .O(gate213inter8));
  nand2 gate1802(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1803(.a(s_179), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1804(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1805(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1806(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1667(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1668(.a(gate214inter0), .b(s_160), .O(gate214inter1));
  and2  gate1669(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1670(.a(s_160), .O(gate214inter3));
  inv1  gate1671(.a(s_161), .O(gate214inter4));
  nand2 gate1672(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1673(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1674(.a(G612), .O(gate214inter7));
  inv1  gate1675(.a(G672), .O(gate214inter8));
  nand2 gate1676(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1677(.a(s_161), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1678(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1679(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1680(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate673(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate674(.a(gate218inter0), .b(s_18), .O(gate218inter1));
  and2  gate675(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate676(.a(s_18), .O(gate218inter3));
  inv1  gate677(.a(s_19), .O(gate218inter4));
  nand2 gate678(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate679(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate680(.a(G627), .O(gate218inter7));
  inv1  gate681(.a(G678), .O(gate218inter8));
  nand2 gate682(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate683(.a(s_19), .b(gate218inter3), .O(gate218inter10));
  nor2  gate684(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate685(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate686(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate631(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate632(.a(gate221inter0), .b(s_12), .O(gate221inter1));
  and2  gate633(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate634(.a(s_12), .O(gate221inter3));
  inv1  gate635(.a(s_13), .O(gate221inter4));
  nand2 gate636(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate637(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate638(.a(G622), .O(gate221inter7));
  inv1  gate639(.a(G684), .O(gate221inter8));
  nand2 gate640(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate641(.a(s_13), .b(gate221inter3), .O(gate221inter10));
  nor2  gate642(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate643(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate644(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1555(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1556(.a(gate224inter0), .b(s_144), .O(gate224inter1));
  and2  gate1557(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1558(.a(s_144), .O(gate224inter3));
  inv1  gate1559(.a(s_145), .O(gate224inter4));
  nand2 gate1560(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1561(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1562(.a(G637), .O(gate224inter7));
  inv1  gate1563(.a(G687), .O(gate224inter8));
  nand2 gate1564(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1565(.a(s_145), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1566(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1567(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1568(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1751(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1752(.a(gate228inter0), .b(s_172), .O(gate228inter1));
  and2  gate1753(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1754(.a(s_172), .O(gate228inter3));
  inv1  gate1755(.a(s_173), .O(gate228inter4));
  nand2 gate1756(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1757(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1758(.a(G696), .O(gate228inter7));
  inv1  gate1759(.a(G697), .O(gate228inter8));
  nand2 gate1760(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1761(.a(s_173), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1762(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1763(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1764(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1149(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1150(.a(gate229inter0), .b(s_86), .O(gate229inter1));
  and2  gate1151(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1152(.a(s_86), .O(gate229inter3));
  inv1  gate1153(.a(s_87), .O(gate229inter4));
  nand2 gate1154(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1155(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1156(.a(G698), .O(gate229inter7));
  inv1  gate1157(.a(G699), .O(gate229inter8));
  nand2 gate1158(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1159(.a(s_87), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1160(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1161(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1162(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1681(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1682(.a(gate235inter0), .b(s_162), .O(gate235inter1));
  and2  gate1683(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1684(.a(s_162), .O(gate235inter3));
  inv1  gate1685(.a(s_163), .O(gate235inter4));
  nand2 gate1686(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1687(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1688(.a(G248), .O(gate235inter7));
  inv1  gate1689(.a(G724), .O(gate235inter8));
  nand2 gate1690(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1691(.a(s_163), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1692(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1693(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1694(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1387(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1388(.a(gate240inter0), .b(s_120), .O(gate240inter1));
  and2  gate1389(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1390(.a(s_120), .O(gate240inter3));
  inv1  gate1391(.a(s_121), .O(gate240inter4));
  nand2 gate1392(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1393(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1394(.a(G263), .O(gate240inter7));
  inv1  gate1395(.a(G715), .O(gate240inter8));
  nand2 gate1396(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1397(.a(s_121), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1398(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1399(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1400(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2003(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2004(.a(gate244inter0), .b(s_208), .O(gate244inter1));
  and2  gate2005(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2006(.a(s_208), .O(gate244inter3));
  inv1  gate2007(.a(s_209), .O(gate244inter4));
  nand2 gate2008(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2009(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2010(.a(G721), .O(gate244inter7));
  inv1  gate2011(.a(G733), .O(gate244inter8));
  nand2 gate2012(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2013(.a(s_209), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2014(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2015(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2016(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1415(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1416(.a(gate248inter0), .b(s_124), .O(gate248inter1));
  and2  gate1417(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1418(.a(s_124), .O(gate248inter3));
  inv1  gate1419(.a(s_125), .O(gate248inter4));
  nand2 gate1420(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1421(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1422(.a(G727), .O(gate248inter7));
  inv1  gate1423(.a(G739), .O(gate248inter8));
  nand2 gate1424(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1425(.a(s_125), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1426(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1427(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1428(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate547(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate548(.a(gate250inter0), .b(s_0), .O(gate250inter1));
  and2  gate549(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate550(.a(s_0), .O(gate250inter3));
  inv1  gate551(.a(s_1), .O(gate250inter4));
  nand2 gate552(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate553(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate554(.a(G706), .O(gate250inter7));
  inv1  gate555(.a(G742), .O(gate250inter8));
  nand2 gate556(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate557(.a(s_1), .b(gate250inter3), .O(gate250inter10));
  nor2  gate558(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate559(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate560(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2143(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2144(.a(gate253inter0), .b(s_228), .O(gate253inter1));
  and2  gate2145(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2146(.a(s_228), .O(gate253inter3));
  inv1  gate2147(.a(s_229), .O(gate253inter4));
  nand2 gate2148(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2149(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2150(.a(G260), .O(gate253inter7));
  inv1  gate2151(.a(G748), .O(gate253inter8));
  nand2 gate2152(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2153(.a(s_229), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2154(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2155(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2156(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1177(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1178(.a(gate255inter0), .b(s_90), .O(gate255inter1));
  and2  gate1179(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1180(.a(s_90), .O(gate255inter3));
  inv1  gate1181(.a(s_91), .O(gate255inter4));
  nand2 gate1182(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1183(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1184(.a(G263), .O(gate255inter7));
  inv1  gate1185(.a(G751), .O(gate255inter8));
  nand2 gate1186(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1187(.a(s_91), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1188(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1189(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1190(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate2283(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2284(.a(gate256inter0), .b(s_248), .O(gate256inter1));
  and2  gate2285(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2286(.a(s_248), .O(gate256inter3));
  inv1  gate2287(.a(s_249), .O(gate256inter4));
  nand2 gate2288(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2289(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2290(.a(G715), .O(gate256inter7));
  inv1  gate2291(.a(G751), .O(gate256inter8));
  nand2 gate2292(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2293(.a(s_249), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2294(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2295(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2296(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate995(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate996(.a(gate261inter0), .b(s_64), .O(gate261inter1));
  and2  gate997(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate998(.a(s_64), .O(gate261inter3));
  inv1  gate999(.a(s_65), .O(gate261inter4));
  nand2 gate1000(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1001(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1002(.a(G762), .O(gate261inter7));
  inv1  gate1003(.a(G763), .O(gate261inter8));
  nand2 gate1004(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1005(.a(s_65), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1006(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1007(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1008(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate953(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate954(.a(gate262inter0), .b(s_58), .O(gate262inter1));
  and2  gate955(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate956(.a(s_58), .O(gate262inter3));
  inv1  gate957(.a(s_59), .O(gate262inter4));
  nand2 gate958(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate959(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate960(.a(G764), .O(gate262inter7));
  inv1  gate961(.a(G765), .O(gate262inter8));
  nand2 gate962(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate963(.a(s_59), .b(gate262inter3), .O(gate262inter10));
  nor2  gate964(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate965(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate966(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1499(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1500(.a(gate265inter0), .b(s_136), .O(gate265inter1));
  and2  gate1501(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1502(.a(s_136), .O(gate265inter3));
  inv1  gate1503(.a(s_137), .O(gate265inter4));
  nand2 gate1504(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1505(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1506(.a(G642), .O(gate265inter7));
  inv1  gate1507(.a(G770), .O(gate265inter8));
  nand2 gate1508(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1509(.a(s_137), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1510(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1511(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1512(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1275(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1276(.a(gate278inter0), .b(s_104), .O(gate278inter1));
  and2  gate1277(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1278(.a(s_104), .O(gate278inter3));
  inv1  gate1279(.a(s_105), .O(gate278inter4));
  nand2 gate1280(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1281(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1282(.a(G776), .O(gate278inter7));
  inv1  gate1283(.a(G800), .O(gate278inter8));
  nand2 gate1284(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1285(.a(s_105), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1286(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1287(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1288(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1429(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1430(.a(gate280inter0), .b(s_126), .O(gate280inter1));
  and2  gate1431(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1432(.a(s_126), .O(gate280inter3));
  inv1  gate1433(.a(s_127), .O(gate280inter4));
  nand2 gate1434(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1435(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1436(.a(G779), .O(gate280inter7));
  inv1  gate1437(.a(G803), .O(gate280inter8));
  nand2 gate1438(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1439(.a(s_127), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1440(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1441(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1442(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1037(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1038(.a(gate281inter0), .b(s_70), .O(gate281inter1));
  and2  gate1039(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1040(.a(s_70), .O(gate281inter3));
  inv1  gate1041(.a(s_71), .O(gate281inter4));
  nand2 gate1042(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1043(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1044(.a(G654), .O(gate281inter7));
  inv1  gate1045(.a(G806), .O(gate281inter8));
  nand2 gate1046(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1047(.a(s_71), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1048(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1049(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1050(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2437(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2438(.a(gate287inter0), .b(s_270), .O(gate287inter1));
  and2  gate2439(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2440(.a(s_270), .O(gate287inter3));
  inv1  gate2441(.a(s_271), .O(gate287inter4));
  nand2 gate2442(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2443(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2444(.a(G663), .O(gate287inter7));
  inv1  gate2445(.a(G815), .O(gate287inter8));
  nand2 gate2446(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2447(.a(s_271), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2448(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2449(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2450(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1737(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1738(.a(gate288inter0), .b(s_170), .O(gate288inter1));
  and2  gate1739(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1740(.a(s_170), .O(gate288inter3));
  inv1  gate1741(.a(s_171), .O(gate288inter4));
  nand2 gate1742(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1743(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1744(.a(G791), .O(gate288inter7));
  inv1  gate1745(.a(G815), .O(gate288inter8));
  nand2 gate1746(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1747(.a(s_171), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1748(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1749(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1750(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2409(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2410(.a(gate293inter0), .b(s_266), .O(gate293inter1));
  and2  gate2411(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2412(.a(s_266), .O(gate293inter3));
  inv1  gate2413(.a(s_267), .O(gate293inter4));
  nand2 gate2414(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2415(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2416(.a(G828), .O(gate293inter7));
  inv1  gate2417(.a(G829), .O(gate293inter8));
  nand2 gate2418(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2419(.a(s_267), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2420(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2421(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2422(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1709(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1710(.a(gate294inter0), .b(s_166), .O(gate294inter1));
  and2  gate1711(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1712(.a(s_166), .O(gate294inter3));
  inv1  gate1713(.a(s_167), .O(gate294inter4));
  nand2 gate1714(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1715(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1716(.a(G832), .O(gate294inter7));
  inv1  gate1717(.a(G833), .O(gate294inter8));
  nand2 gate1718(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1719(.a(s_167), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1720(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1721(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1722(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2115(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2116(.a(gate387inter0), .b(s_224), .O(gate387inter1));
  and2  gate2117(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2118(.a(s_224), .O(gate387inter3));
  inv1  gate2119(.a(s_225), .O(gate387inter4));
  nand2 gate2120(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2121(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2122(.a(G1), .O(gate387inter7));
  inv1  gate2123(.a(G1036), .O(gate387inter8));
  nand2 gate2124(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2125(.a(s_225), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2126(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2127(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2128(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1219(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1220(.a(gate389inter0), .b(s_96), .O(gate389inter1));
  and2  gate1221(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1222(.a(s_96), .O(gate389inter3));
  inv1  gate1223(.a(s_97), .O(gate389inter4));
  nand2 gate1224(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1225(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1226(.a(G3), .O(gate389inter7));
  inv1  gate1227(.a(G1042), .O(gate389inter8));
  nand2 gate1228(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1229(.a(s_97), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1230(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1231(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1232(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate2017(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2018(.a(gate390inter0), .b(s_210), .O(gate390inter1));
  and2  gate2019(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2020(.a(s_210), .O(gate390inter3));
  inv1  gate2021(.a(s_211), .O(gate390inter4));
  nand2 gate2022(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2023(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2024(.a(G4), .O(gate390inter7));
  inv1  gate2025(.a(G1045), .O(gate390inter8));
  nand2 gate2026(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2027(.a(s_211), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2028(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2029(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2030(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1723(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1724(.a(gate394inter0), .b(s_168), .O(gate394inter1));
  and2  gate1725(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1726(.a(s_168), .O(gate394inter3));
  inv1  gate1727(.a(s_169), .O(gate394inter4));
  nand2 gate1728(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1729(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1730(.a(G8), .O(gate394inter7));
  inv1  gate1731(.a(G1057), .O(gate394inter8));
  nand2 gate1732(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1733(.a(s_169), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1734(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1735(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1736(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate2311(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2312(.a(gate399inter0), .b(s_252), .O(gate399inter1));
  and2  gate2313(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2314(.a(s_252), .O(gate399inter3));
  inv1  gate2315(.a(s_253), .O(gate399inter4));
  nand2 gate2316(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2317(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2318(.a(G13), .O(gate399inter7));
  inv1  gate2319(.a(G1072), .O(gate399inter8));
  nand2 gate2320(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2321(.a(s_253), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2322(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2323(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2324(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1835(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1836(.a(gate403inter0), .b(s_184), .O(gate403inter1));
  and2  gate1837(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1838(.a(s_184), .O(gate403inter3));
  inv1  gate1839(.a(s_185), .O(gate403inter4));
  nand2 gate1840(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1841(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1842(.a(G17), .O(gate403inter7));
  inv1  gate1843(.a(G1084), .O(gate403inter8));
  nand2 gate1844(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1845(.a(s_185), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1846(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1847(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1848(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate869(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate870(.a(gate411inter0), .b(s_46), .O(gate411inter1));
  and2  gate871(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate872(.a(s_46), .O(gate411inter3));
  inv1  gate873(.a(s_47), .O(gate411inter4));
  nand2 gate874(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate875(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate876(.a(G25), .O(gate411inter7));
  inv1  gate877(.a(G1108), .O(gate411inter8));
  nand2 gate878(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate879(.a(s_47), .b(gate411inter3), .O(gate411inter10));
  nor2  gate880(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate881(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate882(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2297(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2298(.a(gate412inter0), .b(s_250), .O(gate412inter1));
  and2  gate2299(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2300(.a(s_250), .O(gate412inter3));
  inv1  gate2301(.a(s_251), .O(gate412inter4));
  nand2 gate2302(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2303(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2304(.a(G26), .O(gate412inter7));
  inv1  gate2305(.a(G1111), .O(gate412inter8));
  nand2 gate2306(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2307(.a(s_251), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2308(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2309(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2310(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1289(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1290(.a(gate415inter0), .b(s_106), .O(gate415inter1));
  and2  gate1291(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1292(.a(s_106), .O(gate415inter3));
  inv1  gate1293(.a(s_107), .O(gate415inter4));
  nand2 gate1294(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1295(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1296(.a(G29), .O(gate415inter7));
  inv1  gate1297(.a(G1120), .O(gate415inter8));
  nand2 gate1298(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1299(.a(s_107), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1300(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1301(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1302(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2255(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2256(.a(gate417inter0), .b(s_244), .O(gate417inter1));
  and2  gate2257(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2258(.a(s_244), .O(gate417inter3));
  inv1  gate2259(.a(s_245), .O(gate417inter4));
  nand2 gate2260(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2261(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2262(.a(G31), .O(gate417inter7));
  inv1  gate2263(.a(G1126), .O(gate417inter8));
  nand2 gate2264(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2265(.a(s_245), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2266(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2267(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2268(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2465(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2466(.a(gate419inter0), .b(s_274), .O(gate419inter1));
  and2  gate2467(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2468(.a(s_274), .O(gate419inter3));
  inv1  gate2469(.a(s_275), .O(gate419inter4));
  nand2 gate2470(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2471(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2472(.a(G1), .O(gate419inter7));
  inv1  gate2473(.a(G1132), .O(gate419inter8));
  nand2 gate2474(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2475(.a(s_275), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2476(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2477(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2478(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2213(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2214(.a(gate423inter0), .b(s_238), .O(gate423inter1));
  and2  gate2215(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2216(.a(s_238), .O(gate423inter3));
  inv1  gate2217(.a(s_239), .O(gate423inter4));
  nand2 gate2218(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2219(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2220(.a(G3), .O(gate423inter7));
  inv1  gate2221(.a(G1138), .O(gate423inter8));
  nand2 gate2222(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2223(.a(s_239), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2224(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2225(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2226(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2325(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2326(.a(gate425inter0), .b(s_254), .O(gate425inter1));
  and2  gate2327(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2328(.a(s_254), .O(gate425inter3));
  inv1  gate2329(.a(s_255), .O(gate425inter4));
  nand2 gate2330(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2331(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2332(.a(G4), .O(gate425inter7));
  inv1  gate2333(.a(G1141), .O(gate425inter8));
  nand2 gate2334(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2335(.a(s_255), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2336(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2337(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2338(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1093(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1094(.a(gate427inter0), .b(s_78), .O(gate427inter1));
  and2  gate1095(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1096(.a(s_78), .O(gate427inter3));
  inv1  gate1097(.a(s_79), .O(gate427inter4));
  nand2 gate1098(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1099(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1100(.a(G5), .O(gate427inter7));
  inv1  gate1101(.a(G1144), .O(gate427inter8));
  nand2 gate1102(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1103(.a(s_79), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1104(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1105(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1106(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1905(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1906(.a(gate428inter0), .b(s_194), .O(gate428inter1));
  and2  gate1907(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1908(.a(s_194), .O(gate428inter3));
  inv1  gate1909(.a(s_195), .O(gate428inter4));
  nand2 gate1910(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1911(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1912(.a(G1048), .O(gate428inter7));
  inv1  gate1913(.a(G1144), .O(gate428inter8));
  nand2 gate1914(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1915(.a(s_195), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1916(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1917(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1918(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate855(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate856(.a(gate430inter0), .b(s_44), .O(gate430inter1));
  and2  gate857(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate858(.a(s_44), .O(gate430inter3));
  inv1  gate859(.a(s_45), .O(gate430inter4));
  nand2 gate860(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate861(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate862(.a(G1051), .O(gate430inter7));
  inv1  gate863(.a(G1147), .O(gate430inter8));
  nand2 gate864(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate865(.a(s_45), .b(gate430inter3), .O(gate430inter10));
  nor2  gate866(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate867(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate868(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate617(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate618(.a(gate436inter0), .b(s_10), .O(gate436inter1));
  and2  gate619(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate620(.a(s_10), .O(gate436inter3));
  inv1  gate621(.a(s_11), .O(gate436inter4));
  nand2 gate622(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate623(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate624(.a(G1060), .O(gate436inter7));
  inv1  gate625(.a(G1156), .O(gate436inter8));
  nand2 gate626(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate627(.a(s_11), .b(gate436inter3), .O(gate436inter10));
  nor2  gate628(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate629(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate630(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1807(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1808(.a(gate439inter0), .b(s_180), .O(gate439inter1));
  and2  gate1809(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1810(.a(s_180), .O(gate439inter3));
  inv1  gate1811(.a(s_181), .O(gate439inter4));
  nand2 gate1812(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1813(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1814(.a(G11), .O(gate439inter7));
  inv1  gate1815(.a(G1162), .O(gate439inter8));
  nand2 gate1816(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1817(.a(s_181), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1818(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1819(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1820(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate813(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate814(.a(gate440inter0), .b(s_38), .O(gate440inter1));
  and2  gate815(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate816(.a(s_38), .O(gate440inter3));
  inv1  gate817(.a(s_39), .O(gate440inter4));
  nand2 gate818(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate819(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate820(.a(G1066), .O(gate440inter7));
  inv1  gate821(.a(G1162), .O(gate440inter8));
  nand2 gate822(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate823(.a(s_39), .b(gate440inter3), .O(gate440inter10));
  nor2  gate824(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate825(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate826(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2381(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2382(.a(gate442inter0), .b(s_262), .O(gate442inter1));
  and2  gate2383(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2384(.a(s_262), .O(gate442inter3));
  inv1  gate2385(.a(s_263), .O(gate442inter4));
  nand2 gate2386(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2387(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2388(.a(G1069), .O(gate442inter7));
  inv1  gate2389(.a(G1165), .O(gate442inter8));
  nand2 gate2390(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2391(.a(s_263), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2392(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2393(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2394(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate701(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate702(.a(gate445inter0), .b(s_22), .O(gate445inter1));
  and2  gate703(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate704(.a(s_22), .O(gate445inter3));
  inv1  gate705(.a(s_23), .O(gate445inter4));
  nand2 gate706(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate707(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate708(.a(G14), .O(gate445inter7));
  inv1  gate709(.a(G1171), .O(gate445inter8));
  nand2 gate710(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate711(.a(s_23), .b(gate445inter3), .O(gate445inter10));
  nor2  gate712(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate713(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate714(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1233(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1234(.a(gate446inter0), .b(s_98), .O(gate446inter1));
  and2  gate1235(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1236(.a(s_98), .O(gate446inter3));
  inv1  gate1237(.a(s_99), .O(gate446inter4));
  nand2 gate1238(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1239(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1240(.a(G1075), .O(gate446inter7));
  inv1  gate1241(.a(G1171), .O(gate446inter8));
  nand2 gate1242(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1243(.a(s_99), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1244(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1245(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1246(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2353(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2354(.a(gate448inter0), .b(s_258), .O(gate448inter1));
  and2  gate2355(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2356(.a(s_258), .O(gate448inter3));
  inv1  gate2357(.a(s_259), .O(gate448inter4));
  nand2 gate2358(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2359(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2360(.a(G1078), .O(gate448inter7));
  inv1  gate2361(.a(G1174), .O(gate448inter8));
  nand2 gate2362(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2363(.a(s_259), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2364(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2365(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2366(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1961(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1962(.a(gate449inter0), .b(s_202), .O(gate449inter1));
  and2  gate1963(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1964(.a(s_202), .O(gate449inter3));
  inv1  gate1965(.a(s_203), .O(gate449inter4));
  nand2 gate1966(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1967(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1968(.a(G16), .O(gate449inter7));
  inv1  gate1969(.a(G1177), .O(gate449inter8));
  nand2 gate1970(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1971(.a(s_203), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1972(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1973(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1974(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2157(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2158(.a(gate457inter0), .b(s_230), .O(gate457inter1));
  and2  gate2159(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2160(.a(s_230), .O(gate457inter3));
  inv1  gate2161(.a(s_231), .O(gate457inter4));
  nand2 gate2162(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2163(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2164(.a(G20), .O(gate457inter7));
  inv1  gate2165(.a(G1189), .O(gate457inter8));
  nand2 gate2166(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2167(.a(s_231), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2168(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2169(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2170(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate561(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate562(.a(gate460inter0), .b(s_2), .O(gate460inter1));
  and2  gate563(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate564(.a(s_2), .O(gate460inter3));
  inv1  gate565(.a(s_3), .O(gate460inter4));
  nand2 gate566(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate567(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate568(.a(G1096), .O(gate460inter7));
  inv1  gate569(.a(G1192), .O(gate460inter8));
  nand2 gate570(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate571(.a(s_3), .b(gate460inter3), .O(gate460inter10));
  nor2  gate572(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate573(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate574(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1051(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1052(.a(gate469inter0), .b(s_72), .O(gate469inter1));
  and2  gate1053(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1054(.a(s_72), .O(gate469inter3));
  inv1  gate1055(.a(s_73), .O(gate469inter4));
  nand2 gate1056(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1057(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1058(.a(G26), .O(gate469inter7));
  inv1  gate1059(.a(G1207), .O(gate469inter8));
  nand2 gate1060(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1061(.a(s_73), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1062(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1063(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1064(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2367(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2368(.a(gate470inter0), .b(s_260), .O(gate470inter1));
  and2  gate2369(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2370(.a(s_260), .O(gate470inter3));
  inv1  gate2371(.a(s_261), .O(gate470inter4));
  nand2 gate2372(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2373(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2374(.a(G1111), .O(gate470inter7));
  inv1  gate2375(.a(G1207), .O(gate470inter8));
  nand2 gate2376(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2377(.a(s_261), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2378(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2379(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2380(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2269(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2270(.a(gate471inter0), .b(s_246), .O(gate471inter1));
  and2  gate2271(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2272(.a(s_246), .O(gate471inter3));
  inv1  gate2273(.a(s_247), .O(gate471inter4));
  nand2 gate2274(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2275(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2276(.a(G27), .O(gate471inter7));
  inv1  gate2277(.a(G1210), .O(gate471inter8));
  nand2 gate2278(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2279(.a(s_247), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2280(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2281(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2282(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate841(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate842(.a(gate472inter0), .b(s_42), .O(gate472inter1));
  and2  gate843(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate844(.a(s_42), .O(gate472inter3));
  inv1  gate845(.a(s_43), .O(gate472inter4));
  nand2 gate846(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate847(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate848(.a(G1114), .O(gate472inter7));
  inv1  gate849(.a(G1210), .O(gate472inter8));
  nand2 gate850(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate851(.a(s_43), .b(gate472inter3), .O(gate472inter10));
  nor2  gate852(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate853(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate854(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1163(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1164(.a(gate474inter0), .b(s_88), .O(gate474inter1));
  and2  gate1165(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1166(.a(s_88), .O(gate474inter3));
  inv1  gate1167(.a(s_89), .O(gate474inter4));
  nand2 gate1168(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1169(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1170(.a(G1117), .O(gate474inter7));
  inv1  gate1171(.a(G1213), .O(gate474inter8));
  nand2 gate1172(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1173(.a(s_89), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1174(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1175(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1176(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate939(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate940(.a(gate480inter0), .b(s_56), .O(gate480inter1));
  and2  gate941(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate942(.a(s_56), .O(gate480inter3));
  inv1  gate943(.a(s_57), .O(gate480inter4));
  nand2 gate944(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate945(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate946(.a(G1126), .O(gate480inter7));
  inv1  gate947(.a(G1222), .O(gate480inter8));
  nand2 gate948(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate949(.a(s_57), .b(gate480inter3), .O(gate480inter10));
  nor2  gate950(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate951(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate952(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate589(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate590(.a(gate483inter0), .b(s_6), .O(gate483inter1));
  and2  gate591(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate592(.a(s_6), .O(gate483inter3));
  inv1  gate593(.a(s_7), .O(gate483inter4));
  nand2 gate594(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate595(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate596(.a(G1228), .O(gate483inter7));
  inv1  gate597(.a(G1229), .O(gate483inter8));
  nand2 gate598(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate599(.a(s_7), .b(gate483inter3), .O(gate483inter10));
  nor2  gate600(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate601(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate602(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1597(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1598(.a(gate488inter0), .b(s_150), .O(gate488inter1));
  and2  gate1599(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1600(.a(s_150), .O(gate488inter3));
  inv1  gate1601(.a(s_151), .O(gate488inter4));
  nand2 gate1602(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1603(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1604(.a(G1238), .O(gate488inter7));
  inv1  gate1605(.a(G1239), .O(gate488inter8));
  nand2 gate1606(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1607(.a(s_151), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1608(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1609(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1610(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1569(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1570(.a(gate494inter0), .b(s_146), .O(gate494inter1));
  and2  gate1571(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1572(.a(s_146), .O(gate494inter3));
  inv1  gate1573(.a(s_147), .O(gate494inter4));
  nand2 gate1574(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1575(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1576(.a(G1250), .O(gate494inter7));
  inv1  gate1577(.a(G1251), .O(gate494inter8));
  nand2 gate1578(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1579(.a(s_147), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1580(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1581(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1582(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1527(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1528(.a(gate497inter0), .b(s_140), .O(gate497inter1));
  and2  gate1529(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1530(.a(s_140), .O(gate497inter3));
  inv1  gate1531(.a(s_141), .O(gate497inter4));
  nand2 gate1532(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1533(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1534(.a(G1256), .O(gate497inter7));
  inv1  gate1535(.a(G1257), .O(gate497inter8));
  nand2 gate1536(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1537(.a(s_141), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1538(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1539(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1540(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate799(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate800(.a(gate499inter0), .b(s_36), .O(gate499inter1));
  and2  gate801(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate802(.a(s_36), .O(gate499inter3));
  inv1  gate803(.a(s_37), .O(gate499inter4));
  nand2 gate804(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate805(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate806(.a(G1260), .O(gate499inter7));
  inv1  gate807(.a(G1261), .O(gate499inter8));
  nand2 gate808(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate809(.a(s_37), .b(gate499inter3), .O(gate499inter10));
  nor2  gate810(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate811(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate812(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2423(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2424(.a(gate500inter0), .b(s_268), .O(gate500inter1));
  and2  gate2425(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2426(.a(s_268), .O(gate500inter3));
  inv1  gate2427(.a(s_269), .O(gate500inter4));
  nand2 gate2428(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2429(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2430(.a(G1262), .O(gate500inter7));
  inv1  gate2431(.a(G1263), .O(gate500inter8));
  nand2 gate2432(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2433(.a(s_269), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2434(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2435(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2436(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1947(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1948(.a(gate501inter0), .b(s_200), .O(gate501inter1));
  and2  gate1949(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1950(.a(s_200), .O(gate501inter3));
  inv1  gate1951(.a(s_201), .O(gate501inter4));
  nand2 gate1952(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1953(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1954(.a(G1264), .O(gate501inter7));
  inv1  gate1955(.a(G1265), .O(gate501inter8));
  nand2 gate1956(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1957(.a(s_201), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1958(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1959(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1960(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate883(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate884(.a(gate507inter0), .b(s_48), .O(gate507inter1));
  and2  gate885(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate886(.a(s_48), .O(gate507inter3));
  inv1  gate887(.a(s_49), .O(gate507inter4));
  nand2 gate888(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate889(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate890(.a(G1276), .O(gate507inter7));
  inv1  gate891(.a(G1277), .O(gate507inter8));
  nand2 gate892(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate893(.a(s_49), .b(gate507inter3), .O(gate507inter10));
  nor2  gate894(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate895(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate896(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1821(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1822(.a(gate508inter0), .b(s_182), .O(gate508inter1));
  and2  gate1823(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1824(.a(s_182), .O(gate508inter3));
  inv1  gate1825(.a(s_183), .O(gate508inter4));
  nand2 gate1826(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1827(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1828(.a(G1278), .O(gate508inter7));
  inv1  gate1829(.a(G1279), .O(gate508inter8));
  nand2 gate1830(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1831(.a(s_183), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1832(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1833(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1834(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1695(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1696(.a(gate512inter0), .b(s_164), .O(gate512inter1));
  and2  gate1697(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1698(.a(s_164), .O(gate512inter3));
  inv1  gate1699(.a(s_165), .O(gate512inter4));
  nand2 gate1700(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1701(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1702(.a(G1286), .O(gate512inter7));
  inv1  gate1703(.a(G1287), .O(gate512inter8));
  nand2 gate1704(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1705(.a(s_165), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1706(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1707(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1708(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1345(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1346(.a(gate514inter0), .b(s_114), .O(gate514inter1));
  and2  gate1347(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1348(.a(s_114), .O(gate514inter3));
  inv1  gate1349(.a(s_115), .O(gate514inter4));
  nand2 gate1350(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1351(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1352(.a(G1290), .O(gate514inter7));
  inv1  gate1353(.a(G1291), .O(gate514inter8));
  nand2 gate1354(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1355(.a(s_115), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1356(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1357(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1358(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule