module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1709(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1710(.a(gate9inter0), .b(s_166), .O(gate9inter1));
  and2  gate1711(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1712(.a(s_166), .O(gate9inter3));
  inv1  gate1713(.a(s_167), .O(gate9inter4));
  nand2 gate1714(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1715(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1716(.a(G1), .O(gate9inter7));
  inv1  gate1717(.a(G2), .O(gate9inter8));
  nand2 gate1718(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1719(.a(s_167), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1720(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1721(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1722(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate911(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate912(.a(gate11inter0), .b(s_52), .O(gate11inter1));
  and2  gate913(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate914(.a(s_52), .O(gate11inter3));
  inv1  gate915(.a(s_53), .O(gate11inter4));
  nand2 gate916(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate917(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate918(.a(G5), .O(gate11inter7));
  inv1  gate919(.a(G6), .O(gate11inter8));
  nand2 gate920(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate921(.a(s_53), .b(gate11inter3), .O(gate11inter10));
  nor2  gate922(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate923(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate924(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1723(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1724(.a(gate16inter0), .b(s_168), .O(gate16inter1));
  and2  gate1725(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1726(.a(s_168), .O(gate16inter3));
  inv1  gate1727(.a(s_169), .O(gate16inter4));
  nand2 gate1728(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1729(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1730(.a(G15), .O(gate16inter7));
  inv1  gate1731(.a(G16), .O(gate16inter8));
  nand2 gate1732(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1733(.a(s_169), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1734(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1735(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1736(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1947(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1948(.a(gate18inter0), .b(s_200), .O(gate18inter1));
  and2  gate1949(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1950(.a(s_200), .O(gate18inter3));
  inv1  gate1951(.a(s_201), .O(gate18inter4));
  nand2 gate1952(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1953(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1954(.a(G19), .O(gate18inter7));
  inv1  gate1955(.a(G20), .O(gate18inter8));
  nand2 gate1956(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1957(.a(s_201), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1958(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1959(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1960(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1513(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1514(.a(gate19inter0), .b(s_138), .O(gate19inter1));
  and2  gate1515(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1516(.a(s_138), .O(gate19inter3));
  inv1  gate1517(.a(s_139), .O(gate19inter4));
  nand2 gate1518(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1519(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1520(.a(G21), .O(gate19inter7));
  inv1  gate1521(.a(G22), .O(gate19inter8));
  nand2 gate1522(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1523(.a(s_139), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1524(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1525(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1526(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate575(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate576(.a(gate23inter0), .b(s_4), .O(gate23inter1));
  and2  gate577(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate578(.a(s_4), .O(gate23inter3));
  inv1  gate579(.a(s_5), .O(gate23inter4));
  nand2 gate580(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate581(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate582(.a(G29), .O(gate23inter7));
  inv1  gate583(.a(G30), .O(gate23inter8));
  nand2 gate584(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate585(.a(s_5), .b(gate23inter3), .O(gate23inter10));
  nor2  gate586(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate587(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate588(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate547(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate548(.a(gate24inter0), .b(s_0), .O(gate24inter1));
  and2  gate549(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate550(.a(s_0), .O(gate24inter3));
  inv1  gate551(.a(s_1), .O(gate24inter4));
  nand2 gate552(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate553(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate554(.a(G31), .O(gate24inter7));
  inv1  gate555(.a(G32), .O(gate24inter8));
  nand2 gate556(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate557(.a(s_1), .b(gate24inter3), .O(gate24inter10));
  nor2  gate558(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate559(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate560(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1401(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1402(.a(gate26inter0), .b(s_122), .O(gate26inter1));
  and2  gate1403(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1404(.a(s_122), .O(gate26inter3));
  inv1  gate1405(.a(s_123), .O(gate26inter4));
  nand2 gate1406(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1407(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1408(.a(G9), .O(gate26inter7));
  inv1  gate1409(.a(G13), .O(gate26inter8));
  nand2 gate1410(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1411(.a(s_123), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1412(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1413(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1414(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1135(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1136(.a(gate30inter0), .b(s_84), .O(gate30inter1));
  and2  gate1137(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1138(.a(s_84), .O(gate30inter3));
  inv1  gate1139(.a(s_85), .O(gate30inter4));
  nand2 gate1140(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1141(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1142(.a(G11), .O(gate30inter7));
  inv1  gate1143(.a(G15), .O(gate30inter8));
  nand2 gate1144(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1145(.a(s_85), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1146(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1147(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1148(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1737(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1738(.a(gate36inter0), .b(s_170), .O(gate36inter1));
  and2  gate1739(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1740(.a(s_170), .O(gate36inter3));
  inv1  gate1741(.a(s_171), .O(gate36inter4));
  nand2 gate1742(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1743(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1744(.a(G26), .O(gate36inter7));
  inv1  gate1745(.a(G30), .O(gate36inter8));
  nand2 gate1746(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1747(.a(s_171), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1748(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1749(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1750(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate603(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate604(.a(gate37inter0), .b(s_8), .O(gate37inter1));
  and2  gate605(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate606(.a(s_8), .O(gate37inter3));
  inv1  gate607(.a(s_9), .O(gate37inter4));
  nand2 gate608(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate609(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate610(.a(G19), .O(gate37inter7));
  inv1  gate611(.a(G23), .O(gate37inter8));
  nand2 gate612(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate613(.a(s_9), .b(gate37inter3), .O(gate37inter10));
  nor2  gate614(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate615(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate616(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1807(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1808(.a(gate38inter0), .b(s_180), .O(gate38inter1));
  and2  gate1809(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1810(.a(s_180), .O(gate38inter3));
  inv1  gate1811(.a(s_181), .O(gate38inter4));
  nand2 gate1812(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1813(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1814(.a(G27), .O(gate38inter7));
  inv1  gate1815(.a(G31), .O(gate38inter8));
  nand2 gate1816(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1817(.a(s_181), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1818(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1819(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1820(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1163(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1164(.a(gate40inter0), .b(s_88), .O(gate40inter1));
  and2  gate1165(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1166(.a(s_88), .O(gate40inter3));
  inv1  gate1167(.a(s_89), .O(gate40inter4));
  nand2 gate1168(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1169(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1170(.a(G28), .O(gate40inter7));
  inv1  gate1171(.a(G32), .O(gate40inter8));
  nand2 gate1172(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1173(.a(s_89), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1174(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1175(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1176(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1415(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1416(.a(gate49inter0), .b(s_124), .O(gate49inter1));
  and2  gate1417(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1418(.a(s_124), .O(gate49inter3));
  inv1  gate1419(.a(s_125), .O(gate49inter4));
  nand2 gate1420(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1421(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1422(.a(G9), .O(gate49inter7));
  inv1  gate1423(.a(G278), .O(gate49inter8));
  nand2 gate1424(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1425(.a(s_125), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1426(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1427(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1428(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1275(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1276(.a(gate50inter0), .b(s_104), .O(gate50inter1));
  and2  gate1277(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1278(.a(s_104), .O(gate50inter3));
  inv1  gate1279(.a(s_105), .O(gate50inter4));
  nand2 gate1280(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1281(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1282(.a(G10), .O(gate50inter7));
  inv1  gate1283(.a(G278), .O(gate50inter8));
  nand2 gate1284(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1285(.a(s_105), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1286(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1287(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1288(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate841(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate842(.a(gate57inter0), .b(s_42), .O(gate57inter1));
  and2  gate843(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate844(.a(s_42), .O(gate57inter3));
  inv1  gate845(.a(s_43), .O(gate57inter4));
  nand2 gate846(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate847(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate848(.a(G17), .O(gate57inter7));
  inv1  gate849(.a(G290), .O(gate57inter8));
  nand2 gate850(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate851(.a(s_43), .b(gate57inter3), .O(gate57inter10));
  nor2  gate852(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate853(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate854(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1219(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1220(.a(gate60inter0), .b(s_96), .O(gate60inter1));
  and2  gate1221(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1222(.a(s_96), .O(gate60inter3));
  inv1  gate1223(.a(s_97), .O(gate60inter4));
  nand2 gate1224(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1225(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1226(.a(G20), .O(gate60inter7));
  inv1  gate1227(.a(G293), .O(gate60inter8));
  nand2 gate1228(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1229(.a(s_97), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1230(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1231(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1232(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1835(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1836(.a(gate62inter0), .b(s_184), .O(gate62inter1));
  and2  gate1837(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1838(.a(s_184), .O(gate62inter3));
  inv1  gate1839(.a(s_185), .O(gate62inter4));
  nand2 gate1840(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1841(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1842(.a(G22), .O(gate62inter7));
  inv1  gate1843(.a(G296), .O(gate62inter8));
  nand2 gate1844(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1845(.a(s_185), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1846(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1847(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1848(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2073(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2074(.a(gate74inter0), .b(s_218), .O(gate74inter1));
  and2  gate2075(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2076(.a(s_218), .O(gate74inter3));
  inv1  gate2077(.a(s_219), .O(gate74inter4));
  nand2 gate2078(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2079(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2080(.a(G5), .O(gate74inter7));
  inv1  gate2081(.a(G314), .O(gate74inter8));
  nand2 gate2082(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2083(.a(s_219), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2084(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2085(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2086(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1303(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1304(.a(gate81inter0), .b(s_108), .O(gate81inter1));
  and2  gate1305(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1306(.a(s_108), .O(gate81inter3));
  inv1  gate1307(.a(s_109), .O(gate81inter4));
  nand2 gate1308(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1309(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1310(.a(G3), .O(gate81inter7));
  inv1  gate1311(.a(G326), .O(gate81inter8));
  nand2 gate1312(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1313(.a(s_109), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1314(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1315(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1316(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1597(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1598(.a(gate82inter0), .b(s_150), .O(gate82inter1));
  and2  gate1599(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1600(.a(s_150), .O(gate82inter3));
  inv1  gate1601(.a(s_151), .O(gate82inter4));
  nand2 gate1602(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1603(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1604(.a(G7), .O(gate82inter7));
  inv1  gate1605(.a(G326), .O(gate82inter8));
  nand2 gate1606(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1607(.a(s_151), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1608(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1609(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1610(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate743(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate744(.a(gate86inter0), .b(s_28), .O(gate86inter1));
  and2  gate745(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate746(.a(s_28), .O(gate86inter3));
  inv1  gate747(.a(s_29), .O(gate86inter4));
  nand2 gate748(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate749(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate750(.a(G8), .O(gate86inter7));
  inv1  gate751(.a(G332), .O(gate86inter8));
  nand2 gate752(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate753(.a(s_29), .b(gate86inter3), .O(gate86inter10));
  nor2  gate754(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate755(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate756(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate659(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate660(.a(gate87inter0), .b(s_16), .O(gate87inter1));
  and2  gate661(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate662(.a(s_16), .O(gate87inter3));
  inv1  gate663(.a(s_17), .O(gate87inter4));
  nand2 gate664(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate665(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate666(.a(G12), .O(gate87inter7));
  inv1  gate667(.a(G335), .O(gate87inter8));
  nand2 gate668(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate669(.a(s_17), .b(gate87inter3), .O(gate87inter10));
  nor2  gate670(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate671(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate672(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1541(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1542(.a(gate90inter0), .b(s_142), .O(gate90inter1));
  and2  gate1543(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1544(.a(s_142), .O(gate90inter3));
  inv1  gate1545(.a(s_143), .O(gate90inter4));
  nand2 gate1546(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1547(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1548(.a(G21), .O(gate90inter7));
  inv1  gate1549(.a(G338), .O(gate90inter8));
  nand2 gate1550(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1551(.a(s_143), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1552(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1553(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1554(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1443(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1444(.a(gate91inter0), .b(s_128), .O(gate91inter1));
  and2  gate1445(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1446(.a(s_128), .O(gate91inter3));
  inv1  gate1447(.a(s_129), .O(gate91inter4));
  nand2 gate1448(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1449(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1450(.a(G25), .O(gate91inter7));
  inv1  gate1451(.a(G341), .O(gate91inter8));
  nand2 gate1452(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1453(.a(s_129), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1454(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1455(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1456(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate771(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate772(.a(gate96inter0), .b(s_32), .O(gate96inter1));
  and2  gate773(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate774(.a(s_32), .O(gate96inter3));
  inv1  gate775(.a(s_33), .O(gate96inter4));
  nand2 gate776(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate777(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate778(.a(G30), .O(gate96inter7));
  inv1  gate779(.a(G347), .O(gate96inter8));
  nand2 gate780(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate781(.a(s_33), .b(gate96inter3), .O(gate96inter10));
  nor2  gate782(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate783(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate784(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate883(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate884(.a(gate101inter0), .b(s_48), .O(gate101inter1));
  and2  gate885(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate886(.a(s_48), .O(gate101inter3));
  inv1  gate887(.a(s_49), .O(gate101inter4));
  nand2 gate888(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate889(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate890(.a(G20), .O(gate101inter7));
  inv1  gate891(.a(G356), .O(gate101inter8));
  nand2 gate892(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate893(.a(s_49), .b(gate101inter3), .O(gate101inter10));
  nor2  gate894(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate895(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate896(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate981(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate982(.a(gate108inter0), .b(s_62), .O(gate108inter1));
  and2  gate983(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate984(.a(s_62), .O(gate108inter3));
  inv1  gate985(.a(s_63), .O(gate108inter4));
  nand2 gate986(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate987(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate988(.a(G368), .O(gate108inter7));
  inv1  gate989(.a(G369), .O(gate108inter8));
  nand2 gate990(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate991(.a(s_63), .b(gate108inter3), .O(gate108inter10));
  nor2  gate992(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate993(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate994(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1611(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1612(.a(gate111inter0), .b(s_152), .O(gate111inter1));
  and2  gate1613(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1614(.a(s_152), .O(gate111inter3));
  inv1  gate1615(.a(s_153), .O(gate111inter4));
  nand2 gate1616(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1617(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1618(.a(G374), .O(gate111inter7));
  inv1  gate1619(.a(G375), .O(gate111inter8));
  nand2 gate1620(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1621(.a(s_153), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1622(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1623(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1624(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1569(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1570(.a(gate112inter0), .b(s_146), .O(gate112inter1));
  and2  gate1571(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1572(.a(s_146), .O(gate112inter3));
  inv1  gate1573(.a(s_147), .O(gate112inter4));
  nand2 gate1574(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1575(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1576(.a(G376), .O(gate112inter7));
  inv1  gate1577(.a(G377), .O(gate112inter8));
  nand2 gate1578(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1579(.a(s_147), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1580(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1581(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1582(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1289(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1290(.a(gate113inter0), .b(s_106), .O(gate113inter1));
  and2  gate1291(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1292(.a(s_106), .O(gate113inter3));
  inv1  gate1293(.a(s_107), .O(gate113inter4));
  nand2 gate1294(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1295(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1296(.a(G378), .O(gate113inter7));
  inv1  gate1297(.a(G379), .O(gate113inter8));
  nand2 gate1298(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1299(.a(s_107), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1300(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1301(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1302(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate561(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate562(.a(gate119inter0), .b(s_2), .O(gate119inter1));
  and2  gate563(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate564(.a(s_2), .O(gate119inter3));
  inv1  gate565(.a(s_3), .O(gate119inter4));
  nand2 gate566(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate567(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate568(.a(G390), .O(gate119inter7));
  inv1  gate569(.a(G391), .O(gate119inter8));
  nand2 gate570(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate571(.a(s_3), .b(gate119inter3), .O(gate119inter10));
  nor2  gate572(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate573(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate574(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2157(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2158(.a(gate122inter0), .b(s_230), .O(gate122inter1));
  and2  gate2159(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2160(.a(s_230), .O(gate122inter3));
  inv1  gate2161(.a(s_231), .O(gate122inter4));
  nand2 gate2162(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2163(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2164(.a(G396), .O(gate122inter7));
  inv1  gate2165(.a(G397), .O(gate122inter8));
  nand2 gate2166(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2167(.a(s_231), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2168(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2169(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2170(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1527(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1528(.a(gate123inter0), .b(s_140), .O(gate123inter1));
  and2  gate1529(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1530(.a(s_140), .O(gate123inter3));
  inv1  gate1531(.a(s_141), .O(gate123inter4));
  nand2 gate1532(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1533(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1534(.a(G398), .O(gate123inter7));
  inv1  gate1535(.a(G399), .O(gate123inter8));
  nand2 gate1536(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1537(.a(s_141), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1538(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1539(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1540(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate967(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate968(.a(gate125inter0), .b(s_60), .O(gate125inter1));
  and2  gate969(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate970(.a(s_60), .O(gate125inter3));
  inv1  gate971(.a(s_61), .O(gate125inter4));
  nand2 gate972(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate973(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate974(.a(G402), .O(gate125inter7));
  inv1  gate975(.a(G403), .O(gate125inter8));
  nand2 gate976(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate977(.a(s_61), .b(gate125inter3), .O(gate125inter10));
  nor2  gate978(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate979(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate980(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1065(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1066(.a(gate126inter0), .b(s_74), .O(gate126inter1));
  and2  gate1067(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1068(.a(s_74), .O(gate126inter3));
  inv1  gate1069(.a(s_75), .O(gate126inter4));
  nand2 gate1070(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1071(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1072(.a(G404), .O(gate126inter7));
  inv1  gate1073(.a(G405), .O(gate126inter8));
  nand2 gate1074(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1075(.a(s_75), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1076(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1077(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1078(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1247(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1248(.a(gate128inter0), .b(s_100), .O(gate128inter1));
  and2  gate1249(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1250(.a(s_100), .O(gate128inter3));
  inv1  gate1251(.a(s_101), .O(gate128inter4));
  nand2 gate1252(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1253(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1254(.a(G408), .O(gate128inter7));
  inv1  gate1255(.a(G409), .O(gate128inter8));
  nand2 gate1256(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1257(.a(s_101), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1258(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1259(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1260(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1905(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1906(.a(gate129inter0), .b(s_194), .O(gate129inter1));
  and2  gate1907(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1908(.a(s_194), .O(gate129inter3));
  inv1  gate1909(.a(s_195), .O(gate129inter4));
  nand2 gate1910(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1911(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1912(.a(G410), .O(gate129inter7));
  inv1  gate1913(.a(G411), .O(gate129inter8));
  nand2 gate1914(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1915(.a(s_195), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1916(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1917(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1918(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate757(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate758(.a(gate135inter0), .b(s_30), .O(gate135inter1));
  and2  gate759(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate760(.a(s_30), .O(gate135inter3));
  inv1  gate761(.a(s_31), .O(gate135inter4));
  nand2 gate762(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate763(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate764(.a(G422), .O(gate135inter7));
  inv1  gate765(.a(G423), .O(gate135inter8));
  nand2 gate766(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate767(.a(s_31), .b(gate135inter3), .O(gate135inter10));
  nor2  gate768(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate769(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate770(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1331(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1332(.a(gate136inter0), .b(s_112), .O(gate136inter1));
  and2  gate1333(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1334(.a(s_112), .O(gate136inter3));
  inv1  gate1335(.a(s_113), .O(gate136inter4));
  nand2 gate1336(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1337(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1338(.a(G424), .O(gate136inter7));
  inv1  gate1339(.a(G425), .O(gate136inter8));
  nand2 gate1340(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1341(.a(s_113), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1342(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1343(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1344(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1681(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1682(.a(gate138inter0), .b(s_162), .O(gate138inter1));
  and2  gate1683(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1684(.a(s_162), .O(gate138inter3));
  inv1  gate1685(.a(s_163), .O(gate138inter4));
  nand2 gate1686(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1687(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1688(.a(G432), .O(gate138inter7));
  inv1  gate1689(.a(G435), .O(gate138inter8));
  nand2 gate1690(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1691(.a(s_163), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1692(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1693(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1694(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1009(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1010(.a(gate146inter0), .b(s_66), .O(gate146inter1));
  and2  gate1011(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1012(.a(s_66), .O(gate146inter3));
  inv1  gate1013(.a(s_67), .O(gate146inter4));
  nand2 gate1014(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1015(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1016(.a(G480), .O(gate146inter7));
  inv1  gate1017(.a(G483), .O(gate146inter8));
  nand2 gate1018(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1019(.a(s_67), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1020(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1021(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1022(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1583(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1584(.a(gate149inter0), .b(s_148), .O(gate149inter1));
  and2  gate1585(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1586(.a(s_148), .O(gate149inter3));
  inv1  gate1587(.a(s_149), .O(gate149inter4));
  nand2 gate1588(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1589(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1590(.a(G498), .O(gate149inter7));
  inv1  gate1591(.a(G501), .O(gate149inter8));
  nand2 gate1592(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1593(.a(s_149), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1594(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1595(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1596(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate799(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate800(.a(gate156inter0), .b(s_36), .O(gate156inter1));
  and2  gate801(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate802(.a(s_36), .O(gate156inter3));
  inv1  gate803(.a(s_37), .O(gate156inter4));
  nand2 gate804(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate805(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate806(.a(G435), .O(gate156inter7));
  inv1  gate807(.a(G525), .O(gate156inter8));
  nand2 gate808(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate809(.a(s_37), .b(gate156inter3), .O(gate156inter10));
  nor2  gate810(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate811(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate812(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1261(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1262(.a(gate157inter0), .b(s_102), .O(gate157inter1));
  and2  gate1263(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1264(.a(s_102), .O(gate157inter3));
  inv1  gate1265(.a(s_103), .O(gate157inter4));
  nand2 gate1266(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1267(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1268(.a(G438), .O(gate157inter7));
  inv1  gate1269(.a(G528), .O(gate157inter8));
  nand2 gate1270(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1271(.a(s_103), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1272(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1273(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1274(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1695(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1696(.a(gate159inter0), .b(s_164), .O(gate159inter1));
  and2  gate1697(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1698(.a(s_164), .O(gate159inter3));
  inv1  gate1699(.a(s_165), .O(gate159inter4));
  nand2 gate1700(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1701(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1702(.a(G444), .O(gate159inter7));
  inv1  gate1703(.a(G531), .O(gate159inter8));
  nand2 gate1704(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1705(.a(s_165), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1706(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1707(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1708(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1387(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1388(.a(gate160inter0), .b(s_120), .O(gate160inter1));
  and2  gate1389(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1390(.a(s_120), .O(gate160inter3));
  inv1  gate1391(.a(s_121), .O(gate160inter4));
  nand2 gate1392(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1393(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1394(.a(G447), .O(gate160inter7));
  inv1  gate1395(.a(G531), .O(gate160inter8));
  nand2 gate1396(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1397(.a(s_121), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1398(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1399(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1400(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1359(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1360(.a(gate168inter0), .b(s_116), .O(gate168inter1));
  and2  gate1361(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1362(.a(s_116), .O(gate168inter3));
  inv1  gate1363(.a(s_117), .O(gate168inter4));
  nand2 gate1364(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1365(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1366(.a(G471), .O(gate168inter7));
  inv1  gate1367(.a(G543), .O(gate168inter8));
  nand2 gate1368(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1369(.a(s_117), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1370(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1371(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1372(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1457(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1458(.a(gate169inter0), .b(s_130), .O(gate169inter1));
  and2  gate1459(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1460(.a(s_130), .O(gate169inter3));
  inv1  gate1461(.a(s_131), .O(gate169inter4));
  nand2 gate1462(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1463(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1464(.a(G474), .O(gate169inter7));
  inv1  gate1465(.a(G546), .O(gate169inter8));
  nand2 gate1466(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1467(.a(s_131), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1468(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1469(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1470(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate715(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate716(.a(gate172inter0), .b(s_24), .O(gate172inter1));
  and2  gate717(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate718(.a(s_24), .O(gate172inter3));
  inv1  gate719(.a(s_25), .O(gate172inter4));
  nand2 gate720(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate721(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate722(.a(G483), .O(gate172inter7));
  inv1  gate723(.a(G549), .O(gate172inter8));
  nand2 gate724(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate725(.a(s_25), .b(gate172inter3), .O(gate172inter10));
  nor2  gate726(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate727(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate728(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1205(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1206(.a(gate175inter0), .b(s_94), .O(gate175inter1));
  and2  gate1207(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1208(.a(s_94), .O(gate175inter3));
  inv1  gate1209(.a(s_95), .O(gate175inter4));
  nand2 gate1210(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1211(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1212(.a(G492), .O(gate175inter7));
  inv1  gate1213(.a(G555), .O(gate175inter8));
  nand2 gate1214(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1215(.a(s_95), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1216(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1217(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1218(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2045(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2046(.a(gate180inter0), .b(s_214), .O(gate180inter1));
  and2  gate2047(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2048(.a(s_214), .O(gate180inter3));
  inv1  gate2049(.a(s_215), .O(gate180inter4));
  nand2 gate2050(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2051(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2052(.a(G507), .O(gate180inter7));
  inv1  gate2053(.a(G561), .O(gate180inter8));
  nand2 gate2054(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2055(.a(s_215), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2056(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2057(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2058(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1051(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1052(.a(gate181inter0), .b(s_72), .O(gate181inter1));
  and2  gate1053(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1054(.a(s_72), .O(gate181inter3));
  inv1  gate1055(.a(s_73), .O(gate181inter4));
  nand2 gate1056(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1057(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1058(.a(G510), .O(gate181inter7));
  inv1  gate1059(.a(G564), .O(gate181inter8));
  nand2 gate1060(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1061(.a(s_73), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1062(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1063(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1064(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1485(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1486(.a(gate186inter0), .b(s_134), .O(gate186inter1));
  and2  gate1487(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1488(.a(s_134), .O(gate186inter3));
  inv1  gate1489(.a(s_135), .O(gate186inter4));
  nand2 gate1490(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1491(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1492(.a(G572), .O(gate186inter7));
  inv1  gate1493(.a(G573), .O(gate186inter8));
  nand2 gate1494(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1495(.a(s_135), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1496(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1497(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1498(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1317(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1318(.a(gate187inter0), .b(s_110), .O(gate187inter1));
  and2  gate1319(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1320(.a(s_110), .O(gate187inter3));
  inv1  gate1321(.a(s_111), .O(gate187inter4));
  nand2 gate1322(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1323(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1324(.a(G574), .O(gate187inter7));
  inv1  gate1325(.a(G575), .O(gate187inter8));
  nand2 gate1326(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1327(.a(s_111), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1328(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1329(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1330(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate2129(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2130(.a(gate199inter0), .b(s_226), .O(gate199inter1));
  and2  gate2131(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2132(.a(s_226), .O(gate199inter3));
  inv1  gate2133(.a(s_227), .O(gate199inter4));
  nand2 gate2134(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2135(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2136(.a(G598), .O(gate199inter7));
  inv1  gate2137(.a(G599), .O(gate199inter8));
  nand2 gate2138(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2139(.a(s_227), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2140(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2141(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2142(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1765(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1766(.a(gate203inter0), .b(s_174), .O(gate203inter1));
  and2  gate1767(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1768(.a(s_174), .O(gate203inter3));
  inv1  gate1769(.a(s_175), .O(gate203inter4));
  nand2 gate1770(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1771(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1772(.a(G602), .O(gate203inter7));
  inv1  gate1773(.a(G612), .O(gate203inter8));
  nand2 gate1774(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1775(.a(s_175), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1776(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1777(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1778(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate827(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate828(.a(gate205inter0), .b(s_40), .O(gate205inter1));
  and2  gate829(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate830(.a(s_40), .O(gate205inter3));
  inv1  gate831(.a(s_41), .O(gate205inter4));
  nand2 gate832(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate833(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate834(.a(G622), .O(gate205inter7));
  inv1  gate835(.a(G627), .O(gate205inter8));
  nand2 gate836(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate837(.a(s_41), .b(gate205inter3), .O(gate205inter10));
  nor2  gate838(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate839(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate840(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2101(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2102(.a(gate217inter0), .b(s_222), .O(gate217inter1));
  and2  gate2103(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2104(.a(s_222), .O(gate217inter3));
  inv1  gate2105(.a(s_223), .O(gate217inter4));
  nand2 gate2106(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2107(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2108(.a(G622), .O(gate217inter7));
  inv1  gate2109(.a(G678), .O(gate217inter8));
  nand2 gate2110(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2111(.a(s_223), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2112(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2113(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2114(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate589(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate590(.a(gate218inter0), .b(s_6), .O(gate218inter1));
  and2  gate591(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate592(.a(s_6), .O(gate218inter3));
  inv1  gate593(.a(s_7), .O(gate218inter4));
  nand2 gate594(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate595(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate596(.a(G627), .O(gate218inter7));
  inv1  gate597(.a(G678), .O(gate218inter8));
  nand2 gate598(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate599(.a(s_7), .b(gate218inter3), .O(gate218inter10));
  nor2  gate600(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate601(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate602(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate813(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate814(.a(gate230inter0), .b(s_38), .O(gate230inter1));
  and2  gate815(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate816(.a(s_38), .O(gate230inter3));
  inv1  gate817(.a(s_39), .O(gate230inter4));
  nand2 gate818(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate819(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate820(.a(G700), .O(gate230inter7));
  inv1  gate821(.a(G701), .O(gate230inter8));
  nand2 gate822(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate823(.a(s_39), .b(gate230inter3), .O(gate230inter10));
  nor2  gate824(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate825(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate826(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1653(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1654(.a(gate231inter0), .b(s_158), .O(gate231inter1));
  and2  gate1655(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1656(.a(s_158), .O(gate231inter3));
  inv1  gate1657(.a(s_159), .O(gate231inter4));
  nand2 gate1658(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1659(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1660(.a(G702), .O(gate231inter7));
  inv1  gate1661(.a(G703), .O(gate231inter8));
  nand2 gate1662(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1663(.a(s_159), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1664(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1665(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1666(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate939(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate940(.a(gate236inter0), .b(s_56), .O(gate236inter1));
  and2  gate941(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate942(.a(s_56), .O(gate236inter3));
  inv1  gate943(.a(s_57), .O(gate236inter4));
  nand2 gate944(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate945(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate946(.a(G251), .O(gate236inter7));
  inv1  gate947(.a(G727), .O(gate236inter8));
  nand2 gate948(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate949(.a(s_57), .b(gate236inter3), .O(gate236inter10));
  nor2  gate950(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate951(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate952(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2087(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2088(.a(gate238inter0), .b(s_220), .O(gate238inter1));
  and2  gate2089(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2090(.a(s_220), .O(gate238inter3));
  inv1  gate2091(.a(s_221), .O(gate238inter4));
  nand2 gate2092(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2093(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2094(.a(G257), .O(gate238inter7));
  inv1  gate2095(.a(G709), .O(gate238inter8));
  nand2 gate2096(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2097(.a(s_221), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2098(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2099(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2100(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1975(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1976(.a(gate240inter0), .b(s_204), .O(gate240inter1));
  and2  gate1977(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1978(.a(s_204), .O(gate240inter3));
  inv1  gate1979(.a(s_205), .O(gate240inter4));
  nand2 gate1980(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1981(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1982(.a(G263), .O(gate240inter7));
  inv1  gate1983(.a(G715), .O(gate240inter8));
  nand2 gate1984(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1985(.a(s_205), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1986(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1987(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1988(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate729(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate730(.a(gate242inter0), .b(s_26), .O(gate242inter1));
  and2  gate731(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate732(.a(s_26), .O(gate242inter3));
  inv1  gate733(.a(s_27), .O(gate242inter4));
  nand2 gate734(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate735(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate736(.a(G718), .O(gate242inter7));
  inv1  gate737(.a(G730), .O(gate242inter8));
  nand2 gate738(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate739(.a(s_27), .b(gate242inter3), .O(gate242inter10));
  nor2  gate740(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate741(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate742(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1429(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1430(.a(gate243inter0), .b(s_126), .O(gate243inter1));
  and2  gate1431(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1432(.a(s_126), .O(gate243inter3));
  inv1  gate1433(.a(s_127), .O(gate243inter4));
  nand2 gate1434(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1435(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1436(.a(G245), .O(gate243inter7));
  inv1  gate1437(.a(G733), .O(gate243inter8));
  nand2 gate1438(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1439(.a(s_127), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1440(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1441(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1442(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2143(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2144(.a(gate251inter0), .b(s_228), .O(gate251inter1));
  and2  gate2145(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2146(.a(s_228), .O(gate251inter3));
  inv1  gate2147(.a(s_229), .O(gate251inter4));
  nand2 gate2148(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2149(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2150(.a(G257), .O(gate251inter7));
  inv1  gate2151(.a(G745), .O(gate251inter8));
  nand2 gate2152(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2153(.a(s_229), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2154(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2155(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2156(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate631(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate632(.a(gate257inter0), .b(s_12), .O(gate257inter1));
  and2  gate633(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate634(.a(s_12), .O(gate257inter3));
  inv1  gate635(.a(s_13), .O(gate257inter4));
  nand2 gate636(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate637(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate638(.a(G754), .O(gate257inter7));
  inv1  gate639(.a(G755), .O(gate257inter8));
  nand2 gate640(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate641(.a(s_13), .b(gate257inter3), .O(gate257inter10));
  nor2  gate642(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate643(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate644(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate925(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate926(.a(gate259inter0), .b(s_54), .O(gate259inter1));
  and2  gate927(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate928(.a(s_54), .O(gate259inter3));
  inv1  gate929(.a(s_55), .O(gate259inter4));
  nand2 gate930(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate931(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate932(.a(G758), .O(gate259inter7));
  inv1  gate933(.a(G759), .O(gate259inter8));
  nand2 gate934(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate935(.a(s_55), .b(gate259inter3), .O(gate259inter10));
  nor2  gate936(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate937(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate938(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate673(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate674(.a(gate262inter0), .b(s_18), .O(gate262inter1));
  and2  gate675(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate676(.a(s_18), .O(gate262inter3));
  inv1  gate677(.a(s_19), .O(gate262inter4));
  nand2 gate678(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate679(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate680(.a(G764), .O(gate262inter7));
  inv1  gate681(.a(G765), .O(gate262inter8));
  nand2 gate682(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate683(.a(s_19), .b(gate262inter3), .O(gate262inter10));
  nor2  gate684(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate685(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate686(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1639(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1640(.a(gate268inter0), .b(s_156), .O(gate268inter1));
  and2  gate1641(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1642(.a(s_156), .O(gate268inter3));
  inv1  gate1643(.a(s_157), .O(gate268inter4));
  nand2 gate1644(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1645(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1646(.a(G651), .O(gate268inter7));
  inv1  gate1647(.a(G779), .O(gate268inter8));
  nand2 gate1648(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1649(.a(s_157), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1650(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1651(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1652(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1037(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1038(.a(gate270inter0), .b(s_70), .O(gate270inter1));
  and2  gate1039(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1040(.a(s_70), .O(gate270inter3));
  inv1  gate1041(.a(s_71), .O(gate270inter4));
  nand2 gate1042(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1043(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1044(.a(G657), .O(gate270inter7));
  inv1  gate1045(.a(G785), .O(gate270inter8));
  nand2 gate1046(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1047(.a(s_71), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1048(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1049(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1050(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1373(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1374(.a(gate271inter0), .b(s_118), .O(gate271inter1));
  and2  gate1375(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1376(.a(s_118), .O(gate271inter3));
  inv1  gate1377(.a(s_119), .O(gate271inter4));
  nand2 gate1378(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1379(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1380(.a(G660), .O(gate271inter7));
  inv1  gate1381(.a(G788), .O(gate271inter8));
  nand2 gate1382(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1383(.a(s_119), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1384(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1385(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1386(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate645(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate646(.a(gate278inter0), .b(s_14), .O(gate278inter1));
  and2  gate647(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate648(.a(s_14), .O(gate278inter3));
  inv1  gate649(.a(s_15), .O(gate278inter4));
  nand2 gate650(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate651(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate652(.a(G776), .O(gate278inter7));
  inv1  gate653(.a(G800), .O(gate278inter8));
  nand2 gate654(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate655(.a(s_15), .b(gate278inter3), .O(gate278inter10));
  nor2  gate656(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate657(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate658(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1779(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1780(.a(gate279inter0), .b(s_176), .O(gate279inter1));
  and2  gate1781(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1782(.a(s_176), .O(gate279inter3));
  inv1  gate1783(.a(s_177), .O(gate279inter4));
  nand2 gate1784(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1785(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1786(.a(G651), .O(gate279inter7));
  inv1  gate1787(.a(G803), .O(gate279inter8));
  nand2 gate1788(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1789(.a(s_177), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1790(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1791(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1792(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1919(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1920(.a(gate283inter0), .b(s_196), .O(gate283inter1));
  and2  gate1921(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1922(.a(s_196), .O(gate283inter3));
  inv1  gate1923(.a(s_197), .O(gate283inter4));
  nand2 gate1924(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1925(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1926(.a(G657), .O(gate283inter7));
  inv1  gate1927(.a(G809), .O(gate283inter8));
  nand2 gate1928(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1929(.a(s_197), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1930(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1931(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1932(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1023(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1024(.a(gate288inter0), .b(s_68), .O(gate288inter1));
  and2  gate1025(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1026(.a(s_68), .O(gate288inter3));
  inv1  gate1027(.a(s_69), .O(gate288inter4));
  nand2 gate1028(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1029(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1030(.a(G791), .O(gate288inter7));
  inv1  gate1031(.a(G815), .O(gate288inter8));
  nand2 gate1032(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1033(.a(s_69), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1034(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1035(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1036(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1191(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1192(.a(gate290inter0), .b(s_92), .O(gate290inter1));
  and2  gate1193(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1194(.a(s_92), .O(gate290inter3));
  inv1  gate1195(.a(s_93), .O(gate290inter4));
  nand2 gate1196(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1197(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1198(.a(G820), .O(gate290inter7));
  inv1  gate1199(.a(G821), .O(gate290inter8));
  nand2 gate1200(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1201(.a(s_93), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1202(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1203(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1204(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1345(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1346(.a(gate292inter0), .b(s_114), .O(gate292inter1));
  and2  gate1347(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1348(.a(s_114), .O(gate292inter3));
  inv1  gate1349(.a(s_115), .O(gate292inter4));
  nand2 gate1350(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1351(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1352(.a(G824), .O(gate292inter7));
  inv1  gate1353(.a(G825), .O(gate292inter8));
  nand2 gate1354(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1355(.a(s_115), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1356(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1357(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1358(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1849(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1850(.a(gate387inter0), .b(s_186), .O(gate387inter1));
  and2  gate1851(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1852(.a(s_186), .O(gate387inter3));
  inv1  gate1853(.a(s_187), .O(gate387inter4));
  nand2 gate1854(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1855(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1856(.a(G1), .O(gate387inter7));
  inv1  gate1857(.a(G1036), .O(gate387inter8));
  nand2 gate1858(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1859(.a(s_187), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1860(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1861(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1862(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate953(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate954(.a(gate389inter0), .b(s_58), .O(gate389inter1));
  and2  gate955(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate956(.a(s_58), .O(gate389inter3));
  inv1  gate957(.a(s_59), .O(gate389inter4));
  nand2 gate958(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate959(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate960(.a(G3), .O(gate389inter7));
  inv1  gate961(.a(G1042), .O(gate389inter8));
  nand2 gate962(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate963(.a(s_59), .b(gate389inter3), .O(gate389inter10));
  nor2  gate964(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate965(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate966(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1989(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1990(.a(gate390inter0), .b(s_206), .O(gate390inter1));
  and2  gate1991(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1992(.a(s_206), .O(gate390inter3));
  inv1  gate1993(.a(s_207), .O(gate390inter4));
  nand2 gate1994(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1995(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1996(.a(G4), .O(gate390inter7));
  inv1  gate1997(.a(G1045), .O(gate390inter8));
  nand2 gate1998(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1999(.a(s_207), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2000(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2001(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2002(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate855(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate856(.a(gate391inter0), .b(s_44), .O(gate391inter1));
  and2  gate857(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate858(.a(s_44), .O(gate391inter3));
  inv1  gate859(.a(s_45), .O(gate391inter4));
  nand2 gate860(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate861(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate862(.a(G5), .O(gate391inter7));
  inv1  gate863(.a(G1048), .O(gate391inter8));
  nand2 gate864(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate865(.a(s_45), .b(gate391inter3), .O(gate391inter10));
  nor2  gate866(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate867(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate868(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2003(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2004(.a(gate409inter0), .b(s_208), .O(gate409inter1));
  and2  gate2005(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2006(.a(s_208), .O(gate409inter3));
  inv1  gate2007(.a(s_209), .O(gate409inter4));
  nand2 gate2008(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2009(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2010(.a(G23), .O(gate409inter7));
  inv1  gate2011(.a(G1102), .O(gate409inter8));
  nand2 gate2012(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2013(.a(s_209), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2014(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2015(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2016(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1751(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1752(.a(gate412inter0), .b(s_172), .O(gate412inter1));
  and2  gate1753(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1754(.a(s_172), .O(gate412inter3));
  inv1  gate1755(.a(s_173), .O(gate412inter4));
  nand2 gate1756(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1757(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1758(.a(G26), .O(gate412inter7));
  inv1  gate1759(.a(G1111), .O(gate412inter8));
  nand2 gate1760(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1761(.a(s_173), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1762(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1763(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1764(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate995(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate996(.a(gate419inter0), .b(s_64), .O(gate419inter1));
  and2  gate997(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate998(.a(s_64), .O(gate419inter3));
  inv1  gate999(.a(s_65), .O(gate419inter4));
  nand2 gate1000(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1001(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1002(.a(G1), .O(gate419inter7));
  inv1  gate1003(.a(G1132), .O(gate419inter8));
  nand2 gate1004(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1005(.a(s_65), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1006(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1007(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1008(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate687(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate688(.a(gate420inter0), .b(s_20), .O(gate420inter1));
  and2  gate689(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate690(.a(s_20), .O(gate420inter3));
  inv1  gate691(.a(s_21), .O(gate420inter4));
  nand2 gate692(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate693(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate694(.a(G1036), .O(gate420inter7));
  inv1  gate695(.a(G1132), .O(gate420inter8));
  nand2 gate696(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate697(.a(s_21), .b(gate420inter3), .O(gate420inter10));
  nor2  gate698(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate699(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate700(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1093(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1094(.a(gate422inter0), .b(s_78), .O(gate422inter1));
  and2  gate1095(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1096(.a(s_78), .O(gate422inter3));
  inv1  gate1097(.a(s_79), .O(gate422inter4));
  nand2 gate1098(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1099(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1100(.a(G1039), .O(gate422inter7));
  inv1  gate1101(.a(G1135), .O(gate422inter8));
  nand2 gate1102(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1103(.a(s_79), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1104(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1105(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1106(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate869(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate870(.a(gate423inter0), .b(s_46), .O(gate423inter1));
  and2  gate871(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate872(.a(s_46), .O(gate423inter3));
  inv1  gate873(.a(s_47), .O(gate423inter4));
  nand2 gate874(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate875(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate876(.a(G3), .O(gate423inter7));
  inv1  gate877(.a(G1138), .O(gate423inter8));
  nand2 gate878(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate879(.a(s_47), .b(gate423inter3), .O(gate423inter10));
  nor2  gate880(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate881(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate882(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate617(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate618(.a(gate428inter0), .b(s_10), .O(gate428inter1));
  and2  gate619(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate620(.a(s_10), .O(gate428inter3));
  inv1  gate621(.a(s_11), .O(gate428inter4));
  nand2 gate622(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate623(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate624(.a(G1048), .O(gate428inter7));
  inv1  gate625(.a(G1144), .O(gate428inter8));
  nand2 gate626(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate627(.a(s_11), .b(gate428inter3), .O(gate428inter10));
  nor2  gate628(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate629(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate630(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1233(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1234(.a(gate429inter0), .b(s_98), .O(gate429inter1));
  and2  gate1235(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1236(.a(s_98), .O(gate429inter3));
  inv1  gate1237(.a(s_99), .O(gate429inter4));
  nand2 gate1238(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1239(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1240(.a(G6), .O(gate429inter7));
  inv1  gate1241(.a(G1147), .O(gate429inter8));
  nand2 gate1242(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1243(.a(s_99), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1244(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1245(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1246(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1149(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1150(.a(gate430inter0), .b(s_86), .O(gate430inter1));
  and2  gate1151(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1152(.a(s_86), .O(gate430inter3));
  inv1  gate1153(.a(s_87), .O(gate430inter4));
  nand2 gate1154(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1155(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1156(.a(G1051), .O(gate430inter7));
  inv1  gate1157(.a(G1147), .O(gate430inter8));
  nand2 gate1158(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1159(.a(s_87), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1160(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1161(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1162(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1821(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1822(.a(gate431inter0), .b(s_182), .O(gate431inter1));
  and2  gate1823(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1824(.a(s_182), .O(gate431inter3));
  inv1  gate1825(.a(s_183), .O(gate431inter4));
  nand2 gate1826(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1827(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1828(.a(G7), .O(gate431inter7));
  inv1  gate1829(.a(G1150), .O(gate431inter8));
  nand2 gate1830(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1831(.a(s_183), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1832(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1833(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1834(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1877(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1878(.a(gate432inter0), .b(s_190), .O(gate432inter1));
  and2  gate1879(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1880(.a(s_190), .O(gate432inter3));
  inv1  gate1881(.a(s_191), .O(gate432inter4));
  nand2 gate1882(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1883(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1884(.a(G1054), .O(gate432inter7));
  inv1  gate1885(.a(G1150), .O(gate432inter8));
  nand2 gate1886(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1887(.a(s_191), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1888(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1889(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1890(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1555(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1556(.a(gate434inter0), .b(s_144), .O(gate434inter1));
  and2  gate1557(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1558(.a(s_144), .O(gate434inter3));
  inv1  gate1559(.a(s_145), .O(gate434inter4));
  nand2 gate1560(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1561(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1562(.a(G1057), .O(gate434inter7));
  inv1  gate1563(.a(G1153), .O(gate434inter8));
  nand2 gate1564(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1565(.a(s_145), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1566(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1567(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1568(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate2017(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2018(.a(gate437inter0), .b(s_210), .O(gate437inter1));
  and2  gate2019(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2020(.a(s_210), .O(gate437inter3));
  inv1  gate2021(.a(s_211), .O(gate437inter4));
  nand2 gate2022(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2023(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2024(.a(G10), .O(gate437inter7));
  inv1  gate2025(.a(G1159), .O(gate437inter8));
  nand2 gate2026(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2027(.a(s_211), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2028(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2029(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2030(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate785(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate786(.a(gate439inter0), .b(s_34), .O(gate439inter1));
  and2  gate787(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate788(.a(s_34), .O(gate439inter3));
  inv1  gate789(.a(s_35), .O(gate439inter4));
  nand2 gate790(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate791(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate792(.a(G11), .O(gate439inter7));
  inv1  gate793(.a(G1162), .O(gate439inter8));
  nand2 gate794(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate795(.a(s_35), .b(gate439inter3), .O(gate439inter10));
  nor2  gate796(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate797(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate798(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1079(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1080(.a(gate440inter0), .b(s_76), .O(gate440inter1));
  and2  gate1081(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1082(.a(s_76), .O(gate440inter3));
  inv1  gate1083(.a(s_77), .O(gate440inter4));
  nand2 gate1084(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1085(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1086(.a(G1066), .O(gate440inter7));
  inv1  gate1087(.a(G1162), .O(gate440inter8));
  nand2 gate1088(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1089(.a(s_77), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1090(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1091(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1092(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2031(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2032(.a(gate442inter0), .b(s_212), .O(gate442inter1));
  and2  gate2033(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2034(.a(s_212), .O(gate442inter3));
  inv1  gate2035(.a(s_213), .O(gate442inter4));
  nand2 gate2036(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2037(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2038(.a(G1069), .O(gate442inter7));
  inv1  gate2039(.a(G1165), .O(gate442inter8));
  nand2 gate2040(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2041(.a(s_213), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2042(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2043(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2044(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2059(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2060(.a(gate444inter0), .b(s_216), .O(gate444inter1));
  and2  gate2061(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2062(.a(s_216), .O(gate444inter3));
  inv1  gate2063(.a(s_217), .O(gate444inter4));
  nand2 gate2064(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2065(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2066(.a(G1072), .O(gate444inter7));
  inv1  gate2067(.a(G1168), .O(gate444inter8));
  nand2 gate2068(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2069(.a(s_217), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2070(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2071(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2072(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1107(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1108(.a(gate449inter0), .b(s_80), .O(gate449inter1));
  and2  gate1109(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1110(.a(s_80), .O(gate449inter3));
  inv1  gate1111(.a(s_81), .O(gate449inter4));
  nand2 gate1112(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1113(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1114(.a(G16), .O(gate449inter7));
  inv1  gate1115(.a(G1177), .O(gate449inter8));
  nand2 gate1116(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1117(.a(s_81), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1118(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1119(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1120(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1891(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1892(.a(gate451inter0), .b(s_192), .O(gate451inter1));
  and2  gate1893(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1894(.a(s_192), .O(gate451inter3));
  inv1  gate1895(.a(s_193), .O(gate451inter4));
  nand2 gate1896(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1897(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1898(.a(G17), .O(gate451inter7));
  inv1  gate1899(.a(G1180), .O(gate451inter8));
  nand2 gate1900(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1901(.a(s_193), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1902(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1903(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1904(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1471(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1472(.a(gate460inter0), .b(s_132), .O(gate460inter1));
  and2  gate1473(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1474(.a(s_132), .O(gate460inter3));
  inv1  gate1475(.a(s_133), .O(gate460inter4));
  nand2 gate1476(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1477(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1478(.a(G1096), .O(gate460inter7));
  inv1  gate1479(.a(G1192), .O(gate460inter8));
  nand2 gate1480(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1481(.a(s_133), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1482(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1483(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1484(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate897(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate898(.a(gate463inter0), .b(s_50), .O(gate463inter1));
  and2  gate899(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate900(.a(s_50), .O(gate463inter3));
  inv1  gate901(.a(s_51), .O(gate463inter4));
  nand2 gate902(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate903(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate904(.a(G23), .O(gate463inter7));
  inv1  gate905(.a(G1198), .O(gate463inter8));
  nand2 gate906(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate907(.a(s_51), .b(gate463inter3), .O(gate463inter10));
  nor2  gate908(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate909(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate910(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1961(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1962(.a(gate466inter0), .b(s_202), .O(gate466inter1));
  and2  gate1963(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1964(.a(s_202), .O(gate466inter3));
  inv1  gate1965(.a(s_203), .O(gate466inter4));
  nand2 gate1966(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1967(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1968(.a(G1105), .O(gate466inter7));
  inv1  gate1969(.a(G1201), .O(gate466inter8));
  nand2 gate1970(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1971(.a(s_203), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1972(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1973(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1974(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1933(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1934(.a(gate469inter0), .b(s_198), .O(gate469inter1));
  and2  gate1935(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1936(.a(s_198), .O(gate469inter3));
  inv1  gate1937(.a(s_199), .O(gate469inter4));
  nand2 gate1938(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1939(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1940(.a(G26), .O(gate469inter7));
  inv1  gate1941(.a(G1207), .O(gate469inter8));
  nand2 gate1942(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1943(.a(s_199), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1944(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1945(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1946(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1863(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1864(.a(gate471inter0), .b(s_188), .O(gate471inter1));
  and2  gate1865(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1866(.a(s_188), .O(gate471inter3));
  inv1  gate1867(.a(s_189), .O(gate471inter4));
  nand2 gate1868(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1869(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1870(.a(G27), .O(gate471inter7));
  inv1  gate1871(.a(G1210), .O(gate471inter8));
  nand2 gate1872(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1873(.a(s_189), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1874(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1875(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1876(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1625(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1626(.a(gate477inter0), .b(s_154), .O(gate477inter1));
  and2  gate1627(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1628(.a(s_154), .O(gate477inter3));
  inv1  gate1629(.a(s_155), .O(gate477inter4));
  nand2 gate1630(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1631(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1632(.a(G30), .O(gate477inter7));
  inv1  gate1633(.a(G1219), .O(gate477inter8));
  nand2 gate1634(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1635(.a(s_155), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1636(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1637(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1638(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate701(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate702(.a(gate478inter0), .b(s_22), .O(gate478inter1));
  and2  gate703(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate704(.a(s_22), .O(gate478inter3));
  inv1  gate705(.a(s_23), .O(gate478inter4));
  nand2 gate706(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate707(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate708(.a(G1123), .O(gate478inter7));
  inv1  gate709(.a(G1219), .O(gate478inter8));
  nand2 gate710(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate711(.a(s_23), .b(gate478inter3), .O(gate478inter10));
  nor2  gate712(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate713(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate714(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1121(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1122(.a(gate500inter0), .b(s_82), .O(gate500inter1));
  and2  gate1123(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1124(.a(s_82), .O(gate500inter3));
  inv1  gate1125(.a(s_83), .O(gate500inter4));
  nand2 gate1126(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1127(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1128(.a(G1262), .O(gate500inter7));
  inv1  gate1129(.a(G1263), .O(gate500inter8));
  nand2 gate1130(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1131(.a(s_83), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1132(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1133(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1134(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1793(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1794(.a(gate501inter0), .b(s_178), .O(gate501inter1));
  and2  gate1795(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1796(.a(s_178), .O(gate501inter3));
  inv1  gate1797(.a(s_179), .O(gate501inter4));
  nand2 gate1798(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1799(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1800(.a(G1264), .O(gate501inter7));
  inv1  gate1801(.a(G1265), .O(gate501inter8));
  nand2 gate1802(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1803(.a(s_179), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1804(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1805(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1806(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1499(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1500(.a(gate503inter0), .b(s_136), .O(gate503inter1));
  and2  gate1501(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1502(.a(s_136), .O(gate503inter3));
  inv1  gate1503(.a(s_137), .O(gate503inter4));
  nand2 gate1504(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1505(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1506(.a(G1268), .O(gate503inter7));
  inv1  gate1507(.a(G1269), .O(gate503inter8));
  nand2 gate1508(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1509(.a(s_137), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1510(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1511(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1512(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1177(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1178(.a(gate508inter0), .b(s_90), .O(gate508inter1));
  and2  gate1179(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1180(.a(s_90), .O(gate508inter3));
  inv1  gate1181(.a(s_91), .O(gate508inter4));
  nand2 gate1182(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1183(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1184(.a(G1278), .O(gate508inter7));
  inv1  gate1185(.a(G1279), .O(gate508inter8));
  nand2 gate1186(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1187(.a(s_91), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1188(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1189(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1190(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2115(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2116(.a(gate511inter0), .b(s_224), .O(gate511inter1));
  and2  gate2117(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2118(.a(s_224), .O(gate511inter3));
  inv1  gate2119(.a(s_225), .O(gate511inter4));
  nand2 gate2120(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2121(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2122(.a(G1284), .O(gate511inter7));
  inv1  gate2123(.a(G1285), .O(gate511inter8));
  nand2 gate2124(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2125(.a(s_225), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2126(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2127(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2128(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1667(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1668(.a(gate512inter0), .b(s_160), .O(gate512inter1));
  and2  gate1669(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1670(.a(s_160), .O(gate512inter3));
  inv1  gate1671(.a(s_161), .O(gate512inter4));
  nand2 gate1672(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1673(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1674(.a(G1286), .O(gate512inter7));
  inv1  gate1675(.a(G1287), .O(gate512inter8));
  nand2 gate1676(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1677(.a(s_161), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1678(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1679(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1680(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule