module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1485(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1486(.a(gate11inter0), .b(s_134), .O(gate11inter1));
  and2  gate1487(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1488(.a(s_134), .O(gate11inter3));
  inv1  gate1489(.a(s_135), .O(gate11inter4));
  nand2 gate1490(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1491(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1492(.a(G5), .O(gate11inter7));
  inv1  gate1493(.a(G6), .O(gate11inter8));
  nand2 gate1494(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1495(.a(s_135), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1496(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1497(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1498(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1975(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1976(.a(gate12inter0), .b(s_204), .O(gate12inter1));
  and2  gate1977(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1978(.a(s_204), .O(gate12inter3));
  inv1  gate1979(.a(s_205), .O(gate12inter4));
  nand2 gate1980(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1981(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1982(.a(G7), .O(gate12inter7));
  inv1  gate1983(.a(G8), .O(gate12inter8));
  nand2 gate1984(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1985(.a(s_205), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1986(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1987(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1988(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2381(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2382(.a(gate13inter0), .b(s_262), .O(gate13inter1));
  and2  gate2383(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2384(.a(s_262), .O(gate13inter3));
  inv1  gate2385(.a(s_263), .O(gate13inter4));
  nand2 gate2386(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2387(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2388(.a(G9), .O(gate13inter7));
  inv1  gate2389(.a(G10), .O(gate13inter8));
  nand2 gate2390(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2391(.a(s_263), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2392(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2393(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2394(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1331(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1332(.a(gate14inter0), .b(s_112), .O(gate14inter1));
  and2  gate1333(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1334(.a(s_112), .O(gate14inter3));
  inv1  gate1335(.a(s_113), .O(gate14inter4));
  nand2 gate1336(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1337(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1338(.a(G11), .O(gate14inter7));
  inv1  gate1339(.a(G12), .O(gate14inter8));
  nand2 gate1340(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1341(.a(s_113), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1342(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1343(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1344(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1779(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1780(.a(gate16inter0), .b(s_176), .O(gate16inter1));
  and2  gate1781(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1782(.a(s_176), .O(gate16inter3));
  inv1  gate1783(.a(s_177), .O(gate16inter4));
  nand2 gate1784(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1785(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1786(.a(G15), .O(gate16inter7));
  inv1  gate1787(.a(G16), .O(gate16inter8));
  nand2 gate1788(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1789(.a(s_177), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1790(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1791(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1792(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1919(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1920(.a(gate21inter0), .b(s_196), .O(gate21inter1));
  and2  gate1921(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1922(.a(s_196), .O(gate21inter3));
  inv1  gate1923(.a(s_197), .O(gate21inter4));
  nand2 gate1924(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1925(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1926(.a(G25), .O(gate21inter7));
  inv1  gate1927(.a(G26), .O(gate21inter8));
  nand2 gate1928(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1929(.a(s_197), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1930(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1931(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1932(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate911(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate912(.a(gate25inter0), .b(s_52), .O(gate25inter1));
  and2  gate913(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate914(.a(s_52), .O(gate25inter3));
  inv1  gate915(.a(s_53), .O(gate25inter4));
  nand2 gate916(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate917(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate918(.a(G1), .O(gate25inter7));
  inv1  gate919(.a(G5), .O(gate25inter8));
  nand2 gate920(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate921(.a(s_53), .b(gate25inter3), .O(gate25inter10));
  nor2  gate922(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate923(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate924(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2059(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2060(.a(gate27inter0), .b(s_216), .O(gate27inter1));
  and2  gate2061(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2062(.a(s_216), .O(gate27inter3));
  inv1  gate2063(.a(s_217), .O(gate27inter4));
  nand2 gate2064(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2065(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2066(.a(G2), .O(gate27inter7));
  inv1  gate2067(.a(G6), .O(gate27inter8));
  nand2 gate2068(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2069(.a(s_217), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2070(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2071(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2072(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate883(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate884(.a(gate29inter0), .b(s_48), .O(gate29inter1));
  and2  gate885(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate886(.a(s_48), .O(gate29inter3));
  inv1  gate887(.a(s_49), .O(gate29inter4));
  nand2 gate888(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate889(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate890(.a(G3), .O(gate29inter7));
  inv1  gate891(.a(G7), .O(gate29inter8));
  nand2 gate892(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate893(.a(s_49), .b(gate29inter3), .O(gate29inter10));
  nor2  gate894(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate895(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate896(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1541(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1542(.a(gate30inter0), .b(s_142), .O(gate30inter1));
  and2  gate1543(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1544(.a(s_142), .O(gate30inter3));
  inv1  gate1545(.a(s_143), .O(gate30inter4));
  nand2 gate1546(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1547(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1548(.a(G11), .O(gate30inter7));
  inv1  gate1549(.a(G15), .O(gate30inter8));
  nand2 gate1550(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1551(.a(s_143), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1552(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1553(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1554(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2227(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2228(.a(gate32inter0), .b(s_240), .O(gate32inter1));
  and2  gate2229(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2230(.a(s_240), .O(gate32inter3));
  inv1  gate2231(.a(s_241), .O(gate32inter4));
  nand2 gate2232(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2233(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2234(.a(G12), .O(gate32inter7));
  inv1  gate2235(.a(G16), .O(gate32inter8));
  nand2 gate2236(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2237(.a(s_241), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2238(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2239(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2240(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2199(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2200(.a(gate36inter0), .b(s_236), .O(gate36inter1));
  and2  gate2201(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2202(.a(s_236), .O(gate36inter3));
  inv1  gate2203(.a(s_237), .O(gate36inter4));
  nand2 gate2204(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2205(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2206(.a(G26), .O(gate36inter7));
  inv1  gate2207(.a(G30), .O(gate36inter8));
  nand2 gate2208(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2209(.a(s_237), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2210(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2211(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2212(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1275(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1276(.a(gate37inter0), .b(s_104), .O(gate37inter1));
  and2  gate1277(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1278(.a(s_104), .O(gate37inter3));
  inv1  gate1279(.a(s_105), .O(gate37inter4));
  nand2 gate1280(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1281(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1282(.a(G19), .O(gate37inter7));
  inv1  gate1283(.a(G23), .O(gate37inter8));
  nand2 gate1284(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1285(.a(s_105), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1286(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1287(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1288(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2395(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2396(.a(gate39inter0), .b(s_264), .O(gate39inter1));
  and2  gate2397(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2398(.a(s_264), .O(gate39inter3));
  inv1  gate2399(.a(s_265), .O(gate39inter4));
  nand2 gate2400(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2401(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2402(.a(G20), .O(gate39inter7));
  inv1  gate2403(.a(G24), .O(gate39inter8));
  nand2 gate2404(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2405(.a(s_265), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2406(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2407(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2408(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate757(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate758(.a(gate51inter0), .b(s_30), .O(gate51inter1));
  and2  gate759(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate760(.a(s_30), .O(gate51inter3));
  inv1  gate761(.a(s_31), .O(gate51inter4));
  nand2 gate762(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate763(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate764(.a(G11), .O(gate51inter7));
  inv1  gate765(.a(G281), .O(gate51inter8));
  nand2 gate766(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate767(.a(s_31), .b(gate51inter3), .O(gate51inter10));
  nor2  gate768(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate769(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate770(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate2409(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2410(.a(gate52inter0), .b(s_266), .O(gate52inter1));
  and2  gate2411(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2412(.a(s_266), .O(gate52inter3));
  inv1  gate2413(.a(s_267), .O(gate52inter4));
  nand2 gate2414(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2415(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2416(.a(G12), .O(gate52inter7));
  inv1  gate2417(.a(G281), .O(gate52inter8));
  nand2 gate2418(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2419(.a(s_267), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2420(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2421(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2422(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2185(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2186(.a(gate54inter0), .b(s_234), .O(gate54inter1));
  and2  gate2187(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2188(.a(s_234), .O(gate54inter3));
  inv1  gate2189(.a(s_235), .O(gate54inter4));
  nand2 gate2190(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2191(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2192(.a(G14), .O(gate54inter7));
  inv1  gate2193(.a(G284), .O(gate54inter8));
  nand2 gate2194(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2195(.a(s_235), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2196(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2197(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2198(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate2129(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2130(.a(gate55inter0), .b(s_226), .O(gate55inter1));
  and2  gate2131(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2132(.a(s_226), .O(gate55inter3));
  inv1  gate2133(.a(s_227), .O(gate55inter4));
  nand2 gate2134(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2135(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2136(.a(G15), .O(gate55inter7));
  inv1  gate2137(.a(G287), .O(gate55inter8));
  nand2 gate2138(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2139(.a(s_227), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2140(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2141(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2142(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1023(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1024(.a(gate58inter0), .b(s_68), .O(gate58inter1));
  and2  gate1025(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1026(.a(s_68), .O(gate58inter3));
  inv1  gate1027(.a(s_69), .O(gate58inter4));
  nand2 gate1028(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1029(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1030(.a(G18), .O(gate58inter7));
  inv1  gate1031(.a(G290), .O(gate58inter8));
  nand2 gate1032(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1033(.a(s_69), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1034(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1035(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1036(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate2017(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2018(.a(gate59inter0), .b(s_210), .O(gate59inter1));
  and2  gate2019(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2020(.a(s_210), .O(gate59inter3));
  inv1  gate2021(.a(s_211), .O(gate59inter4));
  nand2 gate2022(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2023(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2024(.a(G19), .O(gate59inter7));
  inv1  gate2025(.a(G293), .O(gate59inter8));
  nand2 gate2026(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2027(.a(s_211), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2028(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2029(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2030(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate645(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate646(.a(gate62inter0), .b(s_14), .O(gate62inter1));
  and2  gate647(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate648(.a(s_14), .O(gate62inter3));
  inv1  gate649(.a(s_15), .O(gate62inter4));
  nand2 gate650(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate651(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate652(.a(G22), .O(gate62inter7));
  inv1  gate653(.a(G296), .O(gate62inter8));
  nand2 gate654(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate655(.a(s_15), .b(gate62inter3), .O(gate62inter10));
  nor2  gate656(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate657(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate658(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate939(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate940(.a(gate63inter0), .b(s_56), .O(gate63inter1));
  and2  gate941(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate942(.a(s_56), .O(gate63inter3));
  inv1  gate943(.a(s_57), .O(gate63inter4));
  nand2 gate944(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate945(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate946(.a(G23), .O(gate63inter7));
  inv1  gate947(.a(G299), .O(gate63inter8));
  nand2 gate948(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate949(.a(s_57), .b(gate63inter3), .O(gate63inter10));
  nor2  gate950(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate951(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate952(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1681(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1682(.a(gate64inter0), .b(s_162), .O(gate64inter1));
  and2  gate1683(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1684(.a(s_162), .O(gate64inter3));
  inv1  gate1685(.a(s_163), .O(gate64inter4));
  nand2 gate1686(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1687(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1688(.a(G24), .O(gate64inter7));
  inv1  gate1689(.a(G299), .O(gate64inter8));
  nand2 gate1690(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1691(.a(s_163), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1692(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1693(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1694(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1639(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1640(.a(gate68inter0), .b(s_156), .O(gate68inter1));
  and2  gate1641(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1642(.a(s_156), .O(gate68inter3));
  inv1  gate1643(.a(s_157), .O(gate68inter4));
  nand2 gate1644(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1645(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1646(.a(G28), .O(gate68inter7));
  inv1  gate1647(.a(G305), .O(gate68inter8));
  nand2 gate1648(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1649(.a(s_157), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1650(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1651(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1652(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1695(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1696(.a(gate71inter0), .b(s_164), .O(gate71inter1));
  and2  gate1697(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1698(.a(s_164), .O(gate71inter3));
  inv1  gate1699(.a(s_165), .O(gate71inter4));
  nand2 gate1700(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1701(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1702(.a(G31), .O(gate71inter7));
  inv1  gate1703(.a(G311), .O(gate71inter8));
  nand2 gate1704(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1705(.a(s_165), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1706(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1707(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1708(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2283(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2284(.a(gate72inter0), .b(s_248), .O(gate72inter1));
  and2  gate2285(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2286(.a(s_248), .O(gate72inter3));
  inv1  gate2287(.a(s_249), .O(gate72inter4));
  nand2 gate2288(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2289(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2290(.a(G32), .O(gate72inter7));
  inv1  gate2291(.a(G311), .O(gate72inter8));
  nand2 gate2292(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2293(.a(s_249), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2294(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2295(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2296(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1877(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1878(.a(gate73inter0), .b(s_190), .O(gate73inter1));
  and2  gate1879(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1880(.a(s_190), .O(gate73inter3));
  inv1  gate1881(.a(s_191), .O(gate73inter4));
  nand2 gate1882(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1883(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1884(.a(G1), .O(gate73inter7));
  inv1  gate1885(.a(G314), .O(gate73inter8));
  nand2 gate1886(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1887(.a(s_191), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1888(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1889(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1890(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate995(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate996(.a(gate74inter0), .b(s_64), .O(gate74inter1));
  and2  gate997(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate998(.a(s_64), .O(gate74inter3));
  inv1  gate999(.a(s_65), .O(gate74inter4));
  nand2 gate1000(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1001(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1002(.a(G5), .O(gate74inter7));
  inv1  gate1003(.a(G314), .O(gate74inter8));
  nand2 gate1004(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1005(.a(s_65), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1006(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1007(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1008(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1177(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1178(.a(gate75inter0), .b(s_90), .O(gate75inter1));
  and2  gate1179(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1180(.a(s_90), .O(gate75inter3));
  inv1  gate1181(.a(s_91), .O(gate75inter4));
  nand2 gate1182(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1183(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1184(.a(G9), .O(gate75inter7));
  inv1  gate1185(.a(G317), .O(gate75inter8));
  nand2 gate1186(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1187(.a(s_91), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1188(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1189(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1190(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1373(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1374(.a(gate77inter0), .b(s_118), .O(gate77inter1));
  and2  gate1375(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1376(.a(s_118), .O(gate77inter3));
  inv1  gate1377(.a(s_119), .O(gate77inter4));
  nand2 gate1378(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1379(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1380(.a(G2), .O(gate77inter7));
  inv1  gate1381(.a(G320), .O(gate77inter8));
  nand2 gate1382(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1383(.a(s_119), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1384(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1385(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1386(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2297(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2298(.a(gate80inter0), .b(s_250), .O(gate80inter1));
  and2  gate2299(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2300(.a(s_250), .O(gate80inter3));
  inv1  gate2301(.a(s_251), .O(gate80inter4));
  nand2 gate2302(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2303(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2304(.a(G14), .O(gate80inter7));
  inv1  gate2305(.a(G323), .O(gate80inter8));
  nand2 gate2306(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2307(.a(s_251), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2308(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2309(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2310(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2045(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2046(.a(gate81inter0), .b(s_214), .O(gate81inter1));
  and2  gate2047(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2048(.a(s_214), .O(gate81inter3));
  inv1  gate2049(.a(s_215), .O(gate81inter4));
  nand2 gate2050(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2051(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2052(.a(G3), .O(gate81inter7));
  inv1  gate2053(.a(G326), .O(gate81inter8));
  nand2 gate2054(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2055(.a(s_215), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2056(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2057(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2058(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate841(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate842(.a(gate82inter0), .b(s_42), .O(gate82inter1));
  and2  gate843(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate844(.a(s_42), .O(gate82inter3));
  inv1  gate845(.a(s_43), .O(gate82inter4));
  nand2 gate846(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate847(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate848(.a(G7), .O(gate82inter7));
  inv1  gate849(.a(G326), .O(gate82inter8));
  nand2 gate850(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate851(.a(s_43), .b(gate82inter3), .O(gate82inter10));
  nor2  gate852(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate853(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate854(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2255(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2256(.a(gate85inter0), .b(s_244), .O(gate85inter1));
  and2  gate2257(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2258(.a(s_244), .O(gate85inter3));
  inv1  gate2259(.a(s_245), .O(gate85inter4));
  nand2 gate2260(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2261(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2262(.a(G4), .O(gate85inter7));
  inv1  gate2263(.a(G332), .O(gate85inter8));
  nand2 gate2264(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2265(.a(s_245), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2266(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2267(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2268(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1807(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1808(.a(gate88inter0), .b(s_180), .O(gate88inter1));
  and2  gate1809(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1810(.a(s_180), .O(gate88inter3));
  inv1  gate1811(.a(s_181), .O(gate88inter4));
  nand2 gate1812(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1813(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1814(.a(G16), .O(gate88inter7));
  inv1  gate1815(.a(G335), .O(gate88inter8));
  nand2 gate1816(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1817(.a(s_181), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1818(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1819(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1820(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate743(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate744(.a(gate90inter0), .b(s_28), .O(gate90inter1));
  and2  gate745(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate746(.a(s_28), .O(gate90inter3));
  inv1  gate747(.a(s_29), .O(gate90inter4));
  nand2 gate748(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate749(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate750(.a(G21), .O(gate90inter7));
  inv1  gate751(.a(G338), .O(gate90inter8));
  nand2 gate752(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate753(.a(s_29), .b(gate90inter3), .O(gate90inter10));
  nor2  gate754(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate755(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate756(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2143(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2144(.a(gate100inter0), .b(s_228), .O(gate100inter1));
  and2  gate2145(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2146(.a(s_228), .O(gate100inter3));
  inv1  gate2147(.a(s_229), .O(gate100inter4));
  nand2 gate2148(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2149(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2150(.a(G31), .O(gate100inter7));
  inv1  gate2151(.a(G353), .O(gate100inter8));
  nand2 gate2152(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2153(.a(s_229), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2154(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2155(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2156(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate2507(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2508(.a(gate101inter0), .b(s_280), .O(gate101inter1));
  and2  gate2509(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2510(.a(s_280), .O(gate101inter3));
  inv1  gate2511(.a(s_281), .O(gate101inter4));
  nand2 gate2512(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2513(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2514(.a(G20), .O(gate101inter7));
  inv1  gate2515(.a(G356), .O(gate101inter8));
  nand2 gate2516(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2517(.a(s_281), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2518(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2519(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2520(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1457(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1458(.a(gate104inter0), .b(s_130), .O(gate104inter1));
  and2  gate1459(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1460(.a(s_130), .O(gate104inter3));
  inv1  gate1461(.a(s_131), .O(gate104inter4));
  nand2 gate1462(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1463(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1464(.a(G32), .O(gate104inter7));
  inv1  gate1465(.a(G359), .O(gate104inter8));
  nand2 gate1466(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1467(.a(s_131), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1468(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1469(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1470(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate729(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate730(.a(gate109inter0), .b(s_26), .O(gate109inter1));
  and2  gate731(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate732(.a(s_26), .O(gate109inter3));
  inv1  gate733(.a(s_27), .O(gate109inter4));
  nand2 gate734(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate735(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate736(.a(G370), .O(gate109inter7));
  inv1  gate737(.a(G371), .O(gate109inter8));
  nand2 gate738(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate739(.a(s_27), .b(gate109inter3), .O(gate109inter10));
  nor2  gate740(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate741(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate742(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate2353(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2354(.a(gate110inter0), .b(s_258), .O(gate110inter1));
  and2  gate2355(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2356(.a(s_258), .O(gate110inter3));
  inv1  gate2357(.a(s_259), .O(gate110inter4));
  nand2 gate2358(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2359(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2360(.a(G372), .O(gate110inter7));
  inv1  gate2361(.a(G373), .O(gate110inter8));
  nand2 gate2362(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2363(.a(s_259), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2364(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2365(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2366(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2311(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2312(.a(gate111inter0), .b(s_252), .O(gate111inter1));
  and2  gate2313(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2314(.a(s_252), .O(gate111inter3));
  inv1  gate2315(.a(s_253), .O(gate111inter4));
  nand2 gate2316(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2317(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2318(.a(G374), .O(gate111inter7));
  inv1  gate2319(.a(G375), .O(gate111inter8));
  nand2 gate2320(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2321(.a(s_253), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2322(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2323(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2324(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate2339(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2340(.a(gate113inter0), .b(s_256), .O(gate113inter1));
  and2  gate2341(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2342(.a(s_256), .O(gate113inter3));
  inv1  gate2343(.a(s_257), .O(gate113inter4));
  nand2 gate2344(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2345(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2346(.a(G378), .O(gate113inter7));
  inv1  gate2347(.a(G379), .O(gate113inter8));
  nand2 gate2348(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2349(.a(s_257), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2350(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2351(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2352(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1135(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1136(.a(gate116inter0), .b(s_84), .O(gate116inter1));
  and2  gate1137(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1138(.a(s_84), .O(gate116inter3));
  inv1  gate1139(.a(s_85), .O(gate116inter4));
  nand2 gate1140(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1141(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1142(.a(G384), .O(gate116inter7));
  inv1  gate1143(.a(G385), .O(gate116inter8));
  nand2 gate1144(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1145(.a(s_85), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1146(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1147(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1148(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2437(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2438(.a(gate121inter0), .b(s_270), .O(gate121inter1));
  and2  gate2439(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2440(.a(s_270), .O(gate121inter3));
  inv1  gate2441(.a(s_271), .O(gate121inter4));
  nand2 gate2442(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2443(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2444(.a(G394), .O(gate121inter7));
  inv1  gate2445(.a(G395), .O(gate121inter8));
  nand2 gate2446(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2447(.a(s_271), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2448(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2449(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2450(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1835(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1836(.a(gate123inter0), .b(s_184), .O(gate123inter1));
  and2  gate1837(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1838(.a(s_184), .O(gate123inter3));
  inv1  gate1839(.a(s_185), .O(gate123inter4));
  nand2 gate1840(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1841(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1842(.a(G398), .O(gate123inter7));
  inv1  gate1843(.a(G399), .O(gate123inter8));
  nand2 gate1844(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1845(.a(s_185), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1846(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1847(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1848(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate785(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate786(.a(gate124inter0), .b(s_34), .O(gate124inter1));
  and2  gate787(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate788(.a(s_34), .O(gate124inter3));
  inv1  gate789(.a(s_35), .O(gate124inter4));
  nand2 gate790(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate791(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate792(.a(G400), .O(gate124inter7));
  inv1  gate793(.a(G401), .O(gate124inter8));
  nand2 gate794(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate795(.a(s_35), .b(gate124inter3), .O(gate124inter10));
  nor2  gate796(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate797(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate798(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate631(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate632(.a(gate125inter0), .b(s_12), .O(gate125inter1));
  and2  gate633(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate634(.a(s_12), .O(gate125inter3));
  inv1  gate635(.a(s_13), .O(gate125inter4));
  nand2 gate636(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate637(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate638(.a(G402), .O(gate125inter7));
  inv1  gate639(.a(G403), .O(gate125inter8));
  nand2 gate640(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate641(.a(s_13), .b(gate125inter3), .O(gate125inter10));
  nor2  gate642(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate643(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate644(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1905(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1906(.a(gate129inter0), .b(s_194), .O(gate129inter1));
  and2  gate1907(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1908(.a(s_194), .O(gate129inter3));
  inv1  gate1909(.a(s_195), .O(gate129inter4));
  nand2 gate1910(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1911(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1912(.a(G410), .O(gate129inter7));
  inv1  gate1913(.a(G411), .O(gate129inter8));
  nand2 gate1914(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1915(.a(s_195), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1916(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1917(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1918(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate855(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate856(.a(gate133inter0), .b(s_44), .O(gate133inter1));
  and2  gate857(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate858(.a(s_44), .O(gate133inter3));
  inv1  gate859(.a(s_45), .O(gate133inter4));
  nand2 gate860(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate861(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate862(.a(G418), .O(gate133inter7));
  inv1  gate863(.a(G419), .O(gate133inter8));
  nand2 gate864(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate865(.a(s_45), .b(gate133inter3), .O(gate133inter10));
  nor2  gate866(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate867(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate868(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate981(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate982(.a(gate134inter0), .b(s_62), .O(gate134inter1));
  and2  gate983(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate984(.a(s_62), .O(gate134inter3));
  inv1  gate985(.a(s_63), .O(gate134inter4));
  nand2 gate986(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate987(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate988(.a(G420), .O(gate134inter7));
  inv1  gate989(.a(G421), .O(gate134inter8));
  nand2 gate990(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate991(.a(s_63), .b(gate134inter3), .O(gate134inter10));
  nor2  gate992(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate993(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate994(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2451(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2452(.a(gate143inter0), .b(s_272), .O(gate143inter1));
  and2  gate2453(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2454(.a(s_272), .O(gate143inter3));
  inv1  gate2455(.a(s_273), .O(gate143inter4));
  nand2 gate2456(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2457(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2458(.a(G462), .O(gate143inter7));
  inv1  gate2459(.a(G465), .O(gate143inter8));
  nand2 gate2460(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2461(.a(s_273), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2462(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2463(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2464(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1961(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1962(.a(gate144inter0), .b(s_202), .O(gate144inter1));
  and2  gate1963(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1964(.a(s_202), .O(gate144inter3));
  inv1  gate1965(.a(s_203), .O(gate144inter4));
  nand2 gate1966(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1967(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1968(.a(G468), .O(gate144inter7));
  inv1  gate1969(.a(G471), .O(gate144inter8));
  nand2 gate1970(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1971(.a(s_203), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1972(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1973(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1974(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1247(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1248(.a(gate146inter0), .b(s_100), .O(gate146inter1));
  and2  gate1249(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1250(.a(s_100), .O(gate146inter3));
  inv1  gate1251(.a(s_101), .O(gate146inter4));
  nand2 gate1252(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1253(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1254(.a(G480), .O(gate146inter7));
  inv1  gate1255(.a(G483), .O(gate146inter8));
  nand2 gate1256(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1257(.a(s_101), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1258(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1259(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1260(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1163(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1164(.a(gate148inter0), .b(s_88), .O(gate148inter1));
  and2  gate1165(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1166(.a(s_88), .O(gate148inter3));
  inv1  gate1167(.a(s_89), .O(gate148inter4));
  nand2 gate1168(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1169(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1170(.a(G492), .O(gate148inter7));
  inv1  gate1171(.a(G495), .O(gate148inter8));
  nand2 gate1172(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1173(.a(s_89), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1174(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1175(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1176(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1499(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1500(.a(gate150inter0), .b(s_136), .O(gate150inter1));
  and2  gate1501(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1502(.a(s_136), .O(gate150inter3));
  inv1  gate1503(.a(s_137), .O(gate150inter4));
  nand2 gate1504(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1505(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1506(.a(G504), .O(gate150inter7));
  inv1  gate1507(.a(G507), .O(gate150inter8));
  nand2 gate1508(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1509(.a(s_137), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1510(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1511(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1512(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2213(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2214(.a(gate151inter0), .b(s_238), .O(gate151inter1));
  and2  gate2215(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2216(.a(s_238), .O(gate151inter3));
  inv1  gate2217(.a(s_239), .O(gate151inter4));
  nand2 gate2218(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2219(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2220(.a(G510), .O(gate151inter7));
  inv1  gate2221(.a(G513), .O(gate151inter8));
  nand2 gate2222(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2223(.a(s_239), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2224(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2225(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2226(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate701(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate702(.a(gate152inter0), .b(s_22), .O(gate152inter1));
  and2  gate703(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate704(.a(s_22), .O(gate152inter3));
  inv1  gate705(.a(s_23), .O(gate152inter4));
  nand2 gate706(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate707(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate708(.a(G516), .O(gate152inter7));
  inv1  gate709(.a(G519), .O(gate152inter8));
  nand2 gate710(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate711(.a(s_23), .b(gate152inter3), .O(gate152inter10));
  nor2  gate712(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate713(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate714(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate561(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate562(.a(gate157inter0), .b(s_2), .O(gate157inter1));
  and2  gate563(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate564(.a(s_2), .O(gate157inter3));
  inv1  gate565(.a(s_3), .O(gate157inter4));
  nand2 gate566(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate567(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate568(.a(G438), .O(gate157inter7));
  inv1  gate569(.a(G528), .O(gate157inter8));
  nand2 gate570(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate571(.a(s_3), .b(gate157inter3), .O(gate157inter10));
  nor2  gate572(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate573(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate574(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1219(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1220(.a(gate158inter0), .b(s_96), .O(gate158inter1));
  and2  gate1221(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1222(.a(s_96), .O(gate158inter3));
  inv1  gate1223(.a(s_97), .O(gate158inter4));
  nand2 gate1224(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1225(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1226(.a(G441), .O(gate158inter7));
  inv1  gate1227(.a(G528), .O(gate158inter8));
  nand2 gate1228(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1229(.a(s_97), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1230(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1231(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1232(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1429(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1430(.a(gate159inter0), .b(s_126), .O(gate159inter1));
  and2  gate1431(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1432(.a(s_126), .O(gate159inter3));
  inv1  gate1433(.a(s_127), .O(gate159inter4));
  nand2 gate1434(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1435(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1436(.a(G444), .O(gate159inter7));
  inv1  gate1437(.a(G531), .O(gate159inter8));
  nand2 gate1438(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1439(.a(s_127), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1440(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1441(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1442(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2031(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2032(.a(gate165inter0), .b(s_212), .O(gate165inter1));
  and2  gate2033(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2034(.a(s_212), .O(gate165inter3));
  inv1  gate2035(.a(s_213), .O(gate165inter4));
  nand2 gate2036(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2037(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2038(.a(G462), .O(gate165inter7));
  inv1  gate2039(.a(G540), .O(gate165inter8));
  nand2 gate2040(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2041(.a(s_213), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2042(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2043(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2044(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2367(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2368(.a(gate170inter0), .b(s_260), .O(gate170inter1));
  and2  gate2369(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2370(.a(s_260), .O(gate170inter3));
  inv1  gate2371(.a(s_261), .O(gate170inter4));
  nand2 gate2372(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2373(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2374(.a(G477), .O(gate170inter7));
  inv1  gate2375(.a(G546), .O(gate170inter8));
  nand2 gate2376(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2377(.a(s_261), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2378(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2379(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2380(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1471(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1472(.a(gate171inter0), .b(s_132), .O(gate171inter1));
  and2  gate1473(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1474(.a(s_132), .O(gate171inter3));
  inv1  gate1475(.a(s_133), .O(gate171inter4));
  nand2 gate1476(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1477(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1478(.a(G480), .O(gate171inter7));
  inv1  gate1479(.a(G549), .O(gate171inter8));
  nand2 gate1480(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1481(.a(s_133), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1482(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1483(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1484(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2073(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2074(.a(gate173inter0), .b(s_218), .O(gate173inter1));
  and2  gate2075(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2076(.a(s_218), .O(gate173inter3));
  inv1  gate2077(.a(s_219), .O(gate173inter4));
  nand2 gate2078(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2079(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2080(.a(G486), .O(gate173inter7));
  inv1  gate2081(.a(G552), .O(gate173inter8));
  nand2 gate2082(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2083(.a(s_219), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2084(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2085(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2086(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2101(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2102(.a(gate174inter0), .b(s_222), .O(gate174inter1));
  and2  gate2103(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2104(.a(s_222), .O(gate174inter3));
  inv1  gate2105(.a(s_223), .O(gate174inter4));
  nand2 gate2106(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2107(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2108(.a(G489), .O(gate174inter7));
  inv1  gate2109(.a(G552), .O(gate174inter8));
  nand2 gate2110(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2111(.a(s_223), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2112(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2113(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2114(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1107(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1108(.a(gate176inter0), .b(s_80), .O(gate176inter1));
  and2  gate1109(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1110(.a(s_80), .O(gate176inter3));
  inv1  gate1111(.a(s_81), .O(gate176inter4));
  nand2 gate1112(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1113(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1114(.a(G495), .O(gate176inter7));
  inv1  gate1115(.a(G555), .O(gate176inter8));
  nand2 gate1116(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1117(.a(s_81), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1118(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1119(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1120(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1009(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1010(.a(gate179inter0), .b(s_66), .O(gate179inter1));
  and2  gate1011(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1012(.a(s_66), .O(gate179inter3));
  inv1  gate1013(.a(s_67), .O(gate179inter4));
  nand2 gate1014(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1015(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1016(.a(G504), .O(gate179inter7));
  inv1  gate1017(.a(G561), .O(gate179inter8));
  nand2 gate1018(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1019(.a(s_67), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1020(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1021(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1022(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate771(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate772(.a(gate181inter0), .b(s_32), .O(gate181inter1));
  and2  gate773(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate774(.a(s_32), .O(gate181inter3));
  inv1  gate775(.a(s_33), .O(gate181inter4));
  nand2 gate776(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate777(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate778(.a(G510), .O(gate181inter7));
  inv1  gate779(.a(G564), .O(gate181inter8));
  nand2 gate780(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate781(.a(s_33), .b(gate181inter3), .O(gate181inter10));
  nor2  gate782(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate783(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate784(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1555(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1556(.a(gate183inter0), .b(s_144), .O(gate183inter1));
  and2  gate1557(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1558(.a(s_144), .O(gate183inter3));
  inv1  gate1559(.a(s_145), .O(gate183inter4));
  nand2 gate1560(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1561(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1562(.a(G516), .O(gate183inter7));
  inv1  gate1563(.a(G567), .O(gate183inter8));
  nand2 gate1564(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1565(.a(s_145), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1566(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1567(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1568(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1611(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1612(.a(gate186inter0), .b(s_152), .O(gate186inter1));
  and2  gate1613(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1614(.a(s_152), .O(gate186inter3));
  inv1  gate1615(.a(s_153), .O(gate186inter4));
  nand2 gate1616(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1617(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1618(.a(G572), .O(gate186inter7));
  inv1  gate1619(.a(G573), .O(gate186inter8));
  nand2 gate1620(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1621(.a(s_153), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1622(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1623(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1624(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate603(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate604(.a(gate188inter0), .b(s_8), .O(gate188inter1));
  and2  gate605(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate606(.a(s_8), .O(gate188inter3));
  inv1  gate607(.a(s_9), .O(gate188inter4));
  nand2 gate608(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate609(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate610(.a(G576), .O(gate188inter7));
  inv1  gate611(.a(G577), .O(gate188inter8));
  nand2 gate612(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate613(.a(s_9), .b(gate188inter3), .O(gate188inter10));
  nor2  gate614(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate615(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate616(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate547(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate548(.a(gate191inter0), .b(s_0), .O(gate191inter1));
  and2  gate549(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate550(.a(s_0), .O(gate191inter3));
  inv1  gate551(.a(s_1), .O(gate191inter4));
  nand2 gate552(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate553(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate554(.a(G582), .O(gate191inter7));
  inv1  gate555(.a(G583), .O(gate191inter8));
  nand2 gate556(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate557(.a(s_1), .b(gate191inter3), .O(gate191inter10));
  nor2  gate558(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate559(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate560(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2493(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2494(.a(gate194inter0), .b(s_278), .O(gate194inter1));
  and2  gate2495(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2496(.a(s_278), .O(gate194inter3));
  inv1  gate2497(.a(s_279), .O(gate194inter4));
  nand2 gate2498(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2499(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2500(.a(G588), .O(gate194inter7));
  inv1  gate2501(.a(G589), .O(gate194inter8));
  nand2 gate2502(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2503(.a(s_279), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2504(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2505(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2506(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1289(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1290(.a(gate195inter0), .b(s_106), .O(gate195inter1));
  and2  gate1291(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1292(.a(s_106), .O(gate195inter3));
  inv1  gate1293(.a(s_107), .O(gate195inter4));
  nand2 gate1294(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1295(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1296(.a(G590), .O(gate195inter7));
  inv1  gate1297(.a(G591), .O(gate195inter8));
  nand2 gate1298(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1299(.a(s_107), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1300(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1301(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1302(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1821(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1822(.a(gate197inter0), .b(s_182), .O(gate197inter1));
  and2  gate1823(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1824(.a(s_182), .O(gate197inter3));
  inv1  gate1825(.a(s_183), .O(gate197inter4));
  nand2 gate1826(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1827(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1828(.a(G594), .O(gate197inter7));
  inv1  gate1829(.a(G595), .O(gate197inter8));
  nand2 gate1830(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1831(.a(s_183), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1832(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1833(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1834(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate659(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate660(.a(gate203inter0), .b(s_16), .O(gate203inter1));
  and2  gate661(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate662(.a(s_16), .O(gate203inter3));
  inv1  gate663(.a(s_17), .O(gate203inter4));
  nand2 gate664(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate665(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate666(.a(G602), .O(gate203inter7));
  inv1  gate667(.a(G612), .O(gate203inter8));
  nand2 gate668(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate669(.a(s_17), .b(gate203inter3), .O(gate203inter10));
  nor2  gate670(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate671(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate672(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2241(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2242(.a(gate206inter0), .b(s_242), .O(gate206inter1));
  and2  gate2243(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2244(.a(s_242), .O(gate206inter3));
  inv1  gate2245(.a(s_243), .O(gate206inter4));
  nand2 gate2246(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2247(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2248(.a(G632), .O(gate206inter7));
  inv1  gate2249(.a(G637), .O(gate206inter8));
  nand2 gate2250(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2251(.a(s_243), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2252(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2253(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2254(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1751(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1752(.a(gate211inter0), .b(s_172), .O(gate211inter1));
  and2  gate1753(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1754(.a(s_172), .O(gate211inter3));
  inv1  gate1755(.a(s_173), .O(gate211inter4));
  nand2 gate1756(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1757(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1758(.a(G612), .O(gate211inter7));
  inv1  gate1759(.a(G669), .O(gate211inter8));
  nand2 gate1760(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1761(.a(s_173), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1762(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1763(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1764(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate715(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate716(.a(gate214inter0), .b(s_24), .O(gate214inter1));
  and2  gate717(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate718(.a(s_24), .O(gate214inter3));
  inv1  gate719(.a(s_25), .O(gate214inter4));
  nand2 gate720(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate721(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate722(.a(G612), .O(gate214inter7));
  inv1  gate723(.a(G672), .O(gate214inter8));
  nand2 gate724(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate725(.a(s_25), .b(gate214inter3), .O(gate214inter10));
  nor2  gate726(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate727(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate728(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1625(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1626(.a(gate215inter0), .b(s_154), .O(gate215inter1));
  and2  gate1627(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1628(.a(s_154), .O(gate215inter3));
  inv1  gate1629(.a(s_155), .O(gate215inter4));
  nand2 gate1630(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1631(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1632(.a(G607), .O(gate215inter7));
  inv1  gate1633(.a(G675), .O(gate215inter8));
  nand2 gate1634(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1635(.a(s_155), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1636(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1637(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1638(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1793(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1794(.a(gate221inter0), .b(s_178), .O(gate221inter1));
  and2  gate1795(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1796(.a(s_178), .O(gate221inter3));
  inv1  gate1797(.a(s_179), .O(gate221inter4));
  nand2 gate1798(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1799(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1800(.a(G622), .O(gate221inter7));
  inv1  gate1801(.a(G684), .O(gate221inter8));
  nand2 gate1802(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1803(.a(s_179), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1804(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1805(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1806(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1303(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1304(.a(gate226inter0), .b(s_108), .O(gate226inter1));
  and2  gate1305(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1306(.a(s_108), .O(gate226inter3));
  inv1  gate1307(.a(s_109), .O(gate226inter4));
  nand2 gate1308(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1309(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1310(.a(G692), .O(gate226inter7));
  inv1  gate1311(.a(G693), .O(gate226inter8));
  nand2 gate1312(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1313(.a(s_109), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1314(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1315(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1316(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1233(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1234(.a(gate231inter0), .b(s_98), .O(gate231inter1));
  and2  gate1235(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1236(.a(s_98), .O(gate231inter3));
  inv1  gate1237(.a(s_99), .O(gate231inter4));
  nand2 gate1238(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1239(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1240(.a(G702), .O(gate231inter7));
  inv1  gate1241(.a(G703), .O(gate231inter8));
  nand2 gate1242(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1243(.a(s_99), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1244(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1245(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1246(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1765(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1766(.a(gate233inter0), .b(s_174), .O(gate233inter1));
  and2  gate1767(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1768(.a(s_174), .O(gate233inter3));
  inv1  gate1769(.a(s_175), .O(gate233inter4));
  nand2 gate1770(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1771(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1772(.a(G242), .O(gate233inter7));
  inv1  gate1773(.a(G718), .O(gate233inter8));
  nand2 gate1774(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1775(.a(s_175), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1776(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1777(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1778(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1261(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1262(.a(gate237inter0), .b(s_102), .O(gate237inter1));
  and2  gate1263(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1264(.a(s_102), .O(gate237inter3));
  inv1  gate1265(.a(s_103), .O(gate237inter4));
  nand2 gate1266(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1267(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1268(.a(G254), .O(gate237inter7));
  inv1  gate1269(.a(G706), .O(gate237inter8));
  nand2 gate1270(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1271(.a(s_103), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1272(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1273(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1274(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1051(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1052(.a(gate238inter0), .b(s_72), .O(gate238inter1));
  and2  gate1053(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1054(.a(s_72), .O(gate238inter3));
  inv1  gate1055(.a(s_73), .O(gate238inter4));
  nand2 gate1056(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1057(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1058(.a(G257), .O(gate238inter7));
  inv1  gate1059(.a(G709), .O(gate238inter8));
  nand2 gate1060(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1061(.a(s_73), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1062(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1063(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1064(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1401(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1402(.a(gate242inter0), .b(s_122), .O(gate242inter1));
  and2  gate1403(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1404(.a(s_122), .O(gate242inter3));
  inv1  gate1405(.a(s_123), .O(gate242inter4));
  nand2 gate1406(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1407(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1408(.a(G718), .O(gate242inter7));
  inv1  gate1409(.a(G730), .O(gate242inter8));
  nand2 gate1410(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1411(.a(s_123), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1412(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1413(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1414(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1947(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1948(.a(gate243inter0), .b(s_200), .O(gate243inter1));
  and2  gate1949(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1950(.a(s_200), .O(gate243inter3));
  inv1  gate1951(.a(s_201), .O(gate243inter4));
  nand2 gate1952(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1953(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1954(.a(G245), .O(gate243inter7));
  inv1  gate1955(.a(G733), .O(gate243inter8));
  nand2 gate1956(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1957(.a(s_201), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1958(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1959(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1960(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate897(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate898(.a(gate246inter0), .b(s_50), .O(gate246inter1));
  and2  gate899(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate900(.a(s_50), .O(gate246inter3));
  inv1  gate901(.a(s_51), .O(gate246inter4));
  nand2 gate902(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate903(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate904(.a(G724), .O(gate246inter7));
  inv1  gate905(.a(G736), .O(gate246inter8));
  nand2 gate906(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate907(.a(s_51), .b(gate246inter3), .O(gate246inter10));
  nor2  gate908(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate909(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate910(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate953(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate954(.a(gate248inter0), .b(s_58), .O(gate248inter1));
  and2  gate955(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate956(.a(s_58), .O(gate248inter3));
  inv1  gate957(.a(s_59), .O(gate248inter4));
  nand2 gate958(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate959(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate960(.a(G727), .O(gate248inter7));
  inv1  gate961(.a(G739), .O(gate248inter8));
  nand2 gate962(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate963(.a(s_59), .b(gate248inter3), .O(gate248inter10));
  nor2  gate964(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate965(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate966(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate925(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate926(.a(gate249inter0), .b(s_54), .O(gate249inter1));
  and2  gate927(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate928(.a(s_54), .O(gate249inter3));
  inv1  gate929(.a(s_55), .O(gate249inter4));
  nand2 gate930(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate931(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate932(.a(G254), .O(gate249inter7));
  inv1  gate933(.a(G742), .O(gate249inter8));
  nand2 gate934(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate935(.a(s_55), .b(gate249inter3), .O(gate249inter10));
  nor2  gate936(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate937(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate938(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1443(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1444(.a(gate252inter0), .b(s_128), .O(gate252inter1));
  and2  gate1445(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1446(.a(s_128), .O(gate252inter3));
  inv1  gate1447(.a(s_129), .O(gate252inter4));
  nand2 gate1448(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1449(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1450(.a(G709), .O(gate252inter7));
  inv1  gate1451(.a(G745), .O(gate252inter8));
  nand2 gate1452(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1453(.a(s_129), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1454(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1455(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1456(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate1569(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1570(.a(gate253inter0), .b(s_146), .O(gate253inter1));
  and2  gate1571(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1572(.a(s_146), .O(gate253inter3));
  inv1  gate1573(.a(s_147), .O(gate253inter4));
  nand2 gate1574(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1575(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1576(.a(G260), .O(gate253inter7));
  inv1  gate1577(.a(G748), .O(gate253inter8));
  nand2 gate1578(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1579(.a(s_147), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1580(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1581(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1582(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1723(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1724(.a(gate259inter0), .b(s_168), .O(gate259inter1));
  and2  gate1725(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1726(.a(s_168), .O(gate259inter3));
  inv1  gate1727(.a(s_169), .O(gate259inter4));
  nand2 gate1728(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1729(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1730(.a(G758), .O(gate259inter7));
  inv1  gate1731(.a(G759), .O(gate259inter8));
  nand2 gate1732(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1733(.a(s_169), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1734(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1735(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1736(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1037(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1038(.a(gate260inter0), .b(s_70), .O(gate260inter1));
  and2  gate1039(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1040(.a(s_70), .O(gate260inter3));
  inv1  gate1041(.a(s_71), .O(gate260inter4));
  nand2 gate1042(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1043(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1044(.a(G760), .O(gate260inter7));
  inv1  gate1045(.a(G761), .O(gate260inter8));
  nand2 gate1046(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1047(.a(s_71), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1048(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1049(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1050(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2171(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2172(.a(gate262inter0), .b(s_232), .O(gate262inter1));
  and2  gate2173(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2174(.a(s_232), .O(gate262inter3));
  inv1  gate2175(.a(s_233), .O(gate262inter4));
  nand2 gate2176(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2177(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2178(.a(G764), .O(gate262inter7));
  inv1  gate2179(.a(G765), .O(gate262inter8));
  nand2 gate2180(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2181(.a(s_233), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2182(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2183(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2184(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1359(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1360(.a(gate267inter0), .b(s_116), .O(gate267inter1));
  and2  gate1361(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1362(.a(s_116), .O(gate267inter3));
  inv1  gate1363(.a(s_117), .O(gate267inter4));
  nand2 gate1364(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1365(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1366(.a(G648), .O(gate267inter7));
  inv1  gate1367(.a(G776), .O(gate267inter8));
  nand2 gate1368(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1369(.a(s_117), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1370(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1371(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1372(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1317(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1318(.a(gate270inter0), .b(s_110), .O(gate270inter1));
  and2  gate1319(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1320(.a(s_110), .O(gate270inter3));
  inv1  gate1321(.a(s_111), .O(gate270inter4));
  nand2 gate1322(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1323(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1324(.a(G657), .O(gate270inter7));
  inv1  gate1325(.a(G785), .O(gate270inter8));
  nand2 gate1326(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1327(.a(s_111), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1328(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1329(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1330(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1891(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1892(.a(gate277inter0), .b(s_192), .O(gate277inter1));
  and2  gate1893(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1894(.a(s_192), .O(gate277inter3));
  inv1  gate1895(.a(s_193), .O(gate277inter4));
  nand2 gate1896(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1897(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1898(.a(G648), .O(gate277inter7));
  inv1  gate1899(.a(G800), .O(gate277inter8));
  nand2 gate1900(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1901(.a(s_193), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1902(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1903(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1904(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1709(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1710(.a(gate279inter0), .b(s_166), .O(gate279inter1));
  and2  gate1711(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1712(.a(s_166), .O(gate279inter3));
  inv1  gate1713(.a(s_167), .O(gate279inter4));
  nand2 gate1714(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1715(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1716(.a(G651), .O(gate279inter7));
  inv1  gate1717(.a(G803), .O(gate279inter8));
  nand2 gate1718(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1719(.a(s_167), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1720(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1721(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1722(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate687(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate688(.a(gate285inter0), .b(s_20), .O(gate285inter1));
  and2  gate689(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate690(.a(s_20), .O(gate285inter3));
  inv1  gate691(.a(s_21), .O(gate285inter4));
  nand2 gate692(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate693(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate694(.a(G660), .O(gate285inter7));
  inv1  gate695(.a(G812), .O(gate285inter8));
  nand2 gate696(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate697(.a(s_21), .b(gate285inter3), .O(gate285inter10));
  nor2  gate698(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate699(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate700(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1079(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1080(.a(gate294inter0), .b(s_76), .O(gate294inter1));
  and2  gate1081(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1082(.a(s_76), .O(gate294inter3));
  inv1  gate1083(.a(s_77), .O(gate294inter4));
  nand2 gate1084(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1085(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1086(.a(G832), .O(gate294inter7));
  inv1  gate1087(.a(G833), .O(gate294inter8));
  nand2 gate1088(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1089(.a(s_77), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1090(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1091(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1092(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate799(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate800(.a(gate295inter0), .b(s_36), .O(gate295inter1));
  and2  gate801(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate802(.a(s_36), .O(gate295inter3));
  inv1  gate803(.a(s_37), .O(gate295inter4));
  nand2 gate804(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate805(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate806(.a(G830), .O(gate295inter7));
  inv1  gate807(.a(G831), .O(gate295inter8));
  nand2 gate808(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate809(.a(s_37), .b(gate295inter3), .O(gate295inter10));
  nor2  gate810(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate811(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate812(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1065(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1066(.a(gate397inter0), .b(s_74), .O(gate397inter1));
  and2  gate1067(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1068(.a(s_74), .O(gate397inter3));
  inv1  gate1069(.a(s_75), .O(gate397inter4));
  nand2 gate1070(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1071(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1072(.a(G11), .O(gate397inter7));
  inv1  gate1073(.a(G1066), .O(gate397inter8));
  nand2 gate1074(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1075(.a(s_75), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1076(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1077(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1078(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2423(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2424(.a(gate398inter0), .b(s_268), .O(gate398inter1));
  and2  gate2425(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2426(.a(s_268), .O(gate398inter3));
  inv1  gate2427(.a(s_269), .O(gate398inter4));
  nand2 gate2428(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2429(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2430(.a(G12), .O(gate398inter7));
  inv1  gate2431(.a(G1069), .O(gate398inter8));
  nand2 gate2432(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2433(.a(s_269), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2434(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2435(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2436(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate617(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate618(.a(gate402inter0), .b(s_10), .O(gate402inter1));
  and2  gate619(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate620(.a(s_10), .O(gate402inter3));
  inv1  gate621(.a(s_11), .O(gate402inter4));
  nand2 gate622(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate623(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate624(.a(G16), .O(gate402inter7));
  inv1  gate625(.a(G1081), .O(gate402inter8));
  nand2 gate626(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate627(.a(s_11), .b(gate402inter3), .O(gate402inter10));
  nor2  gate628(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate629(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate630(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2479(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2480(.a(gate407inter0), .b(s_276), .O(gate407inter1));
  and2  gate2481(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2482(.a(s_276), .O(gate407inter3));
  inv1  gate2483(.a(s_277), .O(gate407inter4));
  nand2 gate2484(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2485(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2486(.a(G21), .O(gate407inter7));
  inv1  gate2487(.a(G1096), .O(gate407inter8));
  nand2 gate2488(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2489(.a(s_277), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2490(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2491(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2492(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate589(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate590(.a(gate409inter0), .b(s_6), .O(gate409inter1));
  and2  gate591(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate592(.a(s_6), .O(gate409inter3));
  inv1  gate593(.a(s_7), .O(gate409inter4));
  nand2 gate594(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate595(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate596(.a(G23), .O(gate409inter7));
  inv1  gate597(.a(G1102), .O(gate409inter8));
  nand2 gate598(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate599(.a(s_7), .b(gate409inter3), .O(gate409inter10));
  nor2  gate600(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate601(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate602(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate869(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate870(.a(gate410inter0), .b(s_46), .O(gate410inter1));
  and2  gate871(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate872(.a(s_46), .O(gate410inter3));
  inv1  gate873(.a(s_47), .O(gate410inter4));
  nand2 gate874(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate875(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate876(.a(G24), .O(gate410inter7));
  inv1  gate877(.a(G1105), .O(gate410inter8));
  nand2 gate878(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate879(.a(s_47), .b(gate410inter3), .O(gate410inter10));
  nor2  gate880(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate881(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate882(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2465(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2466(.a(gate413inter0), .b(s_274), .O(gate413inter1));
  and2  gate2467(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2468(.a(s_274), .O(gate413inter3));
  inv1  gate2469(.a(s_275), .O(gate413inter4));
  nand2 gate2470(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2471(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2472(.a(G27), .O(gate413inter7));
  inv1  gate2473(.a(G1114), .O(gate413inter8));
  nand2 gate2474(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2475(.a(s_275), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2476(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2477(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2478(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1597(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1598(.a(gate415inter0), .b(s_150), .O(gate415inter1));
  and2  gate1599(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1600(.a(s_150), .O(gate415inter3));
  inv1  gate1601(.a(s_151), .O(gate415inter4));
  nand2 gate1602(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1603(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1604(.a(G29), .O(gate415inter7));
  inv1  gate1605(.a(G1120), .O(gate415inter8));
  nand2 gate1606(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1607(.a(s_151), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1608(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1609(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1610(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1093(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1094(.a(gate416inter0), .b(s_78), .O(gate416inter1));
  and2  gate1095(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1096(.a(s_78), .O(gate416inter3));
  inv1  gate1097(.a(s_79), .O(gate416inter4));
  nand2 gate1098(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1099(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1100(.a(G30), .O(gate416inter7));
  inv1  gate1101(.a(G1123), .O(gate416inter8));
  nand2 gate1102(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1103(.a(s_79), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1104(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1105(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1106(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2003(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2004(.a(gate418inter0), .b(s_208), .O(gate418inter1));
  and2  gate2005(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2006(.a(s_208), .O(gate418inter3));
  inv1  gate2007(.a(s_209), .O(gate418inter4));
  nand2 gate2008(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2009(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2010(.a(G32), .O(gate418inter7));
  inv1  gate2011(.a(G1129), .O(gate418inter8));
  nand2 gate2012(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2013(.a(s_209), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2014(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2015(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2016(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2157(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2158(.a(gate420inter0), .b(s_230), .O(gate420inter1));
  and2  gate2159(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2160(.a(s_230), .O(gate420inter3));
  inv1  gate2161(.a(s_231), .O(gate420inter4));
  nand2 gate2162(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2163(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2164(.a(G1036), .O(gate420inter7));
  inv1  gate2165(.a(G1132), .O(gate420inter8));
  nand2 gate2166(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2167(.a(s_231), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2168(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2169(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2170(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1989(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1990(.a(gate426inter0), .b(s_206), .O(gate426inter1));
  and2  gate1991(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1992(.a(s_206), .O(gate426inter3));
  inv1  gate1993(.a(s_207), .O(gate426inter4));
  nand2 gate1994(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1995(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1996(.a(G1045), .O(gate426inter7));
  inv1  gate1997(.a(G1141), .O(gate426inter8));
  nand2 gate1998(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1999(.a(s_207), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2000(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2001(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2002(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1667(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1668(.a(gate430inter0), .b(s_160), .O(gate430inter1));
  and2  gate1669(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1670(.a(s_160), .O(gate430inter3));
  inv1  gate1671(.a(s_161), .O(gate430inter4));
  nand2 gate1672(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1673(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1674(.a(G1051), .O(gate430inter7));
  inv1  gate1675(.a(G1147), .O(gate430inter8));
  nand2 gate1676(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1677(.a(s_161), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1678(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1679(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1680(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2269(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2270(.a(gate431inter0), .b(s_246), .O(gate431inter1));
  and2  gate2271(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2272(.a(s_246), .O(gate431inter3));
  inv1  gate2273(.a(s_247), .O(gate431inter4));
  nand2 gate2274(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2275(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2276(.a(G7), .O(gate431inter7));
  inv1  gate2277(.a(G1150), .O(gate431inter8));
  nand2 gate2278(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2279(.a(s_247), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2280(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2281(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2282(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1121(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1122(.a(gate432inter0), .b(s_82), .O(gate432inter1));
  and2  gate1123(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1124(.a(s_82), .O(gate432inter3));
  inv1  gate1125(.a(s_83), .O(gate432inter4));
  nand2 gate1126(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1127(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1128(.a(G1054), .O(gate432inter7));
  inv1  gate1129(.a(G1150), .O(gate432inter8));
  nand2 gate1130(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1131(.a(s_83), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1132(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1133(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1134(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1653(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1654(.a(gate434inter0), .b(s_158), .O(gate434inter1));
  and2  gate1655(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1656(.a(s_158), .O(gate434inter3));
  inv1  gate1657(.a(s_159), .O(gate434inter4));
  nand2 gate1658(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1659(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1660(.a(G1057), .O(gate434inter7));
  inv1  gate1661(.a(G1153), .O(gate434inter8));
  nand2 gate1662(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1663(.a(s_159), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1664(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1665(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1666(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1583(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1584(.a(gate436inter0), .b(s_148), .O(gate436inter1));
  and2  gate1585(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1586(.a(s_148), .O(gate436inter3));
  inv1  gate1587(.a(s_149), .O(gate436inter4));
  nand2 gate1588(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1589(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1590(.a(G1060), .O(gate436inter7));
  inv1  gate1591(.a(G1156), .O(gate436inter8));
  nand2 gate1592(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1593(.a(s_149), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1594(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1595(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1596(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1191(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1192(.a(gate437inter0), .b(s_92), .O(gate437inter1));
  and2  gate1193(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1194(.a(s_92), .O(gate437inter3));
  inv1  gate1195(.a(s_93), .O(gate437inter4));
  nand2 gate1196(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1197(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1198(.a(G10), .O(gate437inter7));
  inv1  gate1199(.a(G1159), .O(gate437inter8));
  nand2 gate1200(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1201(.a(s_93), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1202(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1203(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1204(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1513(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1514(.a(gate438inter0), .b(s_138), .O(gate438inter1));
  and2  gate1515(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1516(.a(s_138), .O(gate438inter3));
  inv1  gate1517(.a(s_139), .O(gate438inter4));
  nand2 gate1518(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1519(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1520(.a(G1063), .O(gate438inter7));
  inv1  gate1521(.a(G1159), .O(gate438inter8));
  nand2 gate1522(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1523(.a(s_139), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1524(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1525(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1526(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2325(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2326(.a(gate442inter0), .b(s_254), .O(gate442inter1));
  and2  gate2327(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2328(.a(s_254), .O(gate442inter3));
  inv1  gate2329(.a(s_255), .O(gate442inter4));
  nand2 gate2330(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2331(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2332(.a(G1069), .O(gate442inter7));
  inv1  gate2333(.a(G1165), .O(gate442inter8));
  nand2 gate2334(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2335(.a(s_255), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2336(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2337(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2338(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate2115(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2116(.a(gate443inter0), .b(s_224), .O(gate443inter1));
  and2  gate2117(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2118(.a(s_224), .O(gate443inter3));
  inv1  gate2119(.a(s_225), .O(gate443inter4));
  nand2 gate2120(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2121(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2122(.a(G13), .O(gate443inter7));
  inv1  gate2123(.a(G1168), .O(gate443inter8));
  nand2 gate2124(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2125(.a(s_225), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2126(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2127(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2128(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate575(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate576(.a(gate455inter0), .b(s_4), .O(gate455inter1));
  and2  gate577(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate578(.a(s_4), .O(gate455inter3));
  inv1  gate579(.a(s_5), .O(gate455inter4));
  nand2 gate580(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate581(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate582(.a(G19), .O(gate455inter7));
  inv1  gate583(.a(G1186), .O(gate455inter8));
  nand2 gate584(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate585(.a(s_5), .b(gate455inter3), .O(gate455inter10));
  nor2  gate586(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate587(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate588(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1849(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1850(.a(gate459inter0), .b(s_186), .O(gate459inter1));
  and2  gate1851(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1852(.a(s_186), .O(gate459inter3));
  inv1  gate1853(.a(s_187), .O(gate459inter4));
  nand2 gate1854(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1855(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1856(.a(G21), .O(gate459inter7));
  inv1  gate1857(.a(G1192), .O(gate459inter8));
  nand2 gate1858(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1859(.a(s_187), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1860(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1861(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1862(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate813(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate814(.a(gate464inter0), .b(s_38), .O(gate464inter1));
  and2  gate815(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate816(.a(s_38), .O(gate464inter3));
  inv1  gate817(.a(s_39), .O(gate464inter4));
  nand2 gate818(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate819(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate820(.a(G1102), .O(gate464inter7));
  inv1  gate821(.a(G1198), .O(gate464inter8));
  nand2 gate822(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate823(.a(s_39), .b(gate464inter3), .O(gate464inter10));
  nor2  gate824(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate825(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate826(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate967(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate968(.a(gate470inter0), .b(s_60), .O(gate470inter1));
  and2  gate969(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate970(.a(s_60), .O(gate470inter3));
  inv1  gate971(.a(s_61), .O(gate470inter4));
  nand2 gate972(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate973(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate974(.a(G1111), .O(gate470inter7));
  inv1  gate975(.a(G1207), .O(gate470inter8));
  nand2 gate976(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate977(.a(s_61), .b(gate470inter3), .O(gate470inter10));
  nor2  gate978(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate979(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate980(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1933(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1934(.a(gate479inter0), .b(s_198), .O(gate479inter1));
  and2  gate1935(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1936(.a(s_198), .O(gate479inter3));
  inv1  gate1937(.a(s_199), .O(gate479inter4));
  nand2 gate1938(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1939(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1940(.a(G31), .O(gate479inter7));
  inv1  gate1941(.a(G1222), .O(gate479inter8));
  nand2 gate1942(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1943(.a(s_199), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1944(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1945(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1946(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate2087(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2088(.a(gate480inter0), .b(s_220), .O(gate480inter1));
  and2  gate2089(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2090(.a(s_220), .O(gate480inter3));
  inv1  gate2091(.a(s_221), .O(gate480inter4));
  nand2 gate2092(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2093(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2094(.a(G1126), .O(gate480inter7));
  inv1  gate2095(.a(G1222), .O(gate480inter8));
  nand2 gate2096(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2097(.a(s_221), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2098(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2099(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2100(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate827(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate828(.a(gate481inter0), .b(s_40), .O(gate481inter1));
  and2  gate829(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate830(.a(s_40), .O(gate481inter3));
  inv1  gate831(.a(s_41), .O(gate481inter4));
  nand2 gate832(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate833(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate834(.a(G32), .O(gate481inter7));
  inv1  gate835(.a(G1225), .O(gate481inter8));
  nand2 gate836(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate837(.a(s_41), .b(gate481inter3), .O(gate481inter10));
  nor2  gate838(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate839(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate840(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1863(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1864(.a(gate483inter0), .b(s_188), .O(gate483inter1));
  and2  gate1865(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1866(.a(s_188), .O(gate483inter3));
  inv1  gate1867(.a(s_189), .O(gate483inter4));
  nand2 gate1868(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1869(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1870(.a(G1228), .O(gate483inter7));
  inv1  gate1871(.a(G1229), .O(gate483inter8));
  nand2 gate1872(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1873(.a(s_189), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1874(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1875(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1876(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1387(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1388(.a(gate492inter0), .b(s_120), .O(gate492inter1));
  and2  gate1389(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1390(.a(s_120), .O(gate492inter3));
  inv1  gate1391(.a(s_121), .O(gate492inter4));
  nand2 gate1392(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1393(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1394(.a(G1246), .O(gate492inter7));
  inv1  gate1395(.a(G1247), .O(gate492inter8));
  nand2 gate1396(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1397(.a(s_121), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1398(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1399(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1400(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1527(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1528(.a(gate497inter0), .b(s_140), .O(gate497inter1));
  and2  gate1529(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1530(.a(s_140), .O(gate497inter3));
  inv1  gate1531(.a(s_141), .O(gate497inter4));
  nand2 gate1532(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1533(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1534(.a(G1256), .O(gate497inter7));
  inv1  gate1535(.a(G1257), .O(gate497inter8));
  nand2 gate1536(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1537(.a(s_141), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1538(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1539(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1540(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1415(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1416(.a(gate498inter0), .b(s_124), .O(gate498inter1));
  and2  gate1417(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1418(.a(s_124), .O(gate498inter3));
  inv1  gate1419(.a(s_125), .O(gate498inter4));
  nand2 gate1420(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1421(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1422(.a(G1258), .O(gate498inter7));
  inv1  gate1423(.a(G1259), .O(gate498inter8));
  nand2 gate1424(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1425(.a(s_125), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1426(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1427(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1428(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate673(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate674(.a(gate502inter0), .b(s_18), .O(gate502inter1));
  and2  gate675(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate676(.a(s_18), .O(gate502inter3));
  inv1  gate677(.a(s_19), .O(gate502inter4));
  nand2 gate678(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate679(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate680(.a(G1266), .O(gate502inter7));
  inv1  gate681(.a(G1267), .O(gate502inter8));
  nand2 gate682(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate683(.a(s_19), .b(gate502inter3), .O(gate502inter10));
  nor2  gate684(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate685(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate686(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1737(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1738(.a(gate503inter0), .b(s_170), .O(gate503inter1));
  and2  gate1739(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1740(.a(s_170), .O(gate503inter3));
  inv1  gate1741(.a(s_171), .O(gate503inter4));
  nand2 gate1742(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1743(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1744(.a(G1268), .O(gate503inter7));
  inv1  gate1745(.a(G1269), .O(gate503inter8));
  nand2 gate1746(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1747(.a(s_171), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1748(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1749(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1750(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1205(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1206(.a(gate507inter0), .b(s_94), .O(gate507inter1));
  and2  gate1207(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1208(.a(s_94), .O(gate507inter3));
  inv1  gate1209(.a(s_95), .O(gate507inter4));
  nand2 gate1210(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1211(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1212(.a(G1276), .O(gate507inter7));
  inv1  gate1213(.a(G1277), .O(gate507inter8));
  nand2 gate1214(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1215(.a(s_95), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1216(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1217(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1218(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1149(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1150(.a(gate510inter0), .b(s_86), .O(gate510inter1));
  and2  gate1151(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1152(.a(s_86), .O(gate510inter3));
  inv1  gate1153(.a(s_87), .O(gate510inter4));
  nand2 gate1154(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1155(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1156(.a(G1282), .O(gate510inter7));
  inv1  gate1157(.a(G1283), .O(gate510inter8));
  nand2 gate1158(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1159(.a(s_87), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1160(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1161(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1162(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1345(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1346(.a(gate513inter0), .b(s_114), .O(gate513inter1));
  and2  gate1347(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1348(.a(s_114), .O(gate513inter3));
  inv1  gate1349(.a(s_115), .O(gate513inter4));
  nand2 gate1350(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1351(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1352(.a(G1288), .O(gate513inter7));
  inv1  gate1353(.a(G1289), .O(gate513inter8));
  nand2 gate1354(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1355(.a(s_115), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1356(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1357(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1358(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule