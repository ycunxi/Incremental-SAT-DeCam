module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate310inter0, gate310inter1, gate310inter2, gate310inter3, gate310inter4, gate310inter5, gate310inter6, gate310inter7, gate310inter8, gate310inter9, gate310inter10, gate310inter11, gate310inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate301inter0, gate301inter1, gate301inter2, gate301inter3, gate301inter4, gate301inter5, gate301inter6, gate301inter7, gate301inter8, gate301inter9, gate301inter10, gate301inter11, gate301inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate302inter0, gate302inter1, gate302inter2, gate302inter3, gate302inter4, gate302inter5, gate302inter6, gate302inter7, gate302inter8, gate302inter9, gate302inter10, gate302inter11, gate302inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12;



nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );
nand2 gate20( .a(N91), .b(N96), .O(N301) );
or2 gate21( .a(N91), .b(N96), .O(N302) );
nand2 gate22( .a(N101), .b(N106), .O(N303) );
or2 gate23( .a(N101), .b(N106), .O(N304) );
nand2 gate24( .a(N111), .b(N116), .O(N305) );
or2 gate25( .a(N111), .b(N116), .O(N306) );
nand2 gate26( .a(N121), .b(N126), .O(N307) );
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );

  xor2  gate622(.a(N156), .b(N59), .O(gate33inter0));
  nand2 gate623(.a(gate33inter0), .b(s_34), .O(gate33inter1));
  and2  gate624(.a(N156), .b(N59), .O(gate33inter2));
  inv1  gate625(.a(s_34), .O(gate33inter3));
  inv1  gate626(.a(s_35), .O(gate33inter4));
  nand2 gate627(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate628(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate629(.a(N59), .O(gate33inter7));
  inv1  gate630(.a(N156), .O(gate33inter8));
  nand2 gate631(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate632(.a(s_35), .b(gate33inter3), .O(gate33inter10));
  nor2  gate633(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate634(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate635(.a(gate33inter12), .b(gate33inter1), .O(N319));
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17), .b(N42), .O(N323) );
nand2 gate36( .a(N159), .b(N165), .O(N324) );
or2 gate37( .a(N159), .b(N165), .O(N325) );
nand2 gate38( .a(N171), .b(N177), .O(N326) );
or2 gate39( .a(N171), .b(N177), .O(N327) );

  xor2  gate440(.a(N189), .b(N183), .O(gate40inter0));
  nand2 gate441(.a(gate40inter0), .b(s_8), .O(gate40inter1));
  and2  gate442(.a(N189), .b(N183), .O(gate40inter2));
  inv1  gate443(.a(s_8), .O(gate40inter3));
  inv1  gate444(.a(s_9), .O(gate40inter4));
  nand2 gate445(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate446(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate447(.a(N183), .O(gate40inter7));
  inv1  gate448(.a(N189), .O(gate40inter8));
  nand2 gate449(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate450(.a(s_9), .b(gate40inter3), .O(gate40inter10));
  nor2  gate451(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate452(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate453(.a(gate40inter12), .b(gate40inter1), .O(N328));
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
and2 gate49( .a(N255), .b(N259), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );
nor2 gate60( .a(N280), .b(N284), .O(N348) );
or2 gate61( .a(N280), .b(N285), .O(N349) );
or2 gate62( .a(N280), .b(N286), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );
nand2 gate67( .a(N89), .b(N298), .O(N355) );
and2 gate68( .a(N90), .b(N298), .O(N356) );

  xor2  gate720(.a(N302), .b(N301), .O(gate69inter0));
  nand2 gate721(.a(gate69inter0), .b(s_48), .O(gate69inter1));
  and2  gate722(.a(N302), .b(N301), .O(gate69inter2));
  inv1  gate723(.a(s_48), .O(gate69inter3));
  inv1  gate724(.a(s_49), .O(gate69inter4));
  nand2 gate725(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate726(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate727(.a(N301), .O(gate69inter7));
  inv1  gate728(.a(N302), .O(gate69inter8));
  nand2 gate729(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate730(.a(s_49), .b(gate69inter3), .O(gate69inter10));
  nor2  gate731(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate732(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate733(.a(gate69inter12), .b(gate69inter1), .O(N357));
nand2 gate70( .a(N303), .b(N304), .O(N360) );

  xor2  gate706(.a(N306), .b(N305), .O(gate71inter0));
  nand2 gate707(.a(gate71inter0), .b(s_46), .O(gate71inter1));
  and2  gate708(.a(N306), .b(N305), .O(gate71inter2));
  inv1  gate709(.a(s_46), .O(gate71inter3));
  inv1  gate710(.a(s_47), .O(gate71inter4));
  nand2 gate711(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate712(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate713(.a(N305), .O(gate71inter7));
  inv1  gate714(.a(N306), .O(gate71inter8));
  nand2 gate715(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate716(.a(s_47), .b(gate71inter3), .O(gate71inter10));
  nor2  gate717(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate718(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate719(.a(gate71inter12), .b(gate71inter1), .O(N363));
nand2 gate72( .a(N307), .b(N308), .O(N366) );
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );

  xor2  gate580(.a(N327), .b(N326), .O(gate76inter0));
  nand2 gate581(.a(gate76inter0), .b(s_28), .O(gate76inter1));
  and2  gate582(.a(N327), .b(N326), .O(gate76inter2));
  inv1  gate583(.a(s_28), .O(gate76inter3));
  inv1  gate584(.a(s_29), .O(gate76inter4));
  nand2 gate585(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate586(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate587(.a(N326), .O(gate76inter7));
  inv1  gate588(.a(N327), .O(gate76inter8));
  nand2 gate589(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate590(.a(s_29), .b(gate76inter3), .O(gate76inter10));
  nor2  gate591(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate592(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate593(.a(gate76inter12), .b(gate76inter1), .O(N379));
nand2 gate77( .a(N328), .b(N329), .O(N382) );
nand2 gate78( .a(N330), .b(N331), .O(N385) );
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );

  xor2  gate524(.a(N352), .b(N347), .O(gate96inter0));
  nand2 gate525(.a(gate96inter0), .b(s_20), .O(gate96inter1));
  and2  gate526(.a(N352), .b(N347), .O(gate96inter2));
  inv1  gate527(.a(s_20), .O(gate96inter3));
  inv1  gate528(.a(s_21), .O(gate96inter4));
  nand2 gate529(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate530(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate531(.a(N347), .O(gate96inter7));
  inv1  gate532(.a(N352), .O(gate96inter8));
  nand2 gate533(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate534(.a(s_21), .b(gate96inter3), .O(gate96inter10));
  nor2  gate535(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate536(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate537(.a(gate96inter12), .b(gate96inter1), .O(N410));
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );

  xor2  gate594(.a(N425), .b(N406), .O(gate126inter0));
  nand2 gate595(.a(gate126inter0), .b(s_30), .O(gate126inter1));
  and2  gate596(.a(N425), .b(N406), .O(gate126inter2));
  inv1  gate597(.a(s_30), .O(gate126inter3));
  inv1  gate598(.a(s_31), .O(gate126inter4));
  nand2 gate599(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate600(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate601(.a(N406), .O(gate126inter7));
  inv1  gate602(.a(N425), .O(gate126inter8));
  nand2 gate603(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate604(.a(s_31), .b(gate126inter3), .O(gate126inter10));
  nor2  gate605(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate606(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate607(.a(gate126inter12), .b(gate126inter1), .O(N460));
nor2 gate127( .a(N409), .b(N426), .O(N463) );

  xor2  gate692(.a(N410), .b(N442), .O(gate128inter0));
  nand2 gate693(.a(gate128inter0), .b(s_44), .O(gate128inter1));
  and2  gate694(.a(N410), .b(N442), .O(gate128inter2));
  inv1  gate695(.a(s_44), .O(gate128inter3));
  inv1  gate696(.a(s_45), .O(gate128inter4));
  nand2 gate697(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate698(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate699(.a(N442), .O(gate128inter7));
  inv1  gate700(.a(N410), .O(gate128inter8));
  nand2 gate701(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate702(.a(s_45), .b(gate128inter3), .O(gate128inter10));
  nor2  gate703(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate704(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate705(.a(gate128inter12), .b(gate128inter1), .O(N466));
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );
nand2 gate137( .a(N443), .b(N1), .O(N483) );
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );
nor2 gate142( .a(N413), .b(N444), .O(N492) );

  xor2  gate608(.a(N445), .b(N416), .O(gate143inter0));
  nand2 gate609(.a(gate143inter0), .b(s_32), .O(gate143inter1));
  and2  gate610(.a(N445), .b(N416), .O(gate143inter2));
  inv1  gate611(.a(s_32), .O(gate143inter3));
  inv1  gate612(.a(s_33), .O(gate143inter4));
  nand2 gate613(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate614(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate615(.a(N416), .O(gate143inter7));
  inv1  gate616(.a(N445), .O(gate143inter8));
  nand2 gate617(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate618(.a(s_33), .b(gate143inter3), .O(gate143inter10));
  nor2  gate619(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate620(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate621(.a(gate143inter12), .b(gate143inter1), .O(N495));
nand2 gate144( .a(N130), .b(N460), .O(N498) );
or2 gate145( .a(N130), .b(N460), .O(N499) );
nand2 gate146( .a(N463), .b(N135), .O(N500) );
or2 gate147( .a(N463), .b(N135), .O(N501) );
and2 gate148( .a(N91), .b(N466), .O(N502) );
nor2 gate149( .a(N475), .b(N476), .O(N503) );
and2 gate150( .a(N96), .b(N466), .O(N504) );
nor2 gate151( .a(N477), .b(N478), .O(N505) );
and2 gate152( .a(N101), .b(N466), .O(N506) );

  xor2  gate538(.a(N480), .b(N479), .O(gate153inter0));
  nand2 gate539(.a(gate153inter0), .b(s_22), .O(gate153inter1));
  and2  gate540(.a(N480), .b(N479), .O(gate153inter2));
  inv1  gate541(.a(s_22), .O(gate153inter3));
  inv1  gate542(.a(s_23), .O(gate153inter4));
  nand2 gate543(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate544(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate545(.a(N479), .O(gate153inter7));
  inv1  gate546(.a(N480), .O(gate153inter8));
  nand2 gate547(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate548(.a(s_23), .b(gate153inter3), .O(gate153inter10));
  nor2  gate549(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate550(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate551(.a(gate153inter12), .b(gate153inter1), .O(N507));
and2 gate154( .a(N106), .b(N466), .O(N508) );
nor2 gate155( .a(N481), .b(N482), .O(N509) );
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );
nand2 gate164( .a(N130), .b(N492), .O(N518) );
or2 gate165( .a(N130), .b(N492), .O(N519) );

  xor2  gate664(.a(N207), .b(N495), .O(gate166inter0));
  nand2 gate665(.a(gate166inter0), .b(s_40), .O(gate166inter1));
  and2  gate666(.a(N207), .b(N495), .O(gate166inter2));
  inv1  gate667(.a(s_40), .O(gate166inter3));
  inv1  gate668(.a(s_41), .O(gate166inter4));
  nand2 gate669(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate670(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate671(.a(N495), .O(gate166inter7));
  inv1  gate672(.a(N207), .O(gate166inter8));
  nand2 gate673(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate674(.a(s_41), .b(gate166inter3), .O(gate166inter10));
  nor2  gate675(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate676(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate677(.a(gate166inter12), .b(gate166inter1), .O(N520));
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
and2 gate170( .a(N451), .b(N171), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );
nand2 gate173( .a(N451), .b(N189), .O(N527) );
nand2 gate174( .a(N451), .b(N195), .O(N528) );
nand2 gate175( .a(N451), .b(N201), .O(N529) );

  xor2  gate482(.a(N499), .b(N498), .O(gate176inter0));
  nand2 gate483(.a(gate176inter0), .b(s_14), .O(gate176inter1));
  and2  gate484(.a(N499), .b(N498), .O(gate176inter2));
  inv1  gate485(.a(s_14), .O(gate176inter3));
  inv1  gate486(.a(s_15), .O(gate176inter4));
  nand2 gate487(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate488(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate489(.a(N498), .O(gate176inter7));
  inv1  gate490(.a(N499), .O(gate176inter8));
  nand2 gate491(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate492(.a(s_15), .b(gate176inter3), .O(gate176inter10));
  nor2  gate493(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate494(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate495(.a(gate176inter12), .b(gate176inter1), .O(N530));
nand2 gate177( .a(N500), .b(N501), .O(N533) );
nor2 gate178( .a(N309), .b(N502), .O(N536) );
nor2 gate179( .a(N316), .b(N504), .O(N537) );
nor2 gate180( .a(N317), .b(N506), .O(N538) );
nor2 gate181( .a(N318), .b(N508), .O(N539) );

  xor2  gate454(.a(N511), .b(N510), .O(gate182inter0));
  nand2 gate455(.a(gate182inter0), .b(s_10), .O(gate182inter1));
  and2  gate456(.a(N511), .b(N510), .O(gate182inter2));
  inv1  gate457(.a(s_10), .O(gate182inter3));
  inv1  gate458(.a(s_11), .O(gate182inter4));
  nand2 gate459(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate460(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate461(.a(N510), .O(gate182inter7));
  inv1  gate462(.a(N511), .O(gate182inter8));
  nand2 gate463(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate464(.a(s_11), .b(gate182inter3), .O(gate182inter10));
  nor2  gate465(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate466(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate467(.a(gate182inter12), .b(gate182inter1), .O(N540));
nor2 gate183( .a(N512), .b(N513), .O(N541) );
nor2 gate184( .a(N514), .b(N515), .O(N542) );
nor2 gate185( .a(N516), .b(N517), .O(N543) );
nand2 gate186( .a(N518), .b(N519), .O(N544) );
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );
nand2 gate191( .a(N536), .b(N503), .O(N553) );
nand2 gate192( .a(N537), .b(N505), .O(N557) );
nand2 gate193( .a(N538), .b(N507), .O(N561) );
nand2 gate194( .a(N539), .b(N509), .O(N565) );

  xor2  gate566(.a(N540), .b(N488), .O(gate195inter0));
  nand2 gate567(.a(gate195inter0), .b(s_26), .O(gate195inter1));
  and2  gate568(.a(N540), .b(N488), .O(gate195inter2));
  inv1  gate569(.a(s_26), .O(gate195inter3));
  inv1  gate570(.a(s_27), .O(gate195inter4));
  nand2 gate571(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate572(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate573(.a(N488), .O(gate195inter7));
  inv1  gate574(.a(N540), .O(gate195inter8));
  nand2 gate575(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate576(.a(s_27), .b(gate195inter3), .O(gate195inter10));
  nor2  gate577(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate578(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate579(.a(gate195inter12), .b(gate195inter1), .O(N569));
nand2 gate196( .a(N489), .b(N541), .O(N573) );
nand2 gate197( .a(N490), .b(N542), .O(N577) );
nand2 gate198( .a(N491), .b(N543), .O(N581) );
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );
nand2 gate204( .a(N553), .b(N159), .O(N590) );
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );

  xor2  gate468(.a(N165), .b(N557), .O(gate207inter0));
  nand2 gate469(.a(gate207inter0), .b(s_12), .O(gate207inter1));
  and2  gate470(.a(N165), .b(N557), .O(gate207inter2));
  inv1  gate471(.a(s_12), .O(gate207inter3));
  inv1  gate472(.a(s_13), .O(gate207inter4));
  nand2 gate473(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate474(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate475(.a(N557), .O(gate207inter7));
  inv1  gate476(.a(N165), .O(gate207inter8));
  nand2 gate477(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate478(.a(s_13), .b(gate207inter3), .O(gate207inter10));
  nor2  gate479(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate480(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate481(.a(gate207inter12), .b(gate207inter1), .O(N597));
or2 gate208( .a(N557), .b(N165), .O(N600) );
and2 gate209( .a(N246), .b(N557), .O(N605) );
nand2 gate210( .a(N561), .b(N171), .O(N606) );
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );
nand2 gate213( .a(N565), .b(N177), .O(N616) );
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );
nand2 gate216( .a(N569), .b(N183), .O(N625) );
or2 gate217( .a(N569), .b(N183), .O(N628) );
and2 gate218( .a(N246), .b(N569), .O(N631) );

  xor2  gate650(.a(N189), .b(N573), .O(gate219inter0));
  nand2 gate651(.a(gate219inter0), .b(s_38), .O(gate219inter1));
  and2  gate652(.a(N189), .b(N573), .O(gate219inter2));
  inv1  gate653(.a(s_38), .O(gate219inter3));
  inv1  gate654(.a(s_39), .O(gate219inter4));
  nand2 gate655(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate656(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate657(.a(N573), .O(gate219inter7));
  inv1  gate658(.a(N189), .O(gate219inter8));
  nand2 gate659(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate660(.a(s_39), .b(gate219inter3), .O(gate219inter10));
  nor2  gate661(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate662(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate663(.a(gate219inter12), .b(gate219inter1), .O(N632));
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );

  xor2  gate398(.a(N195), .b(N577), .O(gate222inter0));
  nand2 gate399(.a(gate222inter0), .b(s_2), .O(gate222inter1));
  and2  gate400(.a(N195), .b(N577), .O(gate222inter2));
  inv1  gate401(.a(s_2), .O(gate222inter3));
  inv1  gate402(.a(s_3), .O(gate222inter4));
  nand2 gate403(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate404(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate405(.a(N577), .O(gate222inter7));
  inv1  gate406(.a(N195), .O(gate222inter8));
  nand2 gate407(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate408(.a(s_3), .b(gate222inter3), .O(gate222inter10));
  nor2  gate409(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate410(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate411(.a(gate222inter12), .b(gate222inter1), .O(N641));
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );
nand2 gate225( .a(N581), .b(N201), .O(N651) );
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );
nor2 gate228( .a(N552), .b(N588), .O(N660) );
nor2 gate229( .a(N587), .b(N589), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
and2 gate231( .a(N593), .b(N590), .O(N665) );
nor2 gate232( .a(N596), .b(N522), .O(N669) );
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );
nor2 gate235( .a(N605), .b(N523), .O(N677) );
inv1 gate236( .a(N606), .O(N678) );
and2 gate237( .a(N609), .b(N606), .O(N682) );
nor2 gate238( .a(N615), .b(N524), .O(N686) );
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );

  xor2  gate552(.a(N525), .b(N624), .O(gate241inter0));
  nand2 gate553(.a(gate241inter0), .b(s_24), .O(gate241inter1));
  and2  gate554(.a(N525), .b(N624), .O(gate241inter2));
  inv1  gate555(.a(s_24), .O(gate241inter3));
  inv1  gate556(.a(s_25), .O(gate241inter4));
  nand2 gate557(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate558(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate559(.a(N624), .O(gate241inter7));
  inv1  gate560(.a(N525), .O(gate241inter8));
  nand2 gate561(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate562(.a(s_25), .b(gate241inter3), .O(gate241inter10));
  nor2  gate563(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate564(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate565(.a(gate241inter12), .b(gate241inter1), .O(N696));
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );
nor2 gate244( .a(N631), .b(N526), .O(N704) );
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );
nor2 gate247( .a(N337), .b(N640), .O(N712) );
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );

  xor2  gate510(.a(N650), .b(N339), .O(gate250inter0));
  nand2 gate511(.a(gate250inter0), .b(s_18), .O(gate250inter1));
  and2  gate512(.a(N650), .b(N339), .O(gate250inter2));
  inv1  gate513(.a(s_18), .O(gate250inter3));
  inv1  gate514(.a(s_19), .O(gate250inter4));
  nand2 gate515(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate516(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate517(.a(N339), .O(gate250inter7));
  inv1  gate518(.a(N650), .O(gate250inter8));
  nand2 gate519(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate520(.a(s_19), .b(gate250inter3), .O(gate250inter10));
  nor2  gate521(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate522(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate523(.a(gate250inter12), .b(gate250inter1), .O(N721));
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );

  xor2  gate734(.a(N659), .b(N341), .O(gate253inter0));
  nand2 gate735(.a(gate253inter0), .b(s_50), .O(gate253inter1));
  and2  gate736(.a(N659), .b(N341), .O(gate253inter2));
  inv1  gate737(.a(s_50), .O(gate253inter3));
  inv1  gate738(.a(s_51), .O(gate253inter4));
  nand2 gate739(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate740(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate741(.a(N341), .O(gate253inter7));
  inv1  gate742(.a(N659), .O(gate253inter8));
  nand2 gate743(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate744(.a(s_51), .b(gate253inter3), .O(gate253inter10));
  nor2  gate745(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate746(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate747(.a(gate253inter12), .b(gate253inter1), .O(N731));
nand2 gate254( .a(N654), .b(N261), .O(N732) );
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
and2 gate273( .a(N228), .b(N708), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );

  xor2  gate384(.a(N261), .b(N727), .O(gate279inter0));
  nand2 gate385(.a(gate279inter0), .b(s_0), .O(gate279inter1));
  and2  gate386(.a(N261), .b(N727), .O(gate279inter2));
  inv1  gate387(.a(s_0), .O(gate279inter3));
  inv1  gate388(.a(s_1), .O(gate279inter4));
  nand2 gate389(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate390(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate391(.a(N727), .O(gate279inter7));
  inv1  gate392(.a(N261), .O(gate279inter8));
  nand2 gate393(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate394(.a(s_1), .b(gate279inter3), .O(gate279inter10));
  nor2  gate395(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate396(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate397(.a(gate279inter12), .b(gate279inter1), .O(N757));
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );
nand2 gate284( .a(N635), .b(N713), .O(N762) );
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );
nor2 gate291( .a(N736), .b(N737), .O(N769) );
nor2 gate292( .a(N739), .b(N740), .O(N770) );

  xor2  gate412(.a(N743), .b(N742), .O(gate293inter0));
  nand2 gate413(.a(gate293inter0), .b(s_4), .O(gate293inter1));
  and2  gate414(.a(N743), .b(N742), .O(gate293inter2));
  inv1  gate415(.a(s_4), .O(gate293inter3));
  inv1  gate416(.a(s_5), .O(gate293inter4));
  nand2 gate417(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate418(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate419(.a(N742), .O(gate293inter7));
  inv1  gate420(.a(N743), .O(gate293inter8));
  nand2 gate421(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate422(.a(s_5), .b(gate293inter3), .O(gate293inter10));
  nor2  gate423(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate424(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate425(.a(gate293inter12), .b(gate293inter1), .O(N771));
nor2 gate294( .a(N745), .b(N746), .O(N772) );
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );
nor2 gate296( .a(N748), .b(N749), .O(N777) );
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );
nor2 gate298( .a(N751), .b(N752), .O(N781) );
nand2 gate299( .a(N756), .b(N732), .O(N782) );
nor2 gate300( .a(N754), .b(N755), .O(N785) );

  xor2  gate636(.a(N758), .b(N757), .O(gate301inter0));
  nand2 gate637(.a(gate301inter0), .b(s_36), .O(gate301inter1));
  and2  gate638(.a(N758), .b(N757), .O(gate301inter2));
  inv1  gate639(.a(s_36), .O(gate301inter3));
  inv1  gate640(.a(s_37), .O(gate301inter4));
  nand2 gate641(.a(gate301inter4), .b(gate301inter3), .O(gate301inter5));
  nor2  gate642(.a(gate301inter5), .b(gate301inter2), .O(gate301inter6));
  inv1  gate643(.a(N757), .O(gate301inter7));
  inv1  gate644(.a(N758), .O(gate301inter8));
  nand2 gate645(.a(gate301inter8), .b(gate301inter7), .O(gate301inter9));
  nand2 gate646(.a(s_37), .b(gate301inter3), .O(gate301inter10));
  nor2  gate647(.a(gate301inter10), .b(gate301inter9), .O(gate301inter11));
  nor2  gate648(.a(gate301inter11), .b(gate301inter6), .O(gate301inter12));
  nand2 gate649(.a(gate301inter12), .b(gate301inter1), .O(N786));

  xor2  gate678(.a(N760), .b(N759), .O(gate302inter0));
  nand2 gate679(.a(gate302inter0), .b(s_42), .O(gate302inter1));
  and2  gate680(.a(N760), .b(N759), .O(gate302inter2));
  inv1  gate681(.a(s_42), .O(gate302inter3));
  inv1  gate682(.a(s_43), .O(gate302inter4));
  nand2 gate683(.a(gate302inter4), .b(gate302inter3), .O(gate302inter5));
  nor2  gate684(.a(gate302inter5), .b(gate302inter2), .O(gate302inter6));
  inv1  gate685(.a(N759), .O(gate302inter7));
  inv1  gate686(.a(N760), .O(gate302inter8));
  nand2 gate687(.a(gate302inter8), .b(gate302inter7), .O(gate302inter9));
  nand2 gate688(.a(s_43), .b(gate302inter3), .O(gate302inter10));
  nor2  gate689(.a(gate302inter10), .b(gate302inter9), .O(gate302inter11));
  nor2  gate690(.a(gate302inter11), .b(gate302inter6), .O(gate302inter12));
  nand2 gate691(.a(gate302inter12), .b(gate302inter1), .O(N787));
nor2 gate303( .a(N700), .b(N773), .O(N788) );
and2 gate304( .a(N700), .b(N773), .O(N789) );
nor2 gate305( .a(N708), .b(N778), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );
nor2 gate307( .a(N717), .b(N782), .O(N792) );
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );

  xor2  gate426(.a(N773), .b(N628), .O(gate310inter0));
  nand2 gate427(.a(gate310inter0), .b(s_6), .O(gate310inter1));
  and2  gate428(.a(N773), .b(N628), .O(gate310inter2));
  inv1  gate429(.a(s_6), .O(gate310inter3));
  inv1  gate430(.a(s_7), .O(gate310inter4));
  nand2 gate431(.a(gate310inter4), .b(gate310inter3), .O(gate310inter5));
  nor2  gate432(.a(gate310inter5), .b(gate310inter2), .O(gate310inter6));
  inv1  gate433(.a(N628), .O(gate310inter7));
  inv1  gate434(.a(N773), .O(gate310inter8));
  nand2 gate435(.a(gate310inter8), .b(gate310inter7), .O(gate310inter9));
  nand2 gate436(.a(s_7), .b(gate310inter3), .O(gate310inter10));
  nor2  gate437(.a(gate310inter10), .b(gate310inter9), .O(gate310inter11));
  nor2  gate438(.a(gate310inter11), .b(gate310inter6), .O(gate310inter12));
  nand2 gate439(.a(gate310inter12), .b(gate310inter1), .O(N795));
nand2 gate311( .a(N795), .b(N747), .O(N796) );
nor2 gate312( .a(N788), .b(N789), .O(N802) );
nor2 gate313( .a(N790), .b(N791), .O(N803) );

  xor2  gate496(.a(N793), .b(N792), .O(gate314inter0));
  nand2 gate497(.a(gate314inter0), .b(s_16), .O(gate314inter1));
  and2  gate498(.a(N793), .b(N792), .O(gate314inter2));
  inv1  gate499(.a(s_16), .O(gate314inter3));
  inv1  gate500(.a(s_17), .O(gate314inter4));
  nand2 gate501(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate502(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate503(.a(N792), .O(gate314inter7));
  inv1  gate504(.a(N793), .O(gate314inter8));
  nand2 gate505(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate506(.a(s_17), .b(gate314inter3), .O(gate314inter10));
  nor2  gate507(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate508(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate509(.a(gate314inter12), .b(gate314inter1), .O(N804));
nor2 gate315( .a(N340), .b(N794), .O(N805) );
nor2 gate316( .a(N692), .b(N796), .O(N806) );
and2 gate317( .a(N692), .b(N796), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );
nand2 gate322( .a(N619), .b(N796), .O(N812) );
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );
nand2 gate327( .a(N744), .b(N812), .O(N822) );
nor2 gate328( .a(N806), .b(N807), .O(N825) );
nor2 gate329( .a(N335), .b(N808), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );
nor2 gate333( .a(N665), .b(N815), .O(N830) );
and2 gate334( .a(N665), .b(N815), .O(N831) );
nor2 gate335( .a(N673), .b(N819), .O(N832) );
and2 gate336( .a(N673), .b(N819), .O(N833) );
nor2 gate337( .a(N682), .b(N822), .O(N834) );
and2 gate338( .a(N682), .b(N822), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
nand2 gate344( .a(N815), .b(N593), .O(N841) );
nor2 gate345( .a(N830), .b(N831), .O(N842) );
nor2 gate346( .a(N832), .b(N833), .O(N843) );
nor2 gate347( .a(N834), .b(N835), .O(N844) );
nor2 gate348( .a(N334), .b(N836), .O(N845) );
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
and2 gate354( .a(N219), .b(N842), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );
nor2 gate362( .a(N417), .b(N851), .O(N859) );
nor2 gate363( .a(N332), .b(N852), .O(N860) );
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

endmodule